//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G106gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G50gat), .B(G78gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT29), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT78), .A3(G141gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n213), .C1(G141gat), .C2(new_n212), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n218), .B2(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n210), .A2(G148gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n212), .A2(G141gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n218), .A2(new_n215), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n208), .B1(new_n227), .B2(KEYINPUT3), .ZN(new_n228));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G211gat), .A2(G218gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n229), .B1(new_n234), .B2(KEYINPUT73), .ZN(new_n235));
  OR2_X1    g034(.A1(G197gat), .A2(G204gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n236), .A2(new_n237), .B1(new_n232), .B2(new_n231), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT73), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n235), .A2(new_n240), .B1(new_n229), .B2(new_n238), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n228), .B(new_n243), .C1(new_n242), .C2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G228gat), .ZN(new_n246));
  INV_X1    g045(.A(G233gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT84), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT74), .B1(new_n235), .B2(new_n240), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n238), .A2(new_n229), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n241), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n251), .B1(new_n253), .B2(KEYINPUT74), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n250), .B1(new_n254), .B2(KEYINPUT29), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n242), .B1(new_n241), .B2(new_n252), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT84), .B(new_n208), .C1(new_n257), .C2(new_n251), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n249), .B1(new_n259), .B2(new_n227), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT83), .ZN(new_n261));
  INV_X1    g060(.A(new_n252), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n238), .A2(new_n229), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n208), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n227), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n248), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI211_X1 g068(.A(KEYINPUT83), .B(new_n248), .C1(new_n245), .C2(new_n266), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(G22gat), .B1(new_n260), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n258), .A2(new_n256), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n243), .B1(new_n244), .B2(new_n242), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT84), .B1(new_n274), .B2(new_n208), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n227), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n249), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n254), .A2(new_n228), .B1(new_n227), .B2(new_n265), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT83), .B1(new_n279), .B2(new_n248), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n267), .A2(new_n261), .A3(new_n268), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G22gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n278), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI211_X1 g083(.A(KEYINPUT85), .B(new_n207), .C1(new_n272), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n272), .A2(new_n284), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT85), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n206), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n284), .A3(KEYINPUT85), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G15gat), .B(G43gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G71gat), .B(G99gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n297), .A2(KEYINPUT67), .B1(new_n296), .B2(new_n295), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n299), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  OAI211_X1 g104(.A(KEYINPUT66), .B(KEYINPUT28), .C1(new_n305), .C2(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  AOI21_X1  g107(.A(G190gat), .B1(new_n302), .B2(new_n303), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n301), .A2(new_n306), .A3(new_n307), .A4(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(G183gat), .B(G190gat), .C1(KEYINPUT65), .C2(KEYINPUT24), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT65), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n315), .B(new_n318), .C1(new_n307), .C2(new_n314), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n321), .A2(new_n294), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT25), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n318), .A2(KEYINPUT24), .A3(new_n307), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT25), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n325), .B(new_n326), .C1(KEYINPUT24), .C2(new_n307), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n320), .A2(new_n294), .A3(new_n321), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G113gat), .B(G120gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT1), .ZN(new_n333));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT68), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n334), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT68), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n336), .B(new_n337), .C1(KEYINPUT1), .C2(new_n332), .ZN(new_n338));
  XOR2_X1   g137(.A(KEYINPUT69), .B(KEYINPUT1), .Z(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(new_n332), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n335), .A2(new_n338), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n331), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n329), .B1(KEYINPUT25), .B2(new_n323), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n341), .B1(new_n344), .B2(new_n312), .ZN(new_n345));
  OAI211_X1 g144(.A(G227gat), .B(G233gat), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT33), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n293), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n350));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n342), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n344), .A2(new_n341), .A3(new_n312), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT32), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n348), .A2(new_n349), .A3(new_n356), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n346), .B(KEYINPUT32), .C1(new_n347), .C2(new_n293), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT34), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n352), .A2(new_n360), .A3(new_n353), .A4(new_n351), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n361), .A2(KEYINPUT71), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(KEYINPUT71), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n352), .A2(new_n351), .A3(new_n353), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT34), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT72), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n359), .A2(new_n366), .ZN(new_n368));
  INV_X1    g167(.A(new_n366), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n358), .A3(new_n357), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n371), .B2(KEYINPUT72), .ZN(new_n372));
  INV_X1    g171(.A(G226gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(new_n247), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n331), .B2(new_n208), .ZN(new_n375));
  INV_X1    g174(.A(new_n374), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n344), .B2(new_n312), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n254), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n331), .A2(new_n374), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n344), .B2(new_n312), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n379), .B(new_n274), .C1(new_n380), .C2(new_n374), .ZN(new_n381));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT75), .ZN(new_n383));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n378), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT76), .B(KEYINPUT30), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT77), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n390), .A3(new_n387), .ZN(new_n391));
  INV_X1    g190(.A(new_n385), .ZN(new_n392));
  INV_X1    g191(.A(new_n378), .ZN(new_n393));
  INV_X1    g192(.A(new_n381), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n378), .A2(KEYINPUT30), .A3(new_n381), .A4(new_n385), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n389), .A2(new_n391), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n335), .A2(new_n338), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n214), .A2(new_n219), .B1(new_n224), .B2(new_n225), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n340), .A2(new_n334), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT81), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT4), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n341), .B(KEYINPUT79), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n400), .B(KEYINPUT3), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n406), .A2(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(KEYINPUT5), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n404), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n398), .A2(KEYINPUT79), .A3(new_n401), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT79), .B1(new_n398), .B2(new_n401), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n227), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT80), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT80), .B(new_n227), .C1(new_n416), .C2(new_n417), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n411), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n409), .B1(new_n416), .B2(new_n417), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n402), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n411), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT5), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n414), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428));
  INV_X1    g227(.A(G85gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT0), .B(G57gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434));
  INV_X1    g233(.A(new_n432), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(new_n414), .C1(new_n422), .C2(new_n426), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n397), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n290), .A2(new_n372), .A3(new_n439), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n260), .A2(new_n271), .A3(G22gat), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n283), .B1(new_n278), .B2(new_n282), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n287), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n207), .A3(new_n289), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n286), .A2(new_n287), .A3(new_n206), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(new_n371), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n439), .A2(KEYINPUT35), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n202), .A2(new_n440), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT40), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT39), .B1(new_n410), .B2(new_n411), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n418), .A2(new_n419), .ZN(new_n452));
  AND4_X1   g251(.A1(new_n411), .A2(new_n452), .A3(new_n421), .A4(new_n404), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n406), .A2(new_n407), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n423), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT39), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n412), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n435), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n450), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n420), .A2(new_n411), .A3(new_n421), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(KEYINPUT39), .C1(new_n411), .C2(new_n410), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n462), .A2(KEYINPUT40), .A3(new_n435), .A4(new_n458), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n397), .A2(new_n460), .A3(new_n433), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n437), .A2(new_n438), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT37), .B1(new_n393), .B2(new_n394), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT37), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n378), .A2(new_n381), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n392), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT38), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT38), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n466), .A2(new_n471), .A3(new_n392), .A4(new_n468), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n386), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n464), .B1(new_n465), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT87), .B1(new_n474), .B2(new_n446), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n472), .A2(new_n386), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n477), .A2(new_n437), .A3(new_n438), .A4(new_n470), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n290), .A2(new_n476), .A3(new_n478), .A4(new_n464), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT36), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(new_n372), .B2(KEYINPUT36), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n444), .B2(new_n445), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n290), .A2(new_n483), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n439), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n449), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G232gat), .A2(G233gat), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT41), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(G162gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT92), .B(G134gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n496));
  INV_X1    g295(.A(G29gat), .ZN(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT14), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n497), .A3(new_n498), .ZN(new_n502));
  AOI211_X1 g301(.A(new_n496), .B(new_n499), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n502), .A2(new_n500), .B1(G29gat), .B2(G36gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n495), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n507));
  INV_X1    g306(.A(new_n495), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT17), .ZN(new_n511));
  XOR2_X1   g310(.A(G99gat), .B(G106gat), .Z(new_n512));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT8), .ZN(new_n514));
  OR2_X1    g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n514), .A2(KEYINPUT95), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT95), .B1(new_n514), .B2(new_n515), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT94), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(KEYINPUT93), .A2(KEYINPUT94), .A3(KEYINPUT7), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  AND3_X1   g324(.A1(KEYINPUT93), .A2(KEYINPUT94), .A3(KEYINPUT7), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT94), .B1(KEYINPUT93), .B2(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n529));
  OAI22_X1  g328(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n512), .B1(new_n518), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n525), .A2(new_n530), .ZN(new_n533));
  INV_X1    g332(.A(new_n512), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT95), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT8), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n536), .B1(G99gat), .B2(G106gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(G85gat), .A2(G92gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT95), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n533), .A2(new_n534), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n532), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n506), .A2(new_n544), .A3(new_n509), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n511), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT96), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n511), .A2(new_n548), .A3(new_n543), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n490), .A2(KEYINPUT41), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n510), .B2(new_n543), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G190gat), .B(G218gat), .Z(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(new_n557), .A3(new_n553), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n494), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n550), .B2(new_n553), .ZN(new_n560));
  AOI211_X1 g359(.A(new_n555), .B(new_n552), .C1(new_n547), .C2(new_n549), .ZN(new_n561));
  INV_X1    g360(.A(new_n494), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT16), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(G1gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(G1gat), .B2(new_n565), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G8gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  OR2_X1    g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n573), .B(new_n572), .C1(new_n570), .C2(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n569), .B1(KEYINPUT21), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n579), .B(KEYINPUT21), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n569), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT91), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(new_n316), .ZN(new_n586));
  INV_X1    g385(.A(G211gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n583), .B(new_n588), .Z(new_n589));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n589), .B(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n564), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n518), .A2(new_n531), .A3(new_n512), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n534), .B1(new_n533), .B2(new_n541), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n579), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n532), .A2(new_n580), .A3(new_n542), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n532), .A2(new_n542), .A3(KEYINPUT10), .A4(new_n580), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT97), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n601), .A2(new_n603), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n608), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n598), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT99), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT98), .B1(new_n606), .B2(new_n609), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616));
  AOI211_X1 g415(.A(new_n616), .B(new_n608), .C1(new_n604), .C2(new_n605), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n598), .B(new_n612), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(G8gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n568), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n511), .A2(new_n622), .A3(new_n545), .ZN(new_n623));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n510), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n569), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n623), .A2(KEYINPUT18), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n628));
  XNOR2_X1  g427(.A(G113gat), .B(G141gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G169gat), .B(G197gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n624), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n625), .A2(new_n569), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n622), .A2(new_n510), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n627), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT90), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(KEYINPUT90), .A3(new_n641), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n639), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n640), .A2(KEYINPUT89), .A3(new_n641), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT89), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g448(.A1(new_n647), .A2(new_n649), .A3(new_n638), .A4(new_n627), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n646), .B1(new_n650), .B2(new_n633), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n594), .A2(new_n620), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n488), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n465), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT100), .B(G1gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1324gat));
  INV_X1    g455(.A(new_n397), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n621), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT101), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT16), .B(G8gat), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT42), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(G1325gat));
  INV_X1    g463(.A(new_n653), .ZN(new_n665));
  INV_X1    g464(.A(new_n481), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n665), .A2(G15gat), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(G15gat), .B1(new_n665), .B2(new_n372), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(G1326gat));
  NAND2_X1  g468(.A1(new_n485), .A2(new_n486), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT102), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT43), .B(G22gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  INV_X1    g473(.A(new_n564), .ZN(new_n675));
  INV_X1    g474(.A(new_n439), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n444), .A2(new_n483), .A3(new_n445), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n677), .B2(new_n484), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n678), .A2(new_n479), .A3(new_n481), .A4(new_n475), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n679), .B2(new_n449), .ZN(new_n680));
  INV_X1    g479(.A(new_n651), .ZN(new_n681));
  INV_X1    g480(.A(new_n593), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n681), .A2(new_n682), .A3(new_n619), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n465), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n497), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT45), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n488), .B2(new_n564), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n559), .B2(new_n563), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n556), .A2(new_n494), .A3(new_n558), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n562), .B1(new_n560), .B2(new_n561), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT104), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  AOI211_X1 g495(.A(KEYINPUT44), .B(new_n696), .C1(new_n679), .C2(new_n449), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n689), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT103), .Z(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n685), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n687), .B1(new_n701), .B2(new_n497), .ZN(G1328gat));
  NAND3_X1  g501(.A1(new_n684), .A2(new_n498), .A3(new_n397), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT46), .Z(new_n704));
  NAND3_X1  g503(.A1(new_n698), .A2(new_n397), .A3(new_n699), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n498), .B2(new_n706), .ZN(G1329gat));
  INV_X1    g506(.A(G43gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n684), .A2(new_n708), .A3(new_n372), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n666), .B(new_n699), .C1(new_n689), .C2(new_n697), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(new_n708), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1330gat));
  OAI211_X1 g513(.A(new_n446), .B(new_n699), .C1(new_n689), .C2(new_n697), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G50gat), .ZN(new_n716));
  INV_X1    g515(.A(G50gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n684), .A2(new_n717), .A3(new_n670), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(KEYINPUT48), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n716), .A2(KEYINPUT105), .A3(KEYINPUT48), .A4(new_n718), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n670), .B(new_n699), .C1(new_n689), .C2(new_n697), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G50gat), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n724), .A2(new_n718), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n721), .B(new_n722), .C1(KEYINPUT48), .C2(new_n725), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n594), .A2(new_n681), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n679), .B2(new_n449), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n465), .A2(new_n620), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT106), .B(G57gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1332gat));
  INV_X1    g531(.A(KEYINPUT49), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n728), .A2(new_n619), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n657), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(KEYINPUT107), .ZN(new_n737));
  INV_X1    g536(.A(G64gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(KEYINPUT107), .ZN(new_n739));
  AND4_X1   g538(.A1(new_n733), .A2(new_n737), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n737), .A2(new_n739), .B1(new_n733), .B2(new_n738), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(new_n734), .B2(new_n666), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n372), .A2(new_n743), .A3(new_n619), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n728), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n734), .A2(new_n670), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT108), .B(G78gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n682), .A2(new_n651), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n488), .A2(new_n564), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n429), .A3(new_n729), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n620), .A2(new_n682), .A3(new_n651), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n698), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n685), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n755), .B1(new_n759), .B2(new_n429), .ZN(G1336gat));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n752), .A2(new_n761), .A3(KEYINPUT51), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n620), .A2(G92gat), .A3(new_n657), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT109), .B1(new_n680), .B2(new_n751), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n762), .B(new_n763), .C1(KEYINPUT51), .C2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n761), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n753), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n769), .A2(KEYINPUT110), .A3(new_n762), .A4(new_n763), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n397), .B(new_n756), .C1(new_n689), .C2(new_n697), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n767), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(new_n754), .B2(new_n763), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1337gat));
  INV_X1    g576(.A(G99gat), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n754), .A2(new_n778), .A3(new_n372), .A4(new_n619), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n757), .A2(new_n666), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(new_n778), .ZN(G1338gat));
  NOR3_X1   g581(.A1(new_n290), .A2(new_n620), .A3(G106gat), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n769), .A2(new_n762), .A3(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n670), .B(new_n756), .C1(new_n689), .C2(new_n697), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(G106gat), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT53), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT53), .B1(new_n754), .B2(new_n783), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n446), .B(new_n756), .C1(new_n689), .C2(new_n697), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(KEYINPUT111), .ZN(new_n790));
  OAI21_X1  g589(.A(G106gat), .B1(new_n789), .B2(KEYINPUT111), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(new_n792), .ZN(G1339gat));
  NAND3_X1  g592(.A1(new_n604), .A2(new_n608), .A3(new_n605), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(KEYINPUT54), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n615), .B2(new_n617), .ZN(new_n796));
  AOI211_X1 g595(.A(KEYINPUT54), .B(new_n608), .C1(new_n604), .C2(new_n605), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n797), .A2(KEYINPUT112), .A3(new_n598), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n606), .A2(new_n800), .A3(new_n609), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n799), .B1(new_n801), .B2(new_n597), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n796), .B(KEYINPUT55), .C1(new_n798), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n618), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(KEYINPUT113), .A3(new_n618), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT112), .B1(new_n797), .B2(new_n598), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n801), .A2(new_n799), .A3(new_n597), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT55), .B1(new_n810), .B2(new_n796), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n806), .A2(new_n651), .A3(new_n807), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n624), .B1(new_n623), .B2(new_n626), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n636), .A2(new_n637), .A3(new_n635), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n632), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n619), .A2(new_n646), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n695), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n811), .B1(new_n804), .B2(new_n805), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n646), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n646), .B2(new_n816), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND4_X1   g622(.A1(new_n695), .A2(new_n819), .A3(new_n807), .A4(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n593), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n594), .A2(new_n620), .A3(new_n681), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n670), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n465), .A2(new_n397), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(new_n372), .A3(new_n828), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT115), .Z(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n681), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n825), .A2(new_n826), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n447), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n828), .ZN(new_n835));
  INV_X1    g634(.A(G113gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n651), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n837), .ZN(G1340gat));
  OAI21_X1  g637(.A(G120gat), .B1(new_n831), .B2(new_n620), .ZN(new_n839));
  INV_X1    g638(.A(G120gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n835), .A2(new_n840), .A3(new_n619), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(G1341gat));
  AOI21_X1  g641(.A(G127gat), .B1(new_n835), .B2(new_n682), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n682), .A2(G127gat), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n830), .B2(new_n844), .ZN(G1342gat));
  INV_X1    g644(.A(G134gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n835), .A2(new_n846), .A3(new_n564), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT56), .Z(new_n848));
  OAI21_X1  g647(.A(G134gat), .B1(new_n831), .B2(new_n675), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n481), .A2(new_n828), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n290), .B1(new_n825), .B2(new_n826), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(KEYINPUT57), .ZN(new_n855));
  INV_X1    g654(.A(new_n824), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n651), .A2(new_n812), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n817), .B1(new_n857), .B2(new_n804), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n675), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n682), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n826), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n670), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n854), .A2(new_n853), .A3(KEYINPUT57), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n651), .B(new_n852), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G141gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n854), .A2(new_n852), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n210), .A3(new_n651), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT58), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n866), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n212), .A2(KEYINPUT59), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n852), .B1(new_n863), .B2(new_n864), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n620), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n819), .A2(new_n823), .A3(new_n564), .A4(new_n807), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n682), .B1(new_n859), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n878), .B(new_n670), .C1(new_n880), .C2(new_n861), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n854), .B2(new_n878), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n852), .A2(new_n619), .ZN(new_n883));
  OAI21_X1  g682(.A(G148gat), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g683(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n868), .A2(new_n212), .A3(new_n619), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1345gat));
  OAI21_X1  g688(.A(new_n216), .B1(new_n867), .B2(new_n593), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n682), .A2(G155gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n876), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT118), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n876), .B2(new_n696), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n868), .A2(new_n217), .A3(new_n564), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n465), .A2(new_n397), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n834), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(G169gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n651), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n372), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT119), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n827), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904), .B2(new_n681), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n901), .A2(new_n905), .ZN(G1348gat));
  INV_X1    g705(.A(G176gat), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n904), .A2(new_n907), .A3(new_n620), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n899), .A2(new_n619), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n907), .ZN(G1349gat));
  NOR2_X1   g709(.A1(new_n593), .A2(new_n305), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n899), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n827), .A2(new_n682), .A3(new_n903), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G183gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(KEYINPUT121), .A3(KEYINPUT60), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n899), .A2(new_n911), .B1(new_n913), .B2(G183gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT120), .B1(new_n915), .B2(KEYINPUT60), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n918), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  OAI22_X1  g722(.A1(new_n916), .A2(new_n920), .B1(new_n921), .B2(new_n923), .ZN(G1350gat));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925));
  OAI21_X1  g724(.A(G190gat), .B1(new_n904), .B2(new_n675), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n927), .A2(KEYINPUT123), .A3(new_n928), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(new_n926), .B2(KEYINPUT61), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n929), .A2(new_n930), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n899), .A2(new_n317), .A3(new_n695), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1351gat));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n882), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n666), .A2(new_n897), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n882), .A2(new_n937), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n681), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n290), .A2(new_n657), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n481), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n465), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n945), .B2(new_n944), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(new_n833), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n681), .A2(G197gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n942), .B1(new_n952), .B2(new_n953), .ZN(G1352gat));
  INV_X1    g753(.A(G204gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n948), .A2(new_n955), .A3(new_n619), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT62), .Z(new_n957));
  OAI21_X1  g756(.A(G204gat), .B1(new_n941), .B2(new_n620), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1353gat));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n682), .ZN(new_n960));
  OAI21_X1  g759(.A(G211gat), .B1(new_n882), .B2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964));
  OAI211_X1 g763(.A(KEYINPUT63), .B(G211gat), .C1(new_n882), .C2(new_n960), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n965), .A2(new_n964), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n682), .A2(new_n587), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n966), .A2(new_n967), .B1(new_n952), .B2(new_n968), .ZN(G1354gat));
  INV_X1    g768(.A(G218gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n941), .A2(new_n970), .A3(new_n675), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n695), .B1(new_n950), .B2(new_n951), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(new_n970), .B2(new_n972), .ZN(G1355gat));
endmodule


