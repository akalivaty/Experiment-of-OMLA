//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1280, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  OAI21_X1  g0045(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G1), .A3(G13), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(new_n249), .A3(G274), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n246), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n251), .B1(G226), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G223), .A3(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(new_n259), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n262), .B1(G222), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n254), .B1(new_n267), .B2(new_n249), .ZN(new_n268));
  INV_X1    g0068(.A(G169), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n214), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n202), .A2(G50), .ZN(new_n273));
  OR3_X1    g0073(.A1(new_n273), .A2(KEYINPUT68), .A3(new_n206), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(new_n206), .A3(new_n256), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G150), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT68), .B1(new_n273), .B2(new_n206), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n274), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n283));
  INV_X1    g0083(.A(G58), .ZN(new_n284));
  OR3_X1    g0084(.A1(new_n284), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n206), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n272), .B1(new_n281), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G50), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n272), .B1(new_n205), .B2(G20), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(G50), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT69), .B(G179), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n270), .B(new_n294), .C1(new_n296), .C2(new_n268), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n294), .B(KEYINPUT9), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n268), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(G200), .B2(new_n268), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n299), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n298), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT73), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT14), .ZN(new_n309));
  INV_X1    g0109(.A(G232), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G1698), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n311), .B1(G226), .B2(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n249), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n250), .B1(new_n219), .B2(new_n252), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT13), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT13), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n309), .B(G169), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n314), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n249), .A2(G274), .ZN(new_n321));
  AOI22_X1  g0121(.A1(G238), .A2(new_n253), .B1(new_n321), .B2(new_n247), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(G179), .A3(new_n316), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n316), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n309), .B1(new_n327), .B2(G169), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n308), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(G169), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT14), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n331), .A2(KEYINPUT73), .A3(new_n325), .A4(new_n319), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n272), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n278), .A2(G50), .ZN(new_n335));
  INV_X1    g0135(.A(new_n287), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(G77), .B1(G20), .B2(new_n218), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(KEYINPUT11), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(KEYINPUT11), .ZN(new_n340));
  OR3_X1    g0140(.A1(new_n290), .A2(KEYINPUT12), .A3(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT12), .B1(new_n290), .B2(G68), .ZN(new_n342));
  AOI22_X1  g0142(.A1(G68), .A2(new_n292), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n333), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n327), .A2(G200), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n300), .B2(new_n327), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n292), .A2(G77), .ZN(new_n351));
  INV_X1    g0151(.A(new_n290), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n261), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT8), .B(G58), .Z(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT15), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G87), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n356), .A2(KEYINPUT71), .B1(new_n336), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(KEYINPUT71), .B2(new_n356), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n354), .B1(new_n362), .B2(new_n272), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G1698), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n259), .A2(G232), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n259), .A2(G238), .A3(G1698), .ZN(new_n367));
  INV_X1    g0167(.A(G107), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n259), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n249), .B1(new_n369), .B2(KEYINPUT70), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(KEYINPUT70), .B2(new_n369), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n251), .B1(G244), .B2(new_n253), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n364), .B1(G200), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(G190), .A3(new_n372), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n363), .B1(new_n373), .B2(new_n269), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n371), .A2(new_n295), .A3(new_n372), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n374), .A2(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n307), .A2(new_n346), .A3(new_n350), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n284), .A2(new_n218), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(new_n201), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n257), .A2(new_n206), .A3(new_n258), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n258), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n383), .B1(new_n388), .B2(G68), .ZN(new_n389));
  AOI211_X1 g0189(.A(KEYINPUT74), .B(new_n218), .C1(new_n386), .C2(new_n387), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT16), .B(new_n382), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT7), .B1(new_n265), .B2(new_n206), .ZN(new_n392));
  INV_X1    g0192(.A(new_n387), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n382), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(new_n397), .A3(new_n272), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n286), .A2(new_n290), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n286), .B2(new_n292), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT75), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT75), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n399), .B(new_n402), .C1(new_n286), .C2(new_n292), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n250), .B1(new_n310), .B2(new_n252), .ZN(new_n406));
  INV_X1    g0206(.A(G223), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n365), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(G226), .B2(new_n365), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n409), .A2(new_n265), .B1(new_n256), .B2(new_n220), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n406), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n296), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n269), .B2(new_n412), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT18), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n405), .A2(new_n417), .A3(new_n414), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n300), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G200), .B2(new_n412), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n398), .A2(new_n420), .A3(new_n404), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n398), .A2(new_n420), .A3(KEYINPUT17), .A4(new_n404), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n416), .A2(new_n418), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n379), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G116), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n271), .A2(new_n214), .B1(G20), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G283), .ZN(new_n429));
  INV_X1    g0229(.A(G97), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(new_n206), .C1(G33), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT20), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n428), .A2(KEYINPUT20), .A3(new_n431), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n352), .A2(new_n427), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n205), .A2(G33), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n334), .A2(new_n290), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n436), .B(new_n437), .C1(new_n427), .C2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n259), .A2(G264), .A3(G1698), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n259), .A2(G257), .A3(new_n365), .ZN(new_n442));
  INV_X1    g0242(.A(G303), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n259), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n411), .ZN(new_n445));
  INV_X1    g0245(.A(G45), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  AND2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  NOR2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G270), .A3(new_n249), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT5), .B(G41), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(G274), .A3(new_n249), .A4(new_n447), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(KEYINPUT79), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT79), .B1(new_n451), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n445), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n440), .B1(new_n457), .B2(G200), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n300), .B2(new_n457), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT21), .ZN(new_n460));
  INV_X1    g0260(.A(new_n456), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n461), .A2(new_n454), .B1(new_n411), .B2(new_n444), .ZN(new_n462));
  INV_X1    g0262(.A(new_n436), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n437), .B1(new_n439), .B2(new_n427), .ZN(new_n464));
  OAI21_X1  g0264(.A(G169), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n460), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n457), .A2(new_n440), .A3(KEYINPUT21), .A4(G169), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(G179), .A3(new_n440), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n459), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n450), .A2(G257), .A3(new_n249), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n453), .ZN(new_n471));
  OAI211_X1 g0271(.A(G244), .B(new_n365), .C1(new_n263), .C2(new_n264), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n365), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n429), .A4(new_n476), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n300), .B(new_n471), .C1(new_n477), .C2(new_n411), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n278), .A2(G77), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n368), .A2(KEYINPUT6), .A3(G97), .ZN(new_n480));
  XNOR2_X1  g0280(.A(G97), .B(G107), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT6), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n479), .B1(new_n483), .B2(new_n206), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n368), .B1(new_n386), .B2(new_n387), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n272), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n290), .A2(G97), .ZN(new_n487));
  INV_X1    g0287(.A(new_n439), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(G97), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n478), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n477), .A2(new_n411), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT76), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n477), .A2(KEYINPUT76), .A3(new_n411), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n471), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G200), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n491), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n471), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(new_n269), .B1(new_n486), .B2(new_n489), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n477), .A2(KEYINPUT76), .A3(new_n411), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT76), .B1(new_n477), .B2(new_n411), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n295), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G116), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n206), .B2(G107), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n368), .A2(KEYINPUT23), .A3(G20), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n206), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n512), .A2(KEYINPUT22), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(KEYINPUT22), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(KEYINPUT24), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT24), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n512), .B(KEYINPUT22), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(new_n511), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n272), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT25), .B1(new_n352), .B2(new_n368), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n352), .A2(KEYINPUT25), .A3(new_n368), .ZN(new_n523));
  AOI22_X1  g0323(.A1(G107), .A2(new_n488), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XOR2_X1   g0324(.A(KEYINPUT80), .B(G294), .Z(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G33), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n259), .A2(G257), .A3(G1698), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n259), .A2(G250), .A3(new_n365), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n411), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n411), .B1(new_n447), .B2(new_n452), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G264), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n453), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(G190), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n529), .A2(new_n411), .B1(G264), .B2(new_n531), .ZN(new_n535));
  AOI21_X1  g0335(.A(G200), .B1(new_n535), .B2(new_n453), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n520), .B(new_n524), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n498), .A2(new_n505), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n533), .A2(new_n269), .ZN(new_n539));
  INV_X1    g0339(.A(G179), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n540), .A3(new_n453), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n515), .A2(KEYINPUT24), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n518), .A2(new_n517), .A3(new_n511), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n334), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n524), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n539), .B(new_n541), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT77), .ZN(new_n547));
  OAI21_X1  g0347(.A(G250), .B1(new_n446), .B2(G1), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n411), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n221), .B1(new_n205), .B2(G45), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(new_n249), .A3(KEYINPUT77), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n549), .A2(new_n551), .B1(new_n321), .B2(new_n447), .ZN(new_n552));
  OAI211_X1 g0352(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n553));
  OAI211_X1 g0353(.A(G238), .B(new_n365), .C1(new_n263), .C2(new_n264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(new_n506), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n411), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n552), .A2(new_n556), .A3(new_n295), .ZN(new_n557));
  AOI21_X1  g0357(.A(G169), .B1(new_n552), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n488), .A2(new_n360), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT78), .ZN(new_n561));
  NAND3_X1  g0361(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n206), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n220), .A2(new_n430), .A3(new_n368), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n206), .B(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n287), .B2(new_n430), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n272), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n360), .A2(new_n290), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n561), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AOI211_X1 g0373(.A(KEYINPUT78), .B(new_n571), .C1(new_n569), .C2(new_n272), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n560), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n559), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n555), .A2(new_n411), .ZN(new_n577));
  INV_X1    g0377(.A(new_n551), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT77), .B1(new_n550), .B2(new_n249), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n249), .A2(G274), .ZN(new_n580));
  INV_X1    g0380(.A(new_n447), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n578), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n497), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n552), .A2(new_n556), .A3(new_n300), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n570), .A2(new_n572), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n570), .A2(new_n561), .A3(new_n572), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n488), .A2(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n546), .A2(new_n576), .A3(new_n591), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n469), .A2(new_n538), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n426), .A2(new_n593), .ZN(G372));
  AND2_X1   g0394(.A1(new_n416), .A2(new_n418), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n376), .A2(new_n377), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n346), .B1(new_n349), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n423), .A2(new_n424), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n304), .A2(new_n306), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n297), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n426), .ZN(new_n605));
  INV_X1    g0405(.A(new_n546), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT82), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n468), .A2(new_n467), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT82), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n546), .A4(new_n466), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n587), .A2(new_n588), .B1(new_n360), .B2(new_n488), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n552), .A2(new_n556), .A3(new_n295), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n577), .A2(new_n582), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(G169), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n552), .A2(new_n556), .A3(new_n300), .ZN(new_n617));
  AOI21_X1  g0417(.A(G200), .B1(new_n552), .B2(new_n556), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n590), .B1(new_n573), .B2(new_n574), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n613), .A2(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT81), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n491), .B1(new_n504), .B2(new_n501), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT81), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n591), .A2(new_n576), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n622), .A2(new_n625), .A3(new_n537), .A4(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n576), .B1(new_n612), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n621), .A2(new_n505), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT26), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n505), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n622), .A2(new_n633), .A3(new_n627), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n632), .B1(new_n636), .B2(KEYINPUT83), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT83), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n634), .A2(new_n638), .A3(new_n635), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n629), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n604), .B1(new_n605), .B2(new_n640), .ZN(G369));
  NAND3_X1  g0441(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n645), .B(KEYINPUT84), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n607), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n544), .B2(new_n545), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n606), .B1(new_n652), .B2(new_n537), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n546), .A2(new_n649), .ZN(new_n654));
  OR3_X1    g0454(.A1(new_n653), .A2(KEYINPUT85), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(KEYINPUT85), .B1(new_n653), .B2(new_n654), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n654), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n649), .A2(new_n440), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n607), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n469), .B2(new_n660), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n658), .A2(new_n664), .ZN(G399));
  INV_X1    g0465(.A(new_n209), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(G41), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n205), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n564), .A2(G116), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n668), .A2(new_n669), .B1(new_n213), .B2(new_n667), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT28), .Z(new_n671));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n445), .B(G179), .C1(new_n455), .C2(new_n456), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n615), .A2(new_n535), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n471), .B1(new_n477), .B2(new_n411), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT30), .A4(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n615), .A2(new_n296), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n623), .A2(new_n533), .A3(new_n457), .A4(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT30), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n615), .A2(new_n676), .A3(new_n535), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n673), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n677), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT86), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n593), .A2(new_n650), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT31), .B1(new_n683), .B2(new_n649), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n687), .B1(KEYINPUT86), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n672), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n498), .A2(new_n505), .A3(new_n537), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n609), .A2(new_n466), .A3(new_n546), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n691), .A2(new_n622), .A3(new_n627), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n634), .A2(KEYINPUT26), .ZN(new_n694));
  INV_X1    g0494(.A(new_n576), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n630), .B2(new_n635), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n697), .A2(KEYINPUT87), .A3(new_n650), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT87), .B1(new_n697), .B2(new_n650), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT29), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n640), .B2(new_n649), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n690), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n671), .B1(new_n703), .B2(G1), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT88), .Z(G364));
  NAND2_X1  g0505(.A1(new_n206), .A2(G13), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT89), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G45), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n668), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n663), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n662), .A2(G330), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n214), .B1(G20), .B2(new_n269), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n209), .A2(new_n259), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT90), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n721), .A2(G355), .B1(new_n427), .B2(new_n666), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n244), .A2(G45), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n666), .A2(new_n259), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n723), .B(new_n724), .C1(G45), .C2(new_n212), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n719), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n206), .A2(G179), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(G190), .A3(G200), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G87), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n300), .A3(G200), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G190), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G159), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT92), .B(KEYINPUT32), .ZN(new_n736));
  OAI221_X1 g0536(.A(new_n730), .B1(new_n368), .B2(new_n731), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n265), .B(new_n737), .C1(new_n735), .C2(new_n736), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n295), .A2(new_n206), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT91), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n740), .A2(new_n732), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G77), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G50), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n300), .A2(G200), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n743), .B1(new_n744), .B2(new_n745), .C1(new_n284), .C2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n740), .A2(new_n300), .A3(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n746), .A2(new_n540), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n750), .A2(new_n218), .B1(new_n430), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT93), .Z(new_n755));
  INV_X1    g0555(.A(new_n750), .ZN(new_n756));
  XNOR2_X1  g0556(.A(KEYINPUT33), .B(G317), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(new_n747), .B2(G322), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT96), .Z(new_n759));
  XNOR2_X1  g0559(.A(KEYINPUT94), .B(G326), .ZN(new_n760));
  INV_X1    g0560(.A(new_n525), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n745), .A2(new_n760), .B1(new_n761), .B2(new_n753), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT95), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n259), .B1(new_n734), .B2(G329), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n766), .B1(new_n767), .B2(new_n731), .C1(new_n443), .C2(new_n728), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n741), .B2(G311), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n764), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n749), .A2(new_n755), .B1(new_n759), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n726), .B1(new_n771), .B2(new_n717), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n661), .B(new_n716), .C1(new_n469), .C2(new_n660), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n713), .B1(new_n710), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT97), .Z(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(G396));
  AND3_X1   g0577(.A1(new_n591), .A2(new_n626), .A3(new_n576), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n626), .B1(new_n591), .B2(new_n576), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n778), .A2(new_n779), .A3(new_n505), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT83), .B1(new_n780), .B2(KEYINPUT26), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(new_n639), .A3(new_n631), .ZN(new_n782));
  INV_X1    g0582(.A(new_n629), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n649), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n364), .A2(new_n649), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n373), .A2(new_n269), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n786), .A2(new_n364), .A3(new_n377), .A4(new_n649), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT98), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n376), .A2(KEYINPUT98), .A3(new_n377), .A4(new_n649), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n378), .A2(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n784), .B(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n690), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n710), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n717), .A2(new_n714), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n709), .B1(new_n261), .B2(new_n797), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n767), .A2(new_n750), .B1(new_n745), .B2(new_n443), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n265), .B1(new_n733), .B2(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n220), .A2(new_n731), .B1(new_n728), .B2(new_n368), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(G97), .C2(new_n752), .ZN(new_n803));
  INV_X1    g0603(.A(G294), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n748), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n799), .B(new_n805), .C1(G116), .C2(new_n741), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G143), .A2(new_n747), .B1(new_n741), .B2(G159), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  INV_X1    g0608(.A(G150), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n745), .C1(new_n809), .C2(new_n750), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT34), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G50), .A2(new_n729), .B1(new_n752), .B2(G58), .ZN(new_n812));
  INV_X1    g0612(.A(new_n731), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G68), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n265), .B1(new_n734), .B2(G132), .ZN(new_n815));
  AND3_X1   g0615(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n806), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n717), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n798), .B1(new_n715), .B2(new_n792), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n796), .A2(new_n819), .ZN(G384));
  INV_X1    g0620(.A(new_n483), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(KEYINPUT35), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(KEYINPUT35), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n822), .A2(G116), .A3(new_n215), .A4(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT36), .Z(new_n825));
  OR3_X1    g0625(.A1(new_n212), .A2(new_n261), .A3(new_n380), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n744), .A2(G68), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT99), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n205), .B(G13), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT104), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n647), .B1(new_n398), .B2(new_n404), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n425), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n405), .A2(new_n646), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n415), .A2(new_n834), .A3(new_n835), .A4(new_n421), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n415), .A2(new_n834), .A3(new_n421), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(KEYINPUT102), .B1(new_n837), .B2(KEYINPUT37), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n832), .A2(KEYINPUT37), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT102), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n839), .A2(new_n840), .A3(new_n415), .A4(new_n421), .ZN(new_n841));
  AOI22_X1  g0641(.A1(KEYINPUT103), .A2(new_n833), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT103), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n425), .A2(new_n843), .A3(new_n832), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT38), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT39), .ZN(new_n846));
  INV_X1    g0646(.A(new_n836), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n391), .A2(new_n272), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n388), .A2(new_n383), .A3(G68), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT16), .B1(new_n851), .B2(new_n382), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n404), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n414), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n646), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n854), .A2(new_n855), .A3(new_n421), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT101), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n856), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n847), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  INV_X1    g0662(.A(new_n855), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n425), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n846), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n831), .B1(new_n845), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n860), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT101), .B1(new_n856), .B2(KEYINPUT37), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n836), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n425), .A2(new_n863), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n861), .A2(new_n865), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT39), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n833), .A2(KEYINPUT103), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n836), .A2(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n837), .A2(KEYINPUT37), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n841), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(new_n844), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n862), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n870), .A2(new_n864), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(KEYINPUT104), .A3(new_n846), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n867), .A2(new_n874), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n346), .A2(new_n649), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT72), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n344), .B(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n329), .B2(new_n332), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n650), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n888), .A2(new_n349), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n333), .A2(new_n889), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT100), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n889), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n346), .A2(new_n350), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT100), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(new_n896), .A3(new_n891), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n782), .A2(new_n783), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n650), .A3(new_n792), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n597), .A2(new_n649), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n871), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n862), .B1(new_n861), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n881), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n903), .A2(new_n906), .B1(new_n596), .B2(new_n647), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n885), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n700), .A2(new_n426), .A3(new_n702), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT105), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT105), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n700), .A2(new_n702), .A3(new_n911), .A4(new_n426), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n603), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n908), .B(new_n913), .Z(new_n914));
  NOR2_X1   g0714(.A1(new_n469), .A2(new_n592), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(new_n691), .A3(new_n650), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n684), .A2(new_n687), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n791), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n893), .A3(new_n897), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n880), .A2(KEYINPUT106), .A3(new_n881), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT106), .B1(new_n880), .B2(new_n881), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n919), .B1(new_n905), .B2(new_n881), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n924), .B1(KEYINPUT40), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n917), .A2(new_n916), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n426), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n928), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(G330), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n914), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n205), .B2(new_n707), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n914), .A2(new_n931), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n830), .B1(new_n933), .B2(new_n934), .ZN(G367));
  NAND2_X1  g0735(.A1(new_n708), .A2(G1), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n703), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n664), .A2(KEYINPUT109), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n651), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n659), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n654), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n649), .A2(new_n490), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n625), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n633), .A2(new_n649), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n942), .A2(new_n943), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT45), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n658), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n664), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT109), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT44), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n658), .B2(new_n947), .ZN(new_n958));
  INV_X1    g0758(.A(new_n947), .ZN(new_n959));
  OAI211_X1 g0759(.A(KEYINPUT44), .B(new_n959), .C1(new_n657), .C2(new_n654), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n940), .B1(new_n956), .B2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n950), .A2(new_n951), .B1(new_n954), .B2(new_n953), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n939), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n655), .A2(new_n656), .A3(new_n651), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n942), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(new_n663), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n938), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n667), .B(KEYINPUT41), .Z(new_n971));
  OAI21_X1  g0771(.A(new_n937), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n657), .A2(new_n947), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT42), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n625), .A2(new_n606), .A3(new_n944), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n649), .B1(new_n975), .B2(new_n505), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n649), .A2(new_n620), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n778), .A2(new_n779), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n695), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT43), .B1(new_n981), .B2(KEYINPUT107), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(KEYINPUT107), .B2(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n953), .A2(new_n947), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n977), .A2(new_n983), .B1(KEYINPUT108), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n974), .B2(new_n976), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n985), .A2(KEYINPUT108), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n979), .A2(new_n716), .A3(new_n980), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n724), .A2(new_n236), .ZN(new_n994));
  INV_X1    g0794(.A(new_n360), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n718), .C1(new_n209), .C2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n710), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT110), .Z(new_n998));
  AOI21_X1  g0798(.A(new_n259), .B1(new_n734), .B2(G317), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n368), .B2(new_n753), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n728), .A2(new_n427), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT46), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(G97), .C2(new_n813), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n741), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n767), .B2(new_n1004), .C1(new_n443), .C2(new_n748), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n800), .A2(new_n745), .B1(new_n750), .B2(new_n761), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G50), .A2(new_n741), .B1(new_n747), .B2(G150), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n752), .A2(G68), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n284), .B2(new_n728), .C1(new_n808), .C2(new_n733), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n259), .B1(new_n731), .B2(new_n261), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1009), .B1(KEYINPUT111), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1007), .B(new_n1011), .C1(KEYINPUT111), .C2(new_n1010), .ZN(new_n1012));
  INV_X1    g0812(.A(G143), .ZN(new_n1013));
  INV_X1    g0813(.A(G159), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n1013), .A2(new_n745), .B1(new_n750), .B2(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1005), .A2(new_n1006), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT47), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n818), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n998), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n972), .A2(new_n992), .B1(new_n993), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(G387));
  INV_X1    g0822(.A(new_n667), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n969), .B2(new_n703), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n703), .B2(new_n969), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n655), .A2(new_n656), .A3(new_n716), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n233), .A2(G45), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n724), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n721), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1027), .A2(new_n1028), .B1(new_n669), .B2(new_n1029), .ZN(new_n1030));
  OR3_X1    g0830(.A1(new_n282), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1031));
  OAI21_X1  g0831(.A(KEYINPUT50), .B1(new_n282), .B2(G50), .ZN(new_n1032));
  AOI21_X1  g0832(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1031), .A2(new_n669), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1030), .A2(new_n1034), .B1(new_n368), .B2(new_n666), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n710), .B1(new_n1035), .B2(new_n719), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1004), .A2(new_n218), .B1(new_n286), .B2(new_n750), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT112), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n745), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(G159), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n747), .A2(G50), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n259), .B1(new_n733), .B2(new_n809), .C1(new_n430), .C2(new_n731), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n753), .A2(new_n995), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G77), .C2(new_n729), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .A4(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n753), .A2(new_n767), .B1(new_n728), .B2(new_n761), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G303), .A2(new_n741), .B1(new_n747), .B2(G317), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1039), .A2(G322), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n800), .C2(new_n750), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n265), .B1(new_n733), .B2(new_n760), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G116), .B2(new_n813), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1045), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1036), .B1(new_n1058), .B2(new_n717), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n969), .A2(new_n936), .B1(new_n1026), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1025), .A2(new_n1060), .ZN(G393));
  NAND3_X1  g0861(.A1(new_n966), .A2(new_n703), .A3(new_n969), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n969), .A2(new_n703), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n963), .A2(new_n1063), .A3(new_n965), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n667), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n937), .B1(new_n963), .B2(new_n965), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT115), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n241), .A2(new_n1028), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n718), .B1(new_n430), .B2(new_n209), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n710), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n756), .A2(G50), .B1(new_n741), .B2(new_n355), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT113), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT113), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n259), .B1(new_n733), .B2(new_n1013), .C1(new_n220), .C2(new_n731), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n753), .A2(new_n261), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(G68), .C2(new_n729), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1039), .A2(G150), .B1(new_n747), .B2(G159), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1039), .A2(G317), .B1(new_n747), .B2(G311), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n756), .A2(G303), .B1(G116), .B2(new_n752), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT114), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(KEYINPUT114), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n259), .B1(new_n734), .B2(G322), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n368), .B2(new_n731), .C1(new_n767), .C2(new_n728), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n741), .B2(G294), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1078), .A2(new_n1080), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1070), .B1(new_n1090), .B2(new_n717), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n959), .A2(new_n716), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1066), .A2(new_n1067), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n965), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n939), .B1(new_n964), .B2(new_n961), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n936), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT115), .B1(new_n1098), .B2(new_n1093), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1065), .B1(new_n1095), .B2(new_n1099), .ZN(G390));
  NAND2_X1  g0900(.A1(new_n910), .A2(new_n912), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n426), .A2(G330), .A3(new_n927), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n688), .A2(KEYINPUT86), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n687), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n683), .A2(new_n685), .A3(KEYINPUT31), .A4(new_n649), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n916), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1106), .A2(G330), .A3(new_n792), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n898), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n918), .A2(new_n893), .A3(new_n897), .A4(G330), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n900), .A2(new_n902), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n690), .A2(new_n792), .A3(new_n893), .A4(new_n897), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n792), .B1(new_n698), .B2(new_n699), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n927), .A2(G330), .A3(new_n792), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n898), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n902), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1101), .A2(new_n604), .A3(new_n1102), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n884), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n901), .B1(new_n784), .B2(new_n792), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n898), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1123), .A2(new_n867), .A3(new_n874), .A4(new_n882), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n898), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n692), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n696), .B1(new_n628), .B2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n634), .A2(KEYINPUT26), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n650), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT87), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n697), .A2(KEYINPUT87), .A3(new_n650), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n791), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1125), .B1(new_n1133), .B2(new_n901), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1134), .B(new_n1121), .C1(new_n922), .C2(new_n923), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1109), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1124), .A2(new_n1135), .A3(new_n1113), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1120), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1124), .A2(new_n1113), .A3(new_n1135), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1109), .B1(new_n1124), .B2(new_n1135), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1119), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1143), .A3(new_n667), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n883), .A2(new_n715), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G107), .A2(new_n756), .B1(new_n1039), .B2(G283), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1076), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n259), .B1(new_n734), .B2(G294), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1148), .A2(new_n730), .A3(new_n814), .A4(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n747), .B2(G116), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1147), .B(new_n1151), .C1(new_n430), .C2(new_n1004), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n741), .A2(new_n1154), .B1(G159), .B2(new_n752), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n808), .B2(new_n750), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT116), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n259), .B1(new_n733), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n728), .A2(new_n809), .ZN(new_n1160));
  XOR2_X1   g0960(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1161));
  XNOR2_X1  g0961(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1159), .B(new_n1162), .C1(G50), .C2(new_n813), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1039), .A2(G128), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n747), .A2(G132), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1152), .B1(new_n1157), .B2(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1167), .A2(new_n717), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n709), .B(new_n1168), .C1(new_n286), .C2(new_n797), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1145), .A2(new_n936), .B1(new_n1146), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1144), .A2(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(new_n921), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT106), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n845), .B2(new_n873), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n880), .A2(KEYINPUT106), .A3(new_n881), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(G330), .B1(new_n925), .B2(KEYINPUT40), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n294), .A2(new_n646), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n307), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n307), .A2(new_n1178), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OR3_X1    g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1182), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1176), .A2(new_n1177), .A3(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n918), .A2(new_n893), .A3(new_n897), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n872), .B2(new_n873), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n672), .B1(new_n1189), .B2(new_n920), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1185), .B1(new_n924), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n908), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1186), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n924), .A2(new_n1190), .A3(new_n1185), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n885), .A4(new_n907), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n936), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1186), .A2(new_n714), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n797), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n710), .B1(G50), .B2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n259), .A2(G41), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n744), .B1(G33), .B2(G41), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT118), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n430), .A2(new_n750), .B1(new_n745), .B2(new_n427), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n731), .A2(new_n284), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT119), .Z(new_n1207));
  OAI211_X1 g1007(.A(new_n1008), .B(new_n1201), .C1(new_n767), .C2(new_n733), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G77), .B2(new_n729), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1207), .B(new_n1209), .C1(new_n1004), .C2(new_n995), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1205), .B(new_n1210), .C1(G107), .C2(new_n747), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1204), .B1(new_n1211), .B2(KEYINPUT58), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n745), .A2(new_n1158), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n747), .A2(G128), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n729), .A2(new_n1154), .B1(new_n752), .B2(G150), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n1004), .C2(new_n808), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1213), .B(new_n1216), .C1(G132), .C2(new_n756), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n813), .A2(G159), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G33), .B(G41), .C1(new_n734), .C2(G124), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1212), .B1(KEYINPUT58), .B2(new_n1211), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1200), .B1(new_n1224), .B2(new_n717), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1198), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT120), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1197), .A2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1141), .A2(new_n1142), .A3(new_n1119), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1101), .A2(new_n604), .A3(new_n1102), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT121), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n913), .A2(KEYINPUT121), .A3(new_n1102), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1196), .B1(new_n1229), .B2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AND4_X1   g1037(.A1(KEYINPUT121), .A2(new_n1101), .A3(new_n604), .A4(new_n1102), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT121), .B1(new_n913), .B2(new_n1102), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1140), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1236), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1023), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1228), .B1(new_n1237), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(G375));
  INV_X1    g1045(.A(new_n1118), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1230), .A2(new_n1246), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n971), .B(KEYINPUT122), .Z(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1119), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n898), .A2(new_n714), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1199), .A2(G68), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT124), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1207), .A2(new_n259), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1252), .A2(new_n1253), .B1(new_n1039), .B2(G132), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n1252), .B2(new_n1253), .C1(new_n750), .C2(new_n1153), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n741), .A2(G150), .B1(G50), .B2(new_n752), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n729), .A2(G159), .B1(new_n734), .B2(G128), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT125), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1256), .B(new_n1258), .C1(new_n808), .C2(new_n748), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n747), .A2(G283), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n741), .A2(G107), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n259), .B(new_n1043), .C1(G77), .C2(new_n813), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n728), .A2(new_n430), .B1(new_n733), .B2(new_n443), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT123), .Z(new_n1264));
  NAND4_X1  g1064(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n427), .A2(new_n750), .B1(new_n745), .B2(new_n804), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1255), .A2(new_n1259), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n709), .B(new_n1251), .C1(new_n1267), .C2(new_n717), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1118), .A2(new_n936), .B1(new_n1250), .B2(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1249), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(G381));
  NOR2_X1   g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  INV_X1    g1072(.A(G384), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(G387), .A2(G390), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G378), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1244), .A4(new_n1270), .ZN(G407));
  NAND2_X1  g1077(.A1(new_n648), .A2(G213), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1244), .A2(new_n1276), .A3(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G407), .A2(G213), .A3(new_n1280), .ZN(G409));
  AND2_X1   g1081(.A1(new_n1197), .A2(new_n1227), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1229), .A2(new_n1234), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1187), .A2(new_n908), .A3(new_n1191), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1193), .A2(new_n1194), .B1(new_n885), .B2(new_n907), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT57), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n667), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT57), .B1(new_n1241), .B2(new_n1196), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1282), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1241), .A2(new_n1196), .A3(new_n1248), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1196), .A2(new_n936), .B1(new_n1198), .B2(new_n1225), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1276), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1247), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1230), .A2(KEYINPUT60), .A3(new_n1246), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n667), .A3(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(G384), .A3(new_n1269), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G384), .B1(new_n1298), .B2(new_n1269), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1294), .A2(new_n1278), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT62), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1279), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n1307), .A3(new_n1302), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1295), .A2(new_n1247), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1297), .A2(new_n667), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1269), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1273), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1279), .A2(G2897), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1312), .A2(new_n1299), .A3(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1312), .B2(new_n1299), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G378), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(G378), .B2(new_n1244), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1316), .B1(new_n1318), .B2(new_n1279), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1304), .A2(new_n1305), .A3(new_n1308), .A4(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n776), .B1(new_n1025), .B2(new_n1060), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1272), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G390), .A2(new_n1322), .ZN(new_n1323));
  OAI221_X1 g1123(.A(new_n1065), .B1(new_n1272), .B2(new_n1321), .C1(new_n1099), .C2(new_n1095), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1323), .A2(new_n1324), .A3(new_n1021), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1021), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1320), .A2(new_n1328), .ZN(new_n1329));
  OAI211_X1 g1129(.A(G2897), .B(new_n1279), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1312), .A2(new_n1299), .A3(new_n1313), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1327), .B(new_n1305), .C1(new_n1306), .C2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1303), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1337), .B1(new_n1303), .B2(new_n1335), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1306), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(new_n1302), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1334), .A2(new_n1336), .A3(new_n1338), .A4(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1329), .A2(new_n1340), .ZN(G405));
  XNOR2_X1  g1141(.A(new_n1244), .B(G378), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(new_n1302), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1328), .ZN(new_n1344));
  OR2_X1    g1144(.A1(new_n1342), .A2(new_n1302), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1342), .A2(new_n1302), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1345), .A2(new_n1327), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1344), .A2(new_n1347), .ZN(G402));
endmodule


