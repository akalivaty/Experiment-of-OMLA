

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n404) );
  XNOR2_X1 U324 ( .A(n405), .B(n404), .ZN(n411) );
  XNOR2_X1 U325 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U326 ( .A(n308), .B(n307), .ZN(n455) );
  NOR2_X1 U327 ( .A1(n530), .A2(n450), .ZN(n559) );
  XNOR2_X1 U328 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U329 ( .A(n454), .B(n453), .ZN(G1349GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT75), .B(KEYINPUT77), .Z(n293) );
  XOR2_X1 U331 ( .A(G85GAT), .B(G92GAT), .Z(n344) );
  XNOR2_X1 U332 ( .A(G176GAT), .B(G204GAT), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n291), .B(G64GAT), .ZN(n415) );
  XNOR2_X1 U334 ( .A(n344), .B(n415), .ZN(n292) );
  XOR2_X1 U335 ( .A(n293), .B(n292), .Z(n299) );
  XOR2_X1 U336 ( .A(G78GAT), .B(G148GAT), .Z(n295) );
  XNOR2_X1 U337 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n333) );
  XOR2_X1 U339 ( .A(n333), .B(KEYINPUT74), .Z(n297) );
  NAND2_X1 U340 ( .A1(G230GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n308) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(G71GAT), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n300), .B(G120GAT), .ZN(n309) );
  XOR2_X1 U345 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n302) );
  XNOR2_X1 U346 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n371) );
  XNOR2_X1 U348 ( .A(n309), .B(n371), .ZN(n306) );
  XOR2_X1 U349 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n304) );
  XNOR2_X1 U350 ( .A(KEYINPUT31), .B(KEYINPUT78), .ZN(n303) );
  XOR2_X1 U351 ( .A(n304), .B(n303), .Z(n305) );
  XOR2_X1 U352 ( .A(KEYINPUT41), .B(n455), .Z(n547) );
  XOR2_X1 U353 ( .A(n547), .B(KEYINPUT108), .Z(n533) );
  XOR2_X1 U354 ( .A(G43GAT), .B(G134GAT), .Z(n354) );
  XOR2_X1 U355 ( .A(G15GAT), .B(G127GAT), .Z(n376) );
  XNOR2_X1 U356 ( .A(n354), .B(n376), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n315) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n311), .B(KEYINPUT85), .ZN(n435) );
  XOR2_X1 U360 ( .A(n435), .B(KEYINPUT87), .Z(n313) );
  NAND2_X1 U361 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U363 ( .A(n315), .B(n314), .Z(n324) );
  XNOR2_X1 U364 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n316), .B(KEYINPUT18), .ZN(n317) );
  XOR2_X1 U366 ( .A(n317), .B(KEYINPUT19), .Z(n319) );
  XNOR2_X1 U367 ( .A(G169GAT), .B(G190GAT), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n424) );
  XOR2_X1 U369 ( .A(G176GAT), .B(KEYINPUT20), .Z(n321) );
  XNOR2_X1 U370 ( .A(KEYINPUT86), .B(KEYINPUT88), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n424), .B(n322), .ZN(n323) );
  XOR2_X1 U373 ( .A(n324), .B(n323), .Z(n497) );
  INV_X1 U374 ( .A(n497), .ZN(n530) );
  XOR2_X1 U375 ( .A(KEYINPUT90), .B(G218GAT), .Z(n326) );
  XNOR2_X1 U376 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U378 ( .A(G197GAT), .B(n327), .Z(n416) );
  XOR2_X1 U379 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n329) );
  NAND2_X1 U380 ( .A1(G228GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U382 ( .A(n330), .B(KEYINPUT22), .Z(n335) );
  XOR2_X1 U383 ( .A(KEYINPUT91), .B(KEYINPUT3), .Z(n332) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n434) );
  XNOR2_X1 U386 ( .A(n434), .B(n333), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U388 ( .A(G204GAT), .B(KEYINPUT24), .Z(n337) );
  XNOR2_X1 U389 ( .A(KEYINPUT23), .B(KEYINPUT93), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(n339), .B(n338), .Z(n341) );
  XOR2_X1 U392 ( .A(G50GAT), .B(G162GAT), .Z(n343) );
  XOR2_X1 U393 ( .A(G22GAT), .B(G155GAT), .Z(n370) );
  XNOR2_X1 U394 ( .A(n343), .B(n370), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n416), .B(n342), .ZN(n464) );
  XOR2_X1 U397 ( .A(n344), .B(n343), .Z(n346) );
  NAND2_X1 U398 ( .A1(G232GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U400 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n348) );
  XNOR2_X1 U401 ( .A(G190GAT), .B(G106GAT), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U403 ( .A(n350), .B(n349), .Z(n356) );
  XOR2_X1 U404 ( .A(KEYINPUT9), .B(KEYINPUT80), .Z(n352) );
  XNOR2_X1 U405 ( .A(G218GAT), .B(KEYINPUT79), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U409 ( .A(n357), .B(G99GAT), .Z(n361) );
  XOR2_X1 U410 ( .A(G29GAT), .B(KEYINPUT8), .Z(n359) );
  XNOR2_X1 U411 ( .A(KEYINPUT7), .B(KEYINPUT70), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n387) );
  XNOR2_X1 U413 ( .A(n387), .B(G36GAT), .ZN(n360) );
  XOR2_X1 U414 ( .A(n361), .B(n360), .Z(n554) );
  INV_X1 U415 ( .A(n554), .ZN(n558) );
  XOR2_X1 U416 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n363) );
  XNOR2_X1 U417 ( .A(G8GAT), .B(G64GAT), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U419 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n365) );
  XNOR2_X1 U420 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n380) );
  XOR2_X1 U423 ( .A(G78GAT), .B(G211GAT), .Z(n369) );
  XNOR2_X1 U424 ( .A(G183GAT), .B(G71GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n375) );
  XOR2_X1 U426 ( .A(n371), .B(n370), .Z(n373) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U429 ( .A(n375), .B(n374), .Z(n378) );
  XOR2_X1 U430 ( .A(G1GAT), .B(KEYINPUT71), .Z(n386) );
  XNOR2_X1 U431 ( .A(n386), .B(n376), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U433 ( .A(n380), .B(n379), .Z(n551) );
  INV_X1 U434 ( .A(n551), .ZN(n574) );
  XOR2_X1 U435 ( .A(G113GAT), .B(G197GAT), .Z(n382) );
  XNOR2_X1 U436 ( .A(G141GAT), .B(G22GAT), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U438 ( .A(n383), .B(G43GAT), .Z(n385) );
  XOR2_X1 U439 ( .A(G36GAT), .B(G8GAT), .Z(n420) );
  XNOR2_X1 U440 ( .A(n420), .B(G50GAT), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n391) );
  XOR2_X1 U442 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U443 ( .A1(G229GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U445 ( .A(n391), .B(n390), .Z(n399) );
  XOR2_X1 U446 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n393) );
  XNOR2_X1 U447 ( .A(G169GAT), .B(G15GAT), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U449 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n395) );
  XNOR2_X1 U450 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U453 ( .A(n399), .B(n398), .Z(n566) );
  INV_X1 U454 ( .A(n566), .ZN(n544) );
  NOR2_X1 U455 ( .A1(n544), .A2(n547), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n400), .B(KEYINPUT46), .ZN(n401) );
  NOR2_X1 U457 ( .A1(n574), .A2(n401), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n402), .B(KEYINPUT113), .ZN(n403) );
  NOR2_X1 U459 ( .A1(n558), .A2(n403), .ZN(n405) );
  XNOR2_X1 U460 ( .A(KEYINPUT36), .B(n554), .ZN(n581) );
  NOR2_X1 U461 ( .A1(n581), .A2(n551), .ZN(n406) );
  XNOR2_X1 U462 ( .A(KEYINPUT45), .B(n406), .ZN(n407) );
  NAND2_X1 U463 ( .A1(n407), .A2(n455), .ZN(n408) );
  XNOR2_X1 U464 ( .A(KEYINPUT115), .B(n408), .ZN(n409) );
  NAND2_X1 U465 ( .A1(n409), .A2(n544), .ZN(n410) );
  NAND2_X1 U466 ( .A1(n411), .A2(n410), .ZN(n414) );
  XOR2_X1 U467 ( .A(KEYINPUT64), .B(KEYINPUT116), .Z(n412) );
  XNOR2_X1 U468 ( .A(KEYINPUT48), .B(n412), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n526) );
  XOR2_X1 U470 ( .A(KEYINPUT99), .B(n415), .Z(n418) );
  XNOR2_X1 U471 ( .A(n416), .B(G92GAT), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U473 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U476 ( .A(n424), .B(n423), .Z(n494) );
  INV_X1 U477 ( .A(n494), .ZN(n516) );
  NOR2_X1 U478 ( .A1(n526), .A2(n516), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n425), .B(KEYINPUT54), .ZN(n448) );
  XOR2_X1 U480 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n427) );
  XNOR2_X1 U481 ( .A(G57GAT), .B(KEYINPUT98), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n439) );
  XOR2_X1 U483 ( .A(KEYINPUT4), .B(G120GAT), .Z(n429) );
  XNOR2_X1 U484 ( .A(G1GAT), .B(G127GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U486 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n431) );
  XNOR2_X1 U487 ( .A(KEYINPUT1), .B(KEYINPUT95), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n447) );
  NAND2_X1 U493 ( .A1(G225GAT), .A2(G233GAT), .ZN(n445) );
  XOR2_X1 U494 ( .A(G155GAT), .B(G162GAT), .Z(n441) );
  XNOR2_X1 U495 ( .A(G134GAT), .B(G148GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U497 ( .A(G29GAT), .B(G85GAT), .Z(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U500 ( .A(n447), .B(n446), .Z(n490) );
  INV_X1 U501 ( .A(n490), .ZN(n514) );
  NAND2_X1 U502 ( .A1(n448), .A2(n514), .ZN(n564) );
  NOR2_X1 U503 ( .A1(n464), .A2(n564), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  NAND2_X1 U505 ( .A1(n533), .A2(n559), .ZN(n454) );
  XOR2_X1 U506 ( .A(G176GAT), .B(KEYINPUT56), .Z(n452) );
  XNOR2_X1 U507 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n451) );
  INV_X1 U508 ( .A(n455), .ZN(n571) );
  NOR2_X1 U509 ( .A1(n544), .A2(n571), .ZN(n488) );
  XOR2_X1 U510 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n457) );
  NAND2_X1 U511 ( .A1(n574), .A2(n554), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(n473) );
  XNOR2_X1 U513 ( .A(KEYINPUT27), .B(n494), .ZN(n467) );
  NAND2_X1 U514 ( .A1(n490), .A2(n467), .ZN(n525) );
  XOR2_X1 U515 ( .A(KEYINPUT89), .B(n497), .Z(n458) );
  NOR2_X1 U516 ( .A1(n525), .A2(n458), .ZN(n460) );
  XNOR2_X1 U517 ( .A(KEYINPUT28), .B(KEYINPUT65), .ZN(n459) );
  XOR2_X1 U518 ( .A(n459), .B(n464), .Z(n501) );
  INV_X1 U519 ( .A(n501), .ZN(n528) );
  NAND2_X1 U520 ( .A1(n460), .A2(n528), .ZN(n472) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n463) );
  NOR2_X1 U522 ( .A1(n530), .A2(n516), .ZN(n461) );
  NOR2_X1 U523 ( .A1(n464), .A2(n461), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n463), .B(n462), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n464), .A2(n530), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n465), .B(KEYINPUT100), .ZN(n466) );
  XOR2_X1 U527 ( .A(KEYINPUT26), .B(n466), .Z(n562) );
  NAND2_X1 U528 ( .A1(n562), .A2(n467), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n514), .A2(n470), .ZN(n471) );
  NAND2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n484) );
  AND2_X1 U532 ( .A1(n473), .A2(n484), .ZN(n503) );
  NAND2_X1 U533 ( .A1(n488), .A2(n503), .ZN(n482) );
  NOR2_X1 U534 ( .A1(n514), .A2(n482), .ZN(n475) );
  XNOR2_X1 U535 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n476), .Z(G1324GAT) );
  NOR2_X1 U538 ( .A1(n516), .A2(n482), .ZN(n478) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n478), .B(n477), .ZN(G1325GAT) );
  NOR2_X1 U541 ( .A1(n530), .A2(n482), .ZN(n480) );
  XNOR2_X1 U542 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U544 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  NOR2_X1 U545 ( .A1(n528), .A2(n482), .ZN(n483) );
  XOR2_X1 U546 ( .A(G22GAT), .B(n483), .Z(G1327GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT39), .B(KEYINPUT106), .Z(n492) );
  NAND2_X1 U548 ( .A1(n551), .A2(n484), .ZN(n485) );
  NOR2_X1 U549 ( .A1(n581), .A2(n485), .ZN(n487) );
  XNOR2_X1 U550 ( .A(KEYINPUT105), .B(KEYINPUT37), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(n513) );
  NAND2_X1 U552 ( .A1(n488), .A2(n513), .ZN(n489) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(n489), .Z(n500) );
  NAND2_X1 U554 ( .A1(n490), .A2(n500), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  XOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT107), .Z(n496) );
  NAND2_X1 U558 ( .A1(n494), .A2(n500), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n497), .A2(n500), .ZN(n498) );
  XNOR2_X1 U561 ( .A(KEYINPUT40), .B(n498), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NAND2_X1 U563 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n502), .ZN(G1331GAT) );
  AND2_X1 U565 ( .A1(n544), .A2(n533), .ZN(n512) );
  NAND2_X1 U566 ( .A1(n512), .A2(n503), .ZN(n509) );
  NOR2_X1 U567 ( .A1(n514), .A2(n509), .ZN(n504) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n504), .Z(n505) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n516), .A2(n509), .ZN(n506) );
  XOR2_X1 U571 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U572 ( .A1(n530), .A2(n509), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n528), .A2(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n514), .A2(n522), .ZN(n515) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n515), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n522), .ZN(n517) );
  XOR2_X1 U582 ( .A(KEYINPUT110), .B(n517), .Z(n518) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(n518), .ZN(G1337GAT) );
  NOR2_X1 U584 ( .A1(n530), .A2(n522), .ZN(n519) );
  XOR2_X1 U585 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n521) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n524) );
  NOR2_X1 U589 ( .A1(n528), .A2(n522), .ZN(n523) );
  XOR2_X1 U590 ( .A(n524), .B(n523), .Z(G1339GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT117), .B(n527), .Z(n543) );
  NAND2_X1 U593 ( .A1(n543), .A2(n528), .ZN(n529) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n566), .A2(n538), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT118), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U599 ( .A1(n538), .A2(n533), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NAND2_X1 U601 ( .A1(n538), .A2(n574), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(KEYINPUT50), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n558), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT119), .Z(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n562), .A2(n543), .ZN(n553) );
  NOR2_X1 U610 ( .A1(n544), .A2(n553), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT121), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  NOR2_X1 U613 ( .A1(n547), .A2(n553), .ZN(n549) );
  XNOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n553), .ZN(n552) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U620 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  NAND2_X1 U621 ( .A1(n559), .A2(n566), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n559), .A2(n574), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT58), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(n561), .ZN(G1351GAT) );
  INV_X1 U628 ( .A(n562), .ZN(n563) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT123), .B(n565), .ZN(n580) );
  INV_X1 U631 ( .A(n580), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n566), .A2(n575), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U638 ( .A1(n575), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT125), .Z(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n579) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(n583), .B(n582), .Z(G1355GAT) );
endmodule

