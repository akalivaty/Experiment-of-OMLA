

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801;

  XNOR2_X1 U380 ( .A(n430), .B(KEYINPUT0), .ZN(n385) );
  XNOR2_X1 U381 ( .A(n476), .B(n440), .ZN(n782) );
  NOR2_X1 U382 ( .A1(G953), .A2(G237), .ZN(n529) );
  AND2_X1 U383 ( .A1(n409), .A2(G224), .ZN(n402) );
  INV_X1 U384 ( .A(G902), .ZN(n531) );
  XNOR2_X1 U385 ( .A(n507), .B(n506), .ZN(n784) );
  BUF_X1 U386 ( .A(n396), .Z(n770) );
  XNOR2_X2 U387 ( .A(n522), .B(n521), .ZN(n614) );
  NOR2_X1 U388 ( .A1(n622), .A2(n720), .ZN(n623) );
  XNOR2_X2 U389 ( .A(n511), .B(n540), .ZN(n502) );
  INV_X1 U390 ( .A(G953), .ZN(n534) );
  OR2_X1 U391 ( .A1(n577), .A2(n573), .ZN(n717) );
  NAND2_X1 U392 ( .A1(n667), .A2(n358), .ZN(n672) );
  BUF_X1 U393 ( .A(n751), .Z(n378) );
  NOR2_X1 U394 ( .A1(n364), .A2(n363), .ZN(n362) );
  AND2_X1 U395 ( .A1(n448), .A2(n450), .ZN(n653) );
  NOR2_X1 U396 ( .A1(n617), .A2(n690), .ZN(n365) );
  NAND2_X1 U397 ( .A1(n739), .A2(n374), .ZN(n587) );
  XNOR2_X1 U398 ( .A(n447), .B(KEYINPUT41), .ZN(n729) );
  NOR2_X1 U399 ( .A1(n734), .A2(n733), .ZN(n447) );
  XNOR2_X1 U400 ( .A(n377), .B(n639), .ZN(n731) );
  NAND2_X1 U401 ( .A1(n577), .A2(n556), .ZN(n622) );
  BUF_X1 U402 ( .A(n577), .Z(n578) );
  XNOR2_X1 U403 ( .A(n370), .B(n371), .ZN(n577) );
  XNOR2_X1 U404 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U405 ( .A(n465), .B(n432), .ZN(n771) );
  AND2_X1 U406 ( .A1(n546), .A2(G210), .ZN(n358) );
  AND2_X1 U407 ( .A1(n546), .A2(G472), .ZN(n359) );
  XNOR2_X1 U408 ( .A(n389), .B(n459), .ZN(n514) );
  AND2_X1 U409 ( .A1(n438), .A2(n437), .ZN(n400) );
  XNOR2_X1 U410 ( .A(n458), .B(n457), .ZN(n389) );
  NAND2_X1 U411 ( .A1(n446), .A2(n445), .ZN(n444) );
  NAND2_X1 U412 ( .A1(n475), .A2(KEYINPUT3), .ZN(n446) );
  XNOR2_X1 U413 ( .A(n442), .B(n441), .ZN(n440) );
  INV_X1 U414 ( .A(G224), .ZN(n439) );
  XNOR2_X1 U415 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n442) );
  NAND2_X1 U416 ( .A1(G953), .A2(KEYINPUT18), .ZN(n437) );
  INV_X1 U417 ( .A(KEYINPUT18), .ZN(n409) );
  INV_X1 U418 ( .A(KEYINPUT3), .ZN(n474) );
  NAND2_X1 U419 ( .A1(n667), .A2(n359), .ZN(n679) );
  NAND2_X1 U420 ( .A1(n361), .A2(n360), .ZN(n367) );
  AND2_X1 U421 ( .A1(n598), .A2(KEYINPUT44), .ZN(n360) );
  NAND2_X1 U422 ( .A1(n597), .A2(KEYINPUT90), .ZN(n361) );
  NAND2_X1 U423 ( .A1(n366), .A2(n362), .ZN(n621) );
  AND2_X1 U424 ( .A1(n689), .A2(n619), .ZN(n363) );
  NAND2_X1 U425 ( .A1(n618), .A2(n365), .ZN(n364) );
  NAND2_X1 U426 ( .A1(n368), .A2(n367), .ZN(n366) );
  NAND2_X1 U427 ( .A1(n369), .A2(n596), .ZN(n368) );
  NAND2_X1 U428 ( .A1(n593), .A2(n689), .ZN(n369) );
  XNOR2_X2 U429 ( .A(n592), .B(n591), .ZN(n689) );
  XOR2_X1 U430 ( .A(n470), .B(n390), .Z(n370) );
  NOR2_X1 U431 ( .A1(n771), .A2(G902), .ZN(n371) );
  XNOR2_X2 U432 ( .A(n372), .B(n373), .ZN(n560) );
  NOR2_X1 U433 ( .A1(n762), .A2(G902), .ZN(n372) );
  XOR2_X1 U434 ( .A(KEYINPUT71), .B(G469), .Z(n373) );
  INV_X1 U435 ( .A(n613), .ZN(n374) );
  BUF_X1 U436 ( .A(n799), .Z(n375) );
  NAND2_X1 U437 ( .A1(n665), .A2(n664), .ZN(n376) );
  NAND2_X1 U438 ( .A1(n665), .A2(n664), .ZN(n667) );
  XNOR2_X1 U439 ( .A(n552), .B(n551), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n552), .B(n551), .ZN(n566) );
  NAND2_X1 U441 ( .A1(n717), .A2(KEYINPUT109), .ZN(n416) );
  XNOR2_X1 U442 ( .A(n463), .B(G137), .ZN(n497) );
  INV_X1 U443 ( .A(KEYINPUT70), .ZN(n463) );
  OR2_X1 U444 ( .A1(n426), .A2(n419), .ZN(n422) );
  NOR2_X1 U445 ( .A1(n420), .A2(n424), .ZN(n423) );
  NOR2_X1 U446 ( .A1(n632), .A2(n425), .ZN(n424) );
  NOR2_X1 U447 ( .A1(n636), .A2(n421), .ZN(n420) );
  NAND2_X1 U448 ( .A1(KEYINPUT47), .A2(KEYINPUT85), .ZN(n421) );
  INV_X1 U449 ( .A(G953), .ZN(n410) );
  NOR2_X1 U450 ( .A1(n453), .A2(n451), .ZN(n450) );
  NAND2_X1 U451 ( .A1(n474), .A2(G119), .ZN(n445) );
  XNOR2_X1 U452 ( .A(n434), .B(G125), .ZN(n536) );
  INV_X1 U453 ( .A(G146), .ZN(n434) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n734) );
  INV_X1 U455 ( .A(KEYINPUT113), .ZN(n383) );
  INV_X1 U456 ( .A(KEYINPUT30), .ZN(n408) );
  XNOR2_X1 U457 ( .A(n382), .B(KEYINPUT108), .ZN(n733) );
  XNOR2_X1 U458 ( .A(G128), .B(G119), .ZN(n460) );
  XNOR2_X1 U459 ( .A(n387), .B(n497), .ZN(n386) );
  XNOR2_X1 U460 ( .A(n536), .B(n433), .ZN(n790) );
  XNOR2_X1 U461 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n433) );
  XNOR2_X1 U462 ( .A(n527), .B(n381), .ZN(n429) );
  XNOR2_X1 U463 ( .A(G143), .B(G113), .ZN(n525) );
  NAND2_X1 U464 ( .A1(n684), .A2(n531), .ZN(n533) );
  XNOR2_X1 U465 ( .A(n520), .B(n519), .ZN(n768) );
  XNOR2_X1 U466 ( .A(n513), .B(n512), .ZN(n520) );
  AND2_X1 U467 ( .A1(n673), .A2(G953), .ZN(n774) );
  INV_X1 U468 ( .A(KEYINPUT85), .ZN(n425) );
  XNOR2_X1 U469 ( .A(KEYINPUT97), .B(KEYINPUT15), .ZN(n466) );
  NAND2_X1 U470 ( .A1(n415), .A2(n414), .ZN(n413) );
  NOR2_X1 U471 ( .A1(n717), .A2(KEYINPUT109), .ZN(n414) );
  XOR2_X1 U472 ( .A(KEYINPUT104), .B(KEYINPUT76), .Z(n478) );
  XNOR2_X1 U473 ( .A(G137), .B(G131), .ZN(n480) );
  XNOR2_X1 U474 ( .A(n502), .B(n501), .ZN(n411) );
  XNOR2_X1 U475 ( .A(KEYINPUT80), .B(KEYINPUT17), .ZN(n539) );
  XNOR2_X1 U476 ( .A(n399), .B(n535), .ZN(n418) );
  NAND2_X1 U477 ( .A1(n400), .A2(n401), .ZN(n399) );
  XNOR2_X1 U478 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n620) );
  NOR2_X1 U479 ( .A1(G902), .A2(G237), .ZN(n488) );
  INV_X1 U480 ( .A(KEYINPUT48), .ZN(n652) );
  INV_X1 U481 ( .A(G110), .ZN(n506) );
  INV_X1 U482 ( .A(G122), .ZN(n441) );
  XNOR2_X1 U483 ( .A(G116), .B(G107), .ZN(n515) );
  INV_X1 U484 ( .A(KEYINPUT105), .ZN(n512) );
  NOR2_X1 U485 ( .A1(n622), .A2(n602), .ZN(n558) );
  NAND2_X1 U486 ( .A1(n602), .A2(n578), .ZN(n431) );
  AND2_X1 U487 ( .A1(n510), .A2(n627), .ZN(n642) );
  XNOR2_X1 U488 ( .A(n490), .B(n408), .ZN(n407) );
  XOR2_X1 U489 ( .A(KEYINPUT62), .B(n677), .Z(n678) );
  XNOR2_X1 U490 ( .A(n388), .B(n386), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n428), .B(n528), .ZN(n684) );
  XNOR2_X1 U492 ( .A(n530), .B(n429), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n404), .B(n403), .ZN(n769) );
  INV_X1 U494 ( .A(n768), .ZN(n403) );
  NAND2_X1 U495 ( .A1(n770), .A2(G478), .ZN(n404) );
  AND2_X1 U496 ( .A1(n415), .A2(n412), .ZN(n379) );
  AND2_X1 U497 ( .A1(n417), .A2(n416), .ZN(n380) );
  AND2_X1 U498 ( .A1(G214), .A2(n529), .ZN(n381) );
  NAND2_X1 U499 ( .A1(n572), .A2(n614), .ZN(n382) );
  NAND2_X1 U500 ( .A1(n731), .A2(n730), .ZN(n384) );
  INV_X1 U501 ( .A(n385), .ZN(n613) );
  NAND2_X1 U502 ( .A1(n574), .A2(n385), .ZN(n576) );
  XNOR2_X1 U503 ( .A(n464), .B(KEYINPUT101), .ZN(n387) );
  NAND2_X1 U504 ( .A1(n514), .A2(G221), .ZN(n388) );
  INV_X1 U505 ( .A(KEYINPUT102), .ZN(n390) );
  BUF_X1 U506 ( .A(n646), .Z(n391) );
  XNOR2_X1 U507 ( .A(n670), .B(n669), .ZN(n671) );
  INV_X1 U508 ( .A(n739), .ZN(n392) );
  INV_X1 U509 ( .A(n392), .ZN(n393) );
  INV_X1 U510 ( .A(n597), .ZN(n394) );
  BUF_X2 U511 ( .A(n716), .Z(n395) );
  AND2_X2 U512 ( .A1(n376), .A2(n546), .ZN(n396) );
  BUF_X1 U513 ( .A(n603), .Z(n397) );
  NAND2_X1 U514 ( .A1(n603), .A2(n436), .ZN(n435) );
  XNOR2_X1 U515 ( .A(n395), .B(KEYINPUT96), .ZN(n650) );
  NAND2_X1 U516 ( .A1(n799), .A2(n583), .ZN(n398) );
  NAND2_X1 U517 ( .A1(n799), .A2(n583), .ZN(n599) );
  BUF_X1 U518 ( .A(n661), .Z(n775) );
  XNOR2_X1 U519 ( .A(n621), .B(n620), .ZN(n661) );
  XNOR2_X2 U520 ( .A(KEYINPUT67), .B(G101), .ZN(n535) );
  NAND2_X1 U521 ( .A1(n402), .A2(n410), .ZN(n401) );
  NAND2_X1 U522 ( .A1(n406), .A2(n405), .ZN(n665) );
  NOR2_X1 U523 ( .A1(n680), .A2(n774), .ZN(n682) );
  NOR2_X1 U524 ( .A1(n674), .A2(n774), .ZN(n676) );
  NOR2_X1 U525 ( .A1(n687), .A2(n774), .ZN(n688) );
  INV_X1 U526 ( .A(n659), .ZN(n405) );
  INV_X1 U527 ( .A(n660), .ZN(n406) );
  NOR2_X1 U528 ( .A1(n800), .A2(n801), .ZN(n449) );
  XNOR2_X1 U529 ( .A(n645), .B(KEYINPUT40), .ZN(n800) );
  NAND2_X1 U530 ( .A1(n407), .A2(n554), .ZN(n496) );
  NAND2_X1 U531 ( .A1(n439), .A2(KEYINPUT18), .ZN(n438) );
  XNOR2_X1 U532 ( .A(n411), .B(n509), .ZN(n762) );
  XNOR2_X1 U533 ( .A(n411), .B(n790), .ZN(n793) );
  INV_X1 U534 ( .A(n717), .ZN(n412) );
  NAND2_X1 U535 ( .A1(n380), .A2(n413), .ZN(n456) );
  INV_X1 U536 ( .A(n716), .ZN(n415) );
  NAND2_X1 U537 ( .A1(n716), .A2(KEYINPUT109), .ZN(n417) );
  NAND2_X1 U538 ( .A1(n379), .A2(n610), .ZN(n723) );
  XNOR2_X1 U539 ( .A(n418), .B(n536), .ZN(n538) );
  NAND2_X1 U540 ( .A1(n632), .A2(n425), .ZN(n419) );
  NOR2_X1 U541 ( .A1(n636), .A2(n427), .ZN(n426) );
  NAND2_X1 U542 ( .A1(n423), .A2(n422), .ZN(n633) );
  INV_X1 U543 ( .A(n636), .ZN(n735) );
  INV_X1 U544 ( .A(KEYINPUT47), .ZN(n427) );
  NOR2_X2 U545 ( .A1(n629), .A2(n571), .ZN(n430) );
  XNOR2_X2 U546 ( .A(n646), .B(KEYINPUT19), .ZN(n629) );
  XNOR2_X2 U547 ( .A(n567), .B(KEYINPUT93), .ZN(n646) );
  NOR2_X1 U548 ( .A1(n650), .A2(n431), .ZN(n582) );
  XNOR2_X2 U549 ( .A(n435), .B(KEYINPUT32), .ZN(n799) );
  XNOR2_X1 U550 ( .A(n582), .B(KEYINPUT82), .ZN(n436) );
  XNOR2_X2 U551 ( .A(n576), .B(n575), .ZN(n603) );
  XNOR2_X2 U552 ( .A(n444), .B(n443), .ZN(n476) );
  XNOR2_X2 U553 ( .A(G113), .B(G116), .ZN(n443) );
  XNOR2_X1 U554 ( .A(n449), .B(KEYINPUT46), .ZN(n448) );
  XNOR2_X1 U555 ( .A(n452), .B(KEYINPUT86), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n633), .A2(n634), .ZN(n452) );
  OR2_X1 U557 ( .A1(n709), .A2(n638), .ZN(n453) );
  XNOR2_X2 U558 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n540) );
  XNOR2_X2 U559 ( .A(n454), .B(G143), .ZN(n542) );
  XNOR2_X2 U560 ( .A(G128), .B(KEYINPUT84), .ZN(n454) );
  XNOR2_X2 U561 ( .A(n455), .B(n585), .ZN(n739) );
  NAND2_X1 U562 ( .A1(n456), .A2(n581), .ZN(n455) );
  BUF_X1 U563 ( .A(n762), .Z(n763) );
  AND2_X2 U564 ( .A1(n661), .A2(n791), .ZN(n751) );
  INV_X1 U565 ( .A(KEYINPUT5), .ZN(n479) );
  XNOR2_X1 U566 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U567 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U568 ( .A(KEYINPUT87), .ZN(n457) );
  INV_X1 U569 ( .A(KEYINPUT38), .ZN(n639) );
  BUF_X1 U570 ( .A(n668), .Z(n670) );
  NAND2_X1 U571 ( .A1(G234), .A2(n534), .ZN(n458) );
  XOR2_X1 U572 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n459) );
  XOR2_X1 U573 ( .A(G140), .B(G110), .Z(n461) );
  XNOR2_X1 U574 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U575 ( .A(n790), .B(n462), .ZN(n465) );
  XOR2_X1 U576 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n464) );
  XOR2_X1 U577 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n469) );
  XNOR2_X1 U578 ( .A(n466), .B(n531), .ZN(n666) );
  NAND2_X1 U579 ( .A1(G234), .A2(n666), .ZN(n467) );
  XNOR2_X1 U580 ( .A(KEYINPUT20), .B(n467), .ZN(n471) );
  NAND2_X1 U581 ( .A1(n471), .A2(G217), .ZN(n468) );
  XNOR2_X1 U582 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U583 ( .A1(n471), .A2(G221), .ZN(n472) );
  XNOR2_X1 U584 ( .A(KEYINPUT21), .B(n472), .ZN(n714) );
  INV_X1 U585 ( .A(KEYINPUT103), .ZN(n473) );
  XNOR2_X1 U586 ( .A(n714), .B(n473), .ZN(n573) );
  XNOR2_X1 U587 ( .A(n535), .B(G146), .ZN(n505) );
  INV_X1 U588 ( .A(G119), .ZN(n475) );
  XNOR2_X1 U589 ( .A(n505), .B(n476), .ZN(n484) );
  NAND2_X1 U590 ( .A1(n529), .A2(G210), .ZN(n477) );
  XNOR2_X1 U591 ( .A(n478), .B(n477), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X2 U593 ( .A(n542), .B(G134), .ZN(n511) );
  XNOR2_X1 U594 ( .A(n485), .B(n502), .ZN(n677) );
  NAND2_X1 U595 ( .A1(n677), .A2(n531), .ZN(n486) );
  XNOR2_X2 U596 ( .A(n486), .B(G472), .ZN(n610) );
  INV_X1 U597 ( .A(KEYINPUT75), .ZN(n487) );
  XNOR2_X1 U598 ( .A(n488), .B(n487), .ZN(n548) );
  INV_X1 U599 ( .A(G214), .ZN(n489) );
  OR2_X1 U600 ( .A1(n548), .A2(n489), .ZN(n730) );
  NAND2_X1 U601 ( .A1(n610), .A2(n730), .ZN(n490) );
  NAND2_X1 U602 ( .A1(G234), .A2(G237), .ZN(n491) );
  XNOR2_X1 U603 ( .A(n491), .B(KEYINPUT14), .ZN(n494) );
  NAND2_X1 U604 ( .A1(n494), .A2(G902), .ZN(n492) );
  XNOR2_X1 U605 ( .A(n492), .B(KEYINPUT99), .ZN(n568) );
  NAND2_X1 U606 ( .A1(G953), .A2(n568), .ZN(n493) );
  NOR2_X1 U607 ( .A1(G900), .A2(n493), .ZN(n495) );
  AND2_X1 U608 ( .A1(G952), .A2(n494), .ZN(n744) );
  AND2_X1 U609 ( .A1(n744), .A2(n534), .ZN(n569) );
  OR2_X1 U610 ( .A1(n495), .A2(n569), .ZN(n554) );
  NOR2_X1 U611 ( .A1(n717), .A2(n496), .ZN(n510) );
  XNOR2_X1 U612 ( .A(n497), .B(KEYINPUT100), .ZN(n500) );
  INV_X1 U613 ( .A(G140), .ZN(n498) );
  XNOR2_X1 U614 ( .A(n498), .B(G131), .ZN(n523) );
  INV_X1 U615 ( .A(n523), .ZN(n499) );
  XNOR2_X1 U616 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U617 ( .A1(n534), .A2(G227), .ZN(n503) );
  XNOR2_X1 U618 ( .A(n503), .B(KEYINPUT79), .ZN(n504) );
  XNOR2_X1 U619 ( .A(n505), .B(n504), .ZN(n508) );
  XNOR2_X2 U620 ( .A(G104), .B(G107), .ZN(n507) );
  XNOR2_X1 U621 ( .A(n784), .B(KEYINPUT72), .ZN(n537) );
  XNOR2_X1 U622 ( .A(n508), .B(n537), .ZN(n509) );
  INV_X1 U623 ( .A(n560), .ZN(n627) );
  XNOR2_X1 U624 ( .A(n511), .B(KEYINPUT9), .ZN(n513) );
  NAND2_X1 U625 ( .A1(G217), .A2(n514), .ZN(n518) );
  XOR2_X1 U626 ( .A(KEYINPUT7), .B(G122), .Z(n516) );
  XNOR2_X1 U627 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U628 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U629 ( .A1(n768), .A2(n531), .ZN(n522) );
  XOR2_X1 U630 ( .A(KEYINPUT106), .B(G478), .Z(n521) );
  XNOR2_X1 U631 ( .A(n523), .B(KEYINPUT12), .ZN(n524) );
  XNOR2_X1 U632 ( .A(n524), .B(KEYINPUT11), .ZN(n528) );
  XOR2_X1 U633 ( .A(G122), .B(G104), .Z(n526) );
  XNOR2_X1 U634 ( .A(n526), .B(n525), .ZN(n527) );
  INV_X1 U635 ( .A(n790), .ZN(n530) );
  XOR2_X1 U636 ( .A(KEYINPUT13), .B(G475), .Z(n532) );
  XNOR2_X1 U637 ( .A(n533), .B(n532), .ZN(n615) );
  INV_X1 U638 ( .A(n615), .ZN(n572) );
  OR2_X1 U639 ( .A1(n614), .A2(n572), .ZN(n588) );
  XNOR2_X1 U640 ( .A(n538), .B(n537), .ZN(n545) );
  XNOR2_X1 U641 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U642 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U643 ( .A(n543), .B(n782), .ZN(n544) );
  XNOR2_X1 U644 ( .A(n545), .B(n544), .ZN(n668) );
  INV_X1 U645 ( .A(n666), .ZN(n546) );
  OR2_X2 U646 ( .A1(n668), .A2(n546), .ZN(n552) );
  INV_X1 U647 ( .A(G210), .ZN(n547) );
  OR2_X1 U648 ( .A1(n548), .A2(n547), .ZN(n550) );
  INV_X1 U649 ( .A(KEYINPUT98), .ZN(n549) );
  XNOR2_X1 U650 ( .A(n550), .B(n549), .ZN(n551) );
  INV_X1 U651 ( .A(n377), .ZN(n563) );
  NOR2_X1 U652 ( .A1(n588), .A2(n563), .ZN(n553) );
  NAND2_X1 U653 ( .A1(n642), .A2(n553), .ZN(n632) );
  XNOR2_X1 U654 ( .A(n632), .B(G143), .ZN(G45) );
  XNOR2_X1 U655 ( .A(G140), .B(KEYINPUT118), .ZN(n565) );
  NAND2_X1 U656 ( .A1(n615), .A2(n614), .ZN(n644) );
  XNOR2_X1 U657 ( .A(KEYINPUT110), .B(n644), .ZN(n703) );
  INV_X1 U658 ( .A(n554), .ZN(n555) );
  NOR2_X1 U659 ( .A1(n555), .A2(n714), .ZN(n556) );
  INV_X1 U660 ( .A(KEYINPUT6), .ZN(n557) );
  XNOR2_X1 U661 ( .A(n610), .B(n557), .ZN(n581) );
  INV_X1 U662 ( .A(n581), .ZN(n602) );
  XNOR2_X1 U663 ( .A(n558), .B(KEYINPUT111), .ZN(n559) );
  NOR2_X1 U664 ( .A1(n703), .A2(n559), .ZN(n647) );
  AND2_X1 U665 ( .A1(n647), .A2(n730), .ZN(n561) );
  XNOR2_X2 U666 ( .A(n560), .B(KEYINPUT1), .ZN(n716) );
  NAND2_X1 U667 ( .A1(n561), .A2(n395), .ZN(n562) );
  XNOR2_X1 U668 ( .A(n562), .B(KEYINPUT43), .ZN(n564) );
  AND2_X1 U669 ( .A1(n564), .A2(n563), .ZN(n656) );
  XOR2_X1 U670 ( .A(n565), .B(n656), .Z(G42) );
  NAND2_X1 U671 ( .A1(n566), .A2(n730), .ZN(n567) );
  NOR2_X1 U672 ( .A1(G898), .A2(n534), .ZN(n787) );
  AND2_X1 U673 ( .A1(n568), .A2(n787), .ZN(n570) );
  NOR2_X1 U674 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U675 ( .A1(n733), .A2(n573), .ZN(n574) );
  XNOR2_X1 U676 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n575) );
  INV_X1 U677 ( .A(n610), .ZN(n720) );
  NAND2_X1 U678 ( .A1(n578), .A2(n720), .ZN(n579) );
  INV_X1 U679 ( .A(n395), .ZN(n605) );
  NOR2_X1 U680 ( .A1(n579), .A2(n605), .ZN(n580) );
  NAND2_X1 U681 ( .A1(n397), .A2(n580), .ZN(n583) );
  XNOR2_X1 U682 ( .A(n583), .B(G110), .ZN(G12) );
  XNOR2_X1 U683 ( .A(n599), .B(KEYINPUT91), .ZN(n593) );
  INV_X1 U684 ( .A(KEYINPUT95), .ZN(n584) );
  XNOR2_X1 U685 ( .A(n584), .B(KEYINPUT33), .ZN(n585) );
  INV_X1 U686 ( .A(KEYINPUT34), .ZN(n586) );
  XNOR2_X1 U687 ( .A(n587), .B(n586), .ZN(n590) );
  INV_X1 U688 ( .A(n588), .ZN(n589) );
  NAND2_X1 U689 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U690 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n591) );
  INV_X1 U691 ( .A(KEYINPUT44), .ZN(n594) );
  NAND2_X1 U692 ( .A1(n594), .A2(KEYINPUT66), .ZN(n595) );
  INV_X1 U693 ( .A(KEYINPUT90), .ZN(n619) );
  NOR2_X1 U694 ( .A1(n595), .A2(n619), .ZN(n596) );
  INV_X1 U695 ( .A(n689), .ZN(n597) );
  NAND2_X1 U696 ( .A1(n398), .A2(KEYINPUT66), .ZN(n598) );
  INV_X1 U697 ( .A(n398), .ZN(n601) );
  INV_X1 U698 ( .A(KEYINPUT66), .ZN(n600) );
  NAND2_X1 U699 ( .A1(n601), .A2(n600), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U701 ( .A(n604), .B(KEYINPUT89), .ZN(n607) );
  NOR2_X1 U702 ( .A1(n578), .A2(n605), .ZN(n606) );
  AND2_X1 U703 ( .A1(n607), .A2(n606), .ZN(n690) );
  OR2_X1 U704 ( .A1(n613), .A2(n723), .ZN(n609) );
  INV_X1 U705 ( .A(KEYINPUT31), .ZN(n608) );
  XNOR2_X2 U706 ( .A(n609), .B(n608), .ZN(n705) );
  NOR2_X1 U707 ( .A1(n717), .A2(n610), .ZN(n611) );
  NAND2_X1 U708 ( .A1(n611), .A2(n627), .ZN(n612) );
  OR2_X1 U709 ( .A1(n613), .A2(n612), .ZN(n693) );
  NAND2_X1 U710 ( .A1(n705), .A2(n693), .ZN(n616) );
  NOR2_X1 U711 ( .A1(n615), .A2(n614), .ZN(n697) );
  XNOR2_X1 U712 ( .A(KEYINPUT107), .B(n697), .ZN(n654) );
  NAND2_X1 U713 ( .A1(n644), .A2(n654), .ZN(n636) );
  AND2_X1 U714 ( .A1(n616), .A2(n636), .ZN(n617) );
  XNOR2_X1 U715 ( .A(KEYINPUT28), .B(KEYINPUT112), .ZN(n624) );
  NAND2_X1 U716 ( .A1(n624), .A2(n623), .ZN(n626) );
  OR2_X1 U717 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U718 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U719 ( .A1(n628), .A2(n627), .ZN(n640) );
  NOR2_X1 U720 ( .A1(n640), .A2(n629), .ZN(n631) );
  INV_X1 U721 ( .A(KEYINPUT83), .ZN(n630) );
  XNOR2_X1 U722 ( .A(n631), .B(n630), .ZN(n635) );
  OR2_X1 U723 ( .A1(n635), .A2(n427), .ZN(n634) );
  NAND2_X1 U724 ( .A1(n635), .A2(n636), .ZN(n637) );
  NOR2_X1 U725 ( .A1(n637), .A2(KEYINPUT47), .ZN(n638) );
  NOR2_X1 U726 ( .A1(n729), .A2(n640), .ZN(n641) );
  XNOR2_X1 U727 ( .A(KEYINPUT42), .B(n641), .ZN(n801) );
  AND2_X1 U728 ( .A1(n642), .A2(n731), .ZN(n643) );
  XNOR2_X1 U729 ( .A(n643), .B(KEYINPUT39), .ZN(n655) );
  NOR2_X1 U730 ( .A1(n655), .A2(n644), .ZN(n645) );
  NAND2_X1 U731 ( .A1(n647), .A2(n391), .ZN(n649) );
  XNOR2_X1 U732 ( .A(KEYINPUT92), .B(KEYINPUT36), .ZN(n648) );
  XNOR2_X1 U733 ( .A(n649), .B(n648), .ZN(n651) );
  NOR2_X1 U734 ( .A1(n651), .A2(n650), .ZN(n709) );
  XNOR2_X1 U735 ( .A(n653), .B(n652), .ZN(n658) );
  NOR2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n712) );
  OR2_X1 U737 ( .A1(n712), .A2(n656), .ZN(n657) );
  NOR2_X1 U738 ( .A1(n658), .A2(n657), .ZN(n791) );
  XNOR2_X1 U739 ( .A(n751), .B(KEYINPUT2), .ZN(n660) );
  AND2_X1 U740 ( .A1(n751), .A2(KEYINPUT77), .ZN(n659) );
  INV_X1 U741 ( .A(n775), .ZN(n754) );
  INV_X1 U742 ( .A(n791), .ZN(n747) );
  NAND2_X1 U743 ( .A1(n747), .A2(KEYINPUT77), .ZN(n662) );
  NOR2_X1 U744 ( .A1(n754), .A2(n662), .ZN(n663) );
  INV_X1 U745 ( .A(n663), .ZN(n664) );
  XOR2_X1 U746 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n669) );
  XNOR2_X1 U747 ( .A(n672), .B(n671), .ZN(n674) );
  INV_X1 U748 ( .A(G952), .ZN(n673) );
  XNOR2_X1 U749 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n675) );
  XNOR2_X1 U750 ( .A(n676), .B(n675), .ZN(G51) );
  XNOR2_X1 U751 ( .A(n679), .B(n678), .ZN(n680) );
  XOR2_X1 U752 ( .A(KEYINPUT94), .B(KEYINPUT63), .Z(n681) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(G57) );
  NAND2_X1 U754 ( .A1(n396), .A2(G475), .ZN(n686) );
  XOR2_X1 U755 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n683) );
  XNOR2_X1 U756 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U757 ( .A(n688), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U758 ( .A(n394), .B(G122), .ZN(G24) );
  XOR2_X1 U759 ( .A(G101), .B(n690), .Z(G3) );
  NOR2_X1 U760 ( .A1(n703), .A2(n693), .ZN(n691) );
  XOR2_X1 U761 ( .A(KEYINPUT114), .B(n691), .Z(n692) );
  XNOR2_X1 U762 ( .A(G104), .B(n692), .ZN(G6) );
  INV_X1 U763 ( .A(n697), .ZN(n706) );
  NOR2_X1 U764 ( .A1(n706), .A2(n693), .ZN(n695) );
  XNOR2_X1 U765 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n694) );
  XNOR2_X1 U766 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U767 ( .A(G107), .B(n696), .ZN(G9) );
  XOR2_X1 U768 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n699) );
  NAND2_X1 U769 ( .A1(n635), .A2(n697), .ZN(n698) );
  XNOR2_X1 U770 ( .A(n699), .B(n698), .ZN(n700) );
  XOR2_X1 U771 ( .A(G128), .B(n700), .Z(G30) );
  INV_X1 U772 ( .A(n635), .ZN(n701) );
  NOR2_X1 U773 ( .A1(n703), .A2(n701), .ZN(n702) );
  XOR2_X1 U774 ( .A(G146), .B(n702), .Z(G48) );
  NOR2_X1 U775 ( .A1(n703), .A2(n705), .ZN(n704) );
  XOR2_X1 U776 ( .A(G113), .B(n704), .Z(G15) );
  NOR2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U778 ( .A(KEYINPUT116), .B(n707), .Z(n708) );
  XNOR2_X1 U779 ( .A(G116), .B(n708), .ZN(G18) );
  XOR2_X1 U780 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n711) );
  XNOR2_X1 U781 ( .A(G125), .B(n709), .ZN(n710) );
  XNOR2_X1 U782 ( .A(n711), .B(n710), .ZN(G27) );
  XOR2_X1 U783 ( .A(G134), .B(n712), .Z(G36) );
  NOR2_X1 U784 ( .A1(n729), .A2(n392), .ZN(n713) );
  NOR2_X1 U785 ( .A1(n713), .A2(G953), .ZN(n746) );
  NAND2_X1 U786 ( .A1(n714), .A2(n578), .ZN(n715) );
  XNOR2_X1 U787 ( .A(n715), .B(KEYINPUT49), .ZN(n722) );
  NAND2_X1 U788 ( .A1(n717), .A2(n395), .ZN(n718) );
  XNOR2_X1 U789 ( .A(n718), .B(KEYINPUT50), .ZN(n719) );
  NAND2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U791 ( .A1(n722), .A2(n721), .ZN(n725) );
  INV_X1 U792 ( .A(n723), .ZN(n724) );
  NOR2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U794 ( .A(n726), .B(KEYINPUT51), .ZN(n727) );
  XNOR2_X1 U795 ( .A(KEYINPUT119), .B(n727), .ZN(n728) );
  NOR2_X1 U796 ( .A1(n729), .A2(n728), .ZN(n741) );
  NOR2_X1 U797 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U798 ( .A1(n733), .A2(n732), .ZN(n737) );
  NOR2_X1 U799 ( .A1(n735), .A2(n734), .ZN(n736) );
  OR2_X1 U800 ( .A1(n737), .A2(n736), .ZN(n738) );
  AND2_X1 U801 ( .A1(n393), .A2(n738), .ZN(n740) );
  NOR2_X1 U802 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U803 ( .A(KEYINPUT52), .B(n742), .Z(n743) );
  NAND2_X1 U804 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U805 ( .A1(n746), .A2(n745), .ZN(n758) );
  NOR2_X1 U806 ( .A1(n747), .A2(KEYINPUT88), .ZN(n748) );
  NOR2_X1 U807 ( .A1(n378), .A2(n748), .ZN(n749) );
  NOR2_X1 U808 ( .A1(n749), .A2(KEYINPUT2), .ZN(n753) );
  NAND2_X1 U809 ( .A1(KEYINPUT2), .A2(KEYINPUT88), .ZN(n750) );
  NOR2_X1 U810 ( .A1(n378), .A2(n750), .ZN(n752) );
  NOR2_X1 U811 ( .A1(n753), .A2(n752), .ZN(n756) );
  NOR2_X1 U812 ( .A1(n754), .A2(KEYINPUT88), .ZN(n755) );
  NOR2_X1 U813 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U814 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U815 ( .A(KEYINPUT53), .B(n759), .ZN(G75) );
  NAND2_X1 U816 ( .A1(n770), .A2(G469), .ZN(n766) );
  XOR2_X1 U817 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n761) );
  XNOR2_X1 U818 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n760) );
  XNOR2_X1 U819 ( .A(n761), .B(n760), .ZN(n764) );
  XOR2_X1 U820 ( .A(n764), .B(n763), .Z(n765) );
  XNOR2_X1 U821 ( .A(n766), .B(n765), .ZN(n767) );
  NOR2_X1 U822 ( .A1(n774), .A2(n767), .ZN(G54) );
  NOR2_X1 U823 ( .A1(n774), .A2(n769), .ZN(G63) );
  NAND2_X1 U824 ( .A1(n770), .A2(G217), .ZN(n772) );
  XNOR2_X1 U825 ( .A(n772), .B(n771), .ZN(n773) );
  NOR2_X1 U826 ( .A1(n774), .A2(n773), .ZN(G66) );
  NAND2_X1 U827 ( .A1(n775), .A2(n534), .ZN(n781) );
  XOR2_X1 U828 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n777) );
  NAND2_X1 U829 ( .A1(G224), .A2(G953), .ZN(n776) );
  XNOR2_X1 U830 ( .A(n777), .B(n776), .ZN(n778) );
  XNOR2_X1 U831 ( .A(KEYINPUT124), .B(n778), .ZN(n779) );
  NAND2_X1 U832 ( .A1(n779), .A2(G898), .ZN(n780) );
  NAND2_X1 U833 ( .A1(n781), .A2(n780), .ZN(n789) );
  XOR2_X1 U834 ( .A(n782), .B(KEYINPUT126), .Z(n783) );
  XNOR2_X1 U835 ( .A(n784), .B(n783), .ZN(n785) );
  XNOR2_X1 U836 ( .A(n785), .B(G101), .ZN(n786) );
  NOR2_X1 U837 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U838 ( .A(n789), .B(n788), .ZN(G69) );
  XNOR2_X1 U839 ( .A(n791), .B(n793), .ZN(n792) );
  NAND2_X1 U840 ( .A1(n792), .A2(n534), .ZN(n798) );
  XNOR2_X1 U841 ( .A(n793), .B(G227), .ZN(n794) );
  XNOR2_X1 U842 ( .A(n794), .B(KEYINPUT127), .ZN(n795) );
  NAND2_X1 U843 ( .A1(n795), .A2(G900), .ZN(n796) );
  NAND2_X1 U844 ( .A1(n796), .A2(G953), .ZN(n797) );
  NAND2_X1 U845 ( .A1(n798), .A2(n797), .ZN(G72) );
  XNOR2_X1 U846 ( .A(n375), .B(G119), .ZN(G21) );
  XOR2_X1 U847 ( .A(G131), .B(n800), .Z(G33) );
  XOR2_X1 U848 ( .A(G137), .B(n801), .Z(G39) );
endmodule

