

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(n547), .A2(n546), .ZN(G160) );
  BUF_X1 U550 ( .A(n558), .Z(n559) );
  NOR2_X1 U551 ( .A1(G2084), .A2(n733), .ZN(n766) );
  INV_X1 U552 ( .A(n937), .ZN(n775) );
  INV_X1 U553 ( .A(KEYINPUT101), .ZN(n772) );
  XNOR2_X1 U554 ( .A(n773), .B(n772), .ZN(n785) );
  NOR2_X1 U555 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X2 U556 ( .A1(G2105), .A2(n518), .ZN(n858) );
  NOR2_X1 U557 ( .A1(G651), .A2(n648), .ZN(n641) );
  NOR2_X1 U558 ( .A1(n524), .A2(n523), .ZN(G164) );
  NAND2_X1 U559 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  XNOR2_X2 U560 ( .A(n514), .B(KEYINPUT65), .ZN(n862) );
  NAND2_X1 U561 ( .A1(G114), .A2(n862), .ZN(n515) );
  XNOR2_X1 U562 ( .A(n515), .B(KEYINPUT87), .ZN(n524) );
  XNOR2_X1 U563 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n517) );
  NOR2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XNOR2_X1 U565 ( .A(n517), .B(n516), .ZN(n558) );
  NAND2_X1 U566 ( .A1(n558), .A2(G138), .ZN(n522) );
  INV_X1 U567 ( .A(G2104), .ZN(n518) );
  NAND2_X1 U568 ( .A1(G102), .A2(n858), .ZN(n520) );
  AND2_X1 U569 ( .A1(n518), .A2(G2105), .ZN(n861) );
  NAND2_X1 U570 ( .A1(G126), .A2(n861), .ZN(n519) );
  AND2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U573 ( .A(KEYINPUT0), .B(G543), .Z(n648) );
  INV_X1 U574 ( .A(G651), .ZN(n530) );
  NOR2_X1 U575 ( .A1(n648), .A2(n530), .ZN(n635) );
  NAND2_X1 U576 ( .A1(n635), .A2(G76), .ZN(n525) );
  XNOR2_X1 U577 ( .A(KEYINPUT72), .B(n525), .ZN(n528) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n632) );
  NAND2_X1 U579 ( .A1(n632), .A2(G89), .ZN(n526) );
  XNOR2_X1 U580 ( .A(KEYINPUT4), .B(n526), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U582 ( .A(n529), .B(KEYINPUT5), .ZN(n537) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(KEYINPUT73), .ZN(n535) );
  NOR2_X1 U584 ( .A1(G543), .A2(n530), .ZN(n531) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n531), .Z(n647) );
  NAND2_X1 U586 ( .A1(G63), .A2(n647), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G51), .A2(n641), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n535), .B(n534), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U591 ( .A(KEYINPUT7), .B(n538), .ZN(G168) );
  XOR2_X1 U592 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U593 ( .A1(n862), .A2(G113), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n539), .B(KEYINPUT66), .ZN(n547) );
  XOR2_X1 U595 ( .A(KEYINPUT64), .B(KEYINPUT23), .Z(n541) );
  NAND2_X1 U596 ( .A1(G101), .A2(n858), .ZN(n540) );
  XNOR2_X1 U597 ( .A(n541), .B(n540), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G125), .A2(n861), .ZN(n543) );
  NAND2_X1 U599 ( .A1(G137), .A2(n558), .ZN(n542) );
  AND2_X1 U600 ( .A1(n543), .A2(n542), .ZN(n544) );
  AND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U602 ( .A1(G85), .A2(n632), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G60), .A2(n647), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U605 ( .A1(G72), .A2(n635), .ZN(n551) );
  NAND2_X1 U606 ( .A1(G47), .A2(n641), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n552) );
  OR2_X1 U608 ( .A1(n553), .A2(n552), .ZN(G290) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U610 ( .A1(G123), .A2(n861), .ZN(n554) );
  XNOR2_X1 U611 ( .A(n554), .B(KEYINPUT18), .ZN(n557) );
  NAND2_X1 U612 ( .A1(G99), .A2(n858), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n555), .B(KEYINPUT76), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n563) );
  NAND2_X1 U615 ( .A1(G135), .A2(n559), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G111), .A2(n862), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U618 ( .A1(n563), .A2(n562), .ZN(n992) );
  XNOR2_X1 U619 ( .A(n992), .B(G2096), .ZN(n564) );
  XNOR2_X1 U620 ( .A(n564), .B(KEYINPUT77), .ZN(n565) );
  OR2_X1 U621 ( .A1(G2100), .A2(n565), .ZN(G156) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  INV_X1 U624 ( .A(G82), .ZN(G220) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n568) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n566) );
  XOR2_X1 U627 ( .A(n566), .B(KEYINPUT10), .Z(n817) );
  NAND2_X1 U628 ( .A1(G567), .A2(n817), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n568), .B(n567), .ZN(G234) );
  NAND2_X1 U630 ( .A1(n632), .A2(G81), .ZN(n569) );
  XNOR2_X1 U631 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G68), .A2(n635), .ZN(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U634 ( .A(n572), .B(KEYINPUT13), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G43), .A2(n641), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n647), .A2(G56), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n575), .Z(n576) );
  NOR2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n931) );
  INV_X1 U640 ( .A(n931), .ZN(n881) );
  XNOR2_X1 U641 ( .A(G860), .B(KEYINPUT71), .ZN(n605) );
  OR2_X1 U642 ( .A1(n881), .A2(n605), .ZN(G153) );
  NAND2_X1 U643 ( .A1(G90), .A2(n632), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G77), .A2(n635), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(KEYINPUT9), .B(n580), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G64), .A2(n647), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G52), .A2(n641), .ZN(n581) );
  AND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U652 ( .A1(G79), .A2(n635), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G54), .A2(n641), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U655 ( .A1(G92), .A2(n632), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G66), .A2(n647), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U659 ( .A(n591), .B(KEYINPUT15), .Z(n928) );
  INV_X1 U660 ( .A(n928), .ZN(n738) );
  INV_X1 U661 ( .A(G868), .ZN(n660) );
  NAND2_X1 U662 ( .A1(n738), .A2(n660), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G65), .A2(n647), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G53), .A2(n641), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U667 ( .A(KEYINPUT69), .B(n596), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G91), .A2(n632), .ZN(n598) );
  NAND2_X1 U669 ( .A1(G78), .A2(n635), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U671 ( .A(KEYINPUT68), .B(n599), .Z(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(G299) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT74), .ZN(n604) );
  NOR2_X1 U675 ( .A1(n660), .A2(G286), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n606), .A2(n928), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G559), .A2(n660), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n928), .A2(n608), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n609), .B(KEYINPUT75), .ZN(n611) );
  NOR2_X1 U683 ( .A1(n881), .A2(G868), .ZN(n610) );
  NOR2_X1 U684 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G559), .A2(n928), .ZN(n612) );
  XOR2_X1 U686 ( .A(n612), .B(n931), .Z(n656) );
  NOR2_X1 U687 ( .A1(G860), .A2(n656), .ZN(n621) );
  NAND2_X1 U688 ( .A1(G93), .A2(n632), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G80), .A2(n635), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G67), .A2(n647), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G55), .A2(n641), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U694 ( .A(KEYINPUT79), .B(n617), .Z(n618) );
  NOR2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n659) );
  XNOR2_X1 U696 ( .A(n659), .B(KEYINPUT78), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n621), .B(n620), .ZN(G145) );
  NAND2_X1 U698 ( .A1(n632), .A2(G88), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(KEYINPUT84), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G75), .A2(n635), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U702 ( .A(n625), .B(KEYINPUT85), .ZN(n627) );
  NAND2_X1 U703 ( .A1(G50), .A2(n641), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G62), .A2(n647), .ZN(n628) );
  XNOR2_X1 U706 ( .A(KEYINPUT83), .B(n628), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n630), .A2(n629), .ZN(G166) );
  INV_X1 U708 ( .A(G166), .ZN(G303) );
  NAND2_X1 U709 ( .A1(G48), .A2(n641), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n631), .B(KEYINPUT82), .ZN(n640) );
  NAND2_X1 U711 ( .A1(G86), .A2(n632), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G61), .A2(n647), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n635), .A2(G73), .ZN(n636) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U718 ( .A1(G49), .A2(n641), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n642), .B(KEYINPUT80), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n643) );
  XOR2_X1 U721 ( .A(KEYINPUT81), .B(n643), .Z(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(G288) );
  XOR2_X1 U726 ( .A(G303), .B(n659), .Z(n655) );
  XNOR2_X1 U727 ( .A(KEYINPUT19), .B(G299), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n651), .B(G290), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n652), .B(G305), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n653), .B(G288), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n655), .B(n654), .ZN(n882) );
  XOR2_X1 U732 ( .A(n656), .B(n882), .Z(n657) );
  XNOR2_X1 U733 ( .A(KEYINPUT86), .B(n657), .ZN(n658) );
  NOR2_X1 U734 ( .A1(n660), .A2(n658), .ZN(n662) );
  AND2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U736 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U745 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U746 ( .A1(G96), .A2(n669), .ZN(n821) );
  NAND2_X1 U747 ( .A1(n821), .A2(G2106), .ZN(n673) );
  NAND2_X1 U748 ( .A1(G120), .A2(G69), .ZN(n670) );
  NOR2_X1 U749 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U750 ( .A1(G108), .A2(n671), .ZN(n822) );
  NAND2_X1 U751 ( .A1(n822), .A2(G567), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n823) );
  NAND2_X1 U753 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U754 ( .A1(n823), .A2(n674), .ZN(n820) );
  NAND2_X1 U755 ( .A1(n820), .A2(G36), .ZN(G176) );
  INV_X1 U756 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U757 ( .A(G1986), .B(G290), .ZN(n935) );
  NOR2_X1 U758 ( .A1(G164), .A2(G1384), .ZN(n705) );
  NAND2_X1 U759 ( .A1(G160), .A2(G40), .ZN(n675) );
  NOR2_X1 U760 ( .A1(n705), .A2(n675), .ZN(n811) );
  NAND2_X1 U761 ( .A1(n935), .A2(n811), .ZN(n798) );
  XNOR2_X1 U762 ( .A(G2067), .B(KEYINPUT37), .ZN(n799) );
  NAND2_X1 U763 ( .A1(n861), .A2(G128), .ZN(n676) );
  XOR2_X1 U764 ( .A(KEYINPUT89), .B(n676), .Z(n678) );
  NAND2_X1 U765 ( .A1(n862), .A2(G116), .ZN(n677) );
  NAND2_X1 U766 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U767 ( .A(n679), .B(KEYINPUT35), .ZN(n685) );
  NAND2_X1 U768 ( .A1(n858), .A2(G104), .ZN(n680) );
  XNOR2_X1 U769 ( .A(n680), .B(KEYINPUT88), .ZN(n682) );
  NAND2_X1 U770 ( .A1(G140), .A2(n559), .ZN(n681) );
  NAND2_X1 U771 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U772 ( .A(KEYINPUT34), .B(n683), .Z(n684) );
  NAND2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U774 ( .A(n686), .B(KEYINPUT36), .Z(n877) );
  NOR2_X1 U775 ( .A1(n799), .A2(n877), .ZN(n991) );
  NAND2_X1 U776 ( .A1(n811), .A2(n991), .ZN(n806) );
  XOR2_X1 U777 ( .A(KEYINPUT90), .B(G1991), .Z(n909) );
  NAND2_X1 U778 ( .A1(G95), .A2(n858), .ZN(n688) );
  NAND2_X1 U779 ( .A1(G131), .A2(n559), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U781 ( .A1(G119), .A2(n861), .ZN(n690) );
  NAND2_X1 U782 ( .A1(G107), .A2(n862), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n873) );
  NOR2_X1 U785 ( .A1(n909), .A2(n873), .ZN(n701) );
  NAND2_X1 U786 ( .A1(G129), .A2(n861), .ZN(n694) );
  NAND2_X1 U787 ( .A1(G117), .A2(n862), .ZN(n693) );
  NAND2_X1 U788 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n858), .A2(G105), .ZN(n695) );
  XOR2_X1 U790 ( .A(KEYINPUT38), .B(n695), .Z(n696) );
  NOR2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n559), .A2(G141), .ZN(n698) );
  NAND2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n857) );
  AND2_X1 U794 ( .A1(n857), .A2(G1996), .ZN(n700) );
  NOR2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n988) );
  XNOR2_X1 U796 ( .A(KEYINPUT91), .B(n811), .ZN(n702) );
  NOR2_X1 U797 ( .A1(n988), .A2(n702), .ZN(n803) );
  INV_X1 U798 ( .A(n803), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n806), .A2(n703), .ZN(n796) );
  NOR2_X1 U800 ( .A1(G1976), .A2(G288), .ZN(n925) );
  NOR2_X1 U801 ( .A1(G1971), .A2(G303), .ZN(n936) );
  NOR2_X1 U802 ( .A1(n925), .A2(n936), .ZN(n774) );
  INV_X1 U803 ( .A(KEYINPUT93), .ZN(n707) );
  AND2_X1 U804 ( .A1(G160), .A2(G40), .ZN(n704) );
  NAND2_X1 U805 ( .A1(n705), .A2(n704), .ZN(n733) );
  NAND2_X1 U806 ( .A1(G8), .A2(n733), .ZN(n790) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n790), .ZN(n706) );
  XNOR2_X1 U808 ( .A(n707), .B(n706), .ZN(n765) );
  INV_X1 U809 ( .A(KEYINPUT92), .ZN(n708) );
  XNOR2_X1 U810 ( .A(n708), .B(n766), .ZN(n709) );
  NAND2_X1 U811 ( .A1(n709), .A2(G8), .ZN(n710) );
  NOR2_X1 U812 ( .A1(n765), .A2(n710), .ZN(n711) );
  XOR2_X1 U813 ( .A(KEYINPUT30), .B(n711), .Z(n712) );
  NOR2_X1 U814 ( .A1(G168), .A2(n712), .ZN(n717) );
  INV_X1 U815 ( .A(n733), .ZN(n724) );
  NOR2_X1 U816 ( .A1(n724), .A2(G1961), .ZN(n713) );
  XOR2_X1 U817 ( .A(KEYINPUT94), .B(n713), .Z(n715) );
  XNOR2_X1 U818 ( .A(G2078), .B(KEYINPUT25), .ZN(n903) );
  NAND2_X1 U819 ( .A1(n724), .A2(n903), .ZN(n714) );
  NAND2_X1 U820 ( .A1(n715), .A2(n714), .ZN(n750) );
  NOR2_X1 U821 ( .A1(G171), .A2(n750), .ZN(n716) );
  NOR2_X1 U822 ( .A1(n717), .A2(n716), .ZN(n719) );
  XOR2_X1 U823 ( .A(KEYINPUT31), .B(KEYINPUT98), .Z(n718) );
  XNOR2_X1 U824 ( .A(n719), .B(n718), .ZN(n754) );
  NAND2_X1 U825 ( .A1(G1348), .A2(n733), .ZN(n721) );
  NAND2_X1 U826 ( .A1(n724), .A2(G2067), .ZN(n720) );
  NAND2_X1 U827 ( .A1(n721), .A2(n720), .ZN(n739) );
  NAND2_X1 U828 ( .A1(n739), .A2(n738), .ZN(n732) );
  XNOR2_X1 U829 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n725) );
  OR2_X1 U830 ( .A1(n725), .A2(G1996), .ZN(n722) );
  NAND2_X1 U831 ( .A1(n931), .A2(n722), .ZN(n730) );
  INV_X1 U832 ( .A(G1341), .ZN(n932) );
  NAND2_X1 U833 ( .A1(n932), .A2(n725), .ZN(n723) );
  NAND2_X1 U834 ( .A1(n723), .A2(n733), .ZN(n728) );
  AND2_X1 U835 ( .A1(n724), .A2(G1996), .ZN(n726) );
  NAND2_X1 U836 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U837 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U838 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U839 ( .A1(n732), .A2(n731), .ZN(n743) );
  INV_X1 U840 ( .A(G2072), .ZN(n982) );
  NOR2_X1 U841 ( .A1(n733), .A2(n982), .ZN(n735) );
  XOR2_X1 U842 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n734) );
  XNOR2_X1 U843 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U844 ( .A1(n733), .A2(G1956), .ZN(n736) );
  NAND2_X1 U845 ( .A1(n737), .A2(n736), .ZN(n745) );
  NOR2_X1 U846 ( .A1(G299), .A2(n745), .ZN(n741) );
  NOR2_X1 U847 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U848 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U849 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U850 ( .A(KEYINPUT97), .B(n744), .ZN(n748) );
  NAND2_X1 U851 ( .A1(G299), .A2(n745), .ZN(n746) );
  XOR2_X1 U852 ( .A(KEYINPUT28), .B(n746), .Z(n747) );
  NOR2_X1 U853 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U854 ( .A(n749), .B(KEYINPUT29), .ZN(n752) );
  NAND2_X1 U855 ( .A1(G171), .A2(n750), .ZN(n751) );
  NAND2_X1 U856 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U857 ( .A1(n754), .A2(n753), .ZN(n763) );
  NAND2_X1 U858 ( .A1(n763), .A2(G286), .ZN(n759) );
  NOR2_X1 U859 ( .A1(G1971), .A2(n790), .ZN(n756) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n733), .ZN(n755) );
  NOR2_X1 U861 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U862 ( .A1(n757), .A2(G303), .ZN(n758) );
  NAND2_X1 U863 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U864 ( .A(n760), .B(KEYINPUT100), .ZN(n761) );
  NAND2_X1 U865 ( .A1(n761), .A2(G8), .ZN(n762) );
  XNOR2_X1 U866 ( .A(n762), .B(KEYINPUT32), .ZN(n771) );
  XNOR2_X1 U867 ( .A(KEYINPUT99), .B(n763), .ZN(n764) );
  NOR2_X1 U868 ( .A1(n765), .A2(n764), .ZN(n769) );
  XNOR2_X1 U869 ( .A(n766), .B(KEYINPUT92), .ZN(n767) );
  NAND2_X1 U870 ( .A1(G8), .A2(n767), .ZN(n768) );
  NAND2_X1 U871 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U872 ( .A1(n771), .A2(n770), .ZN(n773) );
  NAND2_X1 U873 ( .A1(n774), .A2(n785), .ZN(n777) );
  NAND2_X1 U874 ( .A1(G1976), .A2(G288), .ZN(n937) );
  NOR2_X1 U875 ( .A1(n790), .A2(n775), .ZN(n776) );
  AND2_X1 U876 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U877 ( .A1(KEYINPUT33), .A2(n778), .ZN(n781) );
  NAND2_X1 U878 ( .A1(n925), .A2(KEYINPUT33), .ZN(n779) );
  NOR2_X1 U879 ( .A1(n779), .A2(n790), .ZN(n780) );
  XOR2_X1 U880 ( .A(G1981), .B(G305), .Z(n948) );
  NAND2_X1 U881 ( .A1(n782), .A2(n948), .ZN(n794) );
  NOR2_X1 U882 ( .A1(G2090), .A2(G303), .ZN(n783) );
  XNOR2_X1 U883 ( .A(n783), .B(KEYINPUT102), .ZN(n784) );
  NAND2_X1 U884 ( .A1(n784), .A2(G8), .ZN(n786) );
  NAND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n787) );
  AND2_X1 U886 ( .A1(n787), .A2(n790), .ZN(n792) );
  NOR2_X1 U887 ( .A1(G1981), .A2(G305), .ZN(n788) );
  XOR2_X1 U888 ( .A(n788), .B(KEYINPUT24), .Z(n789) );
  NOR2_X1 U889 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U890 ( .A1(n792), .A2(n791), .ZN(n793) );
  AND2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n815) );
  AND2_X1 U894 ( .A1(n799), .A2(n877), .ZN(n1006) );
  NOR2_X1 U895 ( .A1(G1996), .A2(n857), .ZN(n800) );
  XOR2_X1 U896 ( .A(KEYINPUT103), .B(n800), .Z(n999) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n801) );
  AND2_X1 U898 ( .A1(n909), .A2(n873), .ZN(n993) );
  NOR2_X1 U899 ( .A1(n801), .A2(n993), .ZN(n802) );
  NOR2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n999), .A2(n804), .ZN(n805) );
  XNOR2_X1 U902 ( .A(n805), .B(KEYINPUT39), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U904 ( .A(KEYINPUT104), .B(n808), .Z(n809) );
  NOR2_X1 U905 ( .A1(n1006), .A2(n809), .ZN(n810) );
  XNOR2_X1 U906 ( .A(KEYINPUT105), .B(n810), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U908 ( .A(KEYINPUT106), .B(n813), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n816), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n817), .ZN(G217) );
  INV_X1 U912 ( .A(n817), .ZN(G223) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U914 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(G188) );
  XOR2_X1 U917 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(G325) );
  XNOR2_X1 U919 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(n823), .ZN(G319) );
  XOR2_X1 U924 ( .A(G2096), .B(KEYINPUT43), .Z(n825) );
  XNOR2_X1 U925 ( .A(G2090), .B(G2678), .ZN(n824) );
  XNOR2_X1 U926 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U927 ( .A(n826), .B(KEYINPUT110), .Z(n828) );
  XOR2_X1 U928 ( .A(G2067), .B(n982), .Z(n827) );
  XNOR2_X1 U929 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U930 ( .A(KEYINPUT42), .B(G2100), .Z(n830) );
  XNOR2_X1 U931 ( .A(G2084), .B(G2078), .ZN(n829) );
  XNOR2_X1 U932 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n832), .B(n831), .ZN(G227) );
  XOR2_X1 U934 ( .A(G1976), .B(G1971), .Z(n834) );
  XNOR2_X1 U935 ( .A(G1961), .B(G1956), .ZN(n833) );
  XNOR2_X1 U936 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U937 ( .A(n835), .B(G2474), .Z(n837) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U940 ( .A(KEYINPUT41), .B(G1986), .Z(n839) );
  XNOR2_X1 U941 ( .A(G1966), .B(G1981), .ZN(n838) );
  XNOR2_X1 U942 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(G229) );
  NAND2_X1 U944 ( .A1(G124), .A2(n861), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n842), .B(KEYINPUT44), .ZN(n845) );
  NAND2_X1 U946 ( .A1(G100), .A2(n858), .ZN(n843) );
  XOR2_X1 U947 ( .A(KEYINPUT111), .B(n843), .Z(n844) );
  NAND2_X1 U948 ( .A1(n845), .A2(n844), .ZN(n849) );
  NAND2_X1 U949 ( .A1(G136), .A2(n559), .ZN(n847) );
  NAND2_X1 U950 ( .A1(G112), .A2(n862), .ZN(n846) );
  NAND2_X1 U951 ( .A1(n847), .A2(n846), .ZN(n848) );
  NOR2_X1 U952 ( .A1(n849), .A2(n848), .ZN(G162) );
  NAND2_X1 U953 ( .A1(G130), .A2(n861), .ZN(n851) );
  NAND2_X1 U954 ( .A1(G118), .A2(n862), .ZN(n850) );
  NAND2_X1 U955 ( .A1(n851), .A2(n850), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G106), .A2(n858), .ZN(n853) );
  NAND2_X1 U957 ( .A1(G142), .A2(n559), .ZN(n852) );
  NAND2_X1 U958 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U959 ( .A(KEYINPUT45), .B(n854), .Z(n855) );
  NOR2_X1 U960 ( .A1(n856), .A2(n855), .ZN(n870) );
  XOR2_X1 U961 ( .A(n857), .B(n992), .Z(n868) );
  NAND2_X1 U962 ( .A1(G103), .A2(n858), .ZN(n860) );
  NAND2_X1 U963 ( .A1(G139), .A2(n559), .ZN(n859) );
  NAND2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G127), .A2(n861), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G115), .A2(n862), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(KEYINPUT47), .B(n865), .Z(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n981) );
  XNOR2_X1 U970 ( .A(n868), .B(n981), .ZN(n869) );
  XOR2_X1 U971 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U972 ( .A(G164), .B(G162), .ZN(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n879) );
  XOR2_X1 U974 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n875) );
  XNOR2_X1 U975 ( .A(G160), .B(n873), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n880) );
  NOR2_X1 U979 ( .A1(G37), .A2(n880), .ZN(G395) );
  XOR2_X1 U980 ( .A(n881), .B(G286), .Z(n883) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n885) );
  XOR2_X1 U982 ( .A(n928), .B(G171), .Z(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U984 ( .A1(G37), .A2(n886), .ZN(G397) );
  XOR2_X1 U985 ( .A(G2454), .B(G2435), .Z(n888) );
  XNOR2_X1 U986 ( .A(G2438), .B(G2427), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n895) );
  XOR2_X1 U988 ( .A(KEYINPUT107), .B(G2446), .Z(n890) );
  XNOR2_X1 U989 ( .A(G2443), .B(G2430), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(n891), .B(G2451), .Z(n893) );
  XOR2_X1 U992 ( .A(G1348), .B(n932), .Z(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n896), .A2(G14), .ZN(n902) );
  NAND2_X1 U996 ( .A1(G319), .A2(n902), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n897) );
  XNOR2_X1 U998 ( .A(KEYINPUT49), .B(n897), .ZN(n898) );
  NOR2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  INV_X1 U1004 ( .A(n902), .ZN(G401) );
  XNOR2_X1 U1005 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1018) );
  INV_X1 U1006 ( .A(KEYINPUT55), .ZN(n1008) );
  XNOR2_X1 U1007 ( .A(n1008), .B(KEYINPUT119), .ZN(n923) );
  XNOR2_X1 U1008 ( .A(G2090), .B(G35), .ZN(n918) );
  XOR2_X1 U1009 ( .A(G2067), .B(G26), .Z(n908) );
  XOR2_X1 U1010 ( .A(n903), .B(G27), .Z(n905) );
  XNOR2_X1 U1011 ( .A(G32), .B(G1996), .ZN(n904) );
  NOR2_X1 U1012 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1013 ( .A(n906), .B(KEYINPUT118), .ZN(n907) );
  NAND2_X1 U1014 ( .A1(n908), .A2(n907), .ZN(n915) );
  XOR2_X1 U1015 ( .A(G33), .B(G2072), .Z(n913) );
  XNOR2_X1 U1016 ( .A(n909), .B(G25), .ZN(n910) );
  NAND2_X1 U1017 ( .A1(n910), .A2(G28), .ZN(n911) );
  XNOR2_X1 U1018 ( .A(n911), .B(KEYINPUT117), .ZN(n912) );
  NAND2_X1 U1019 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1020 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1021 ( .A(KEYINPUT53), .B(n916), .ZN(n917) );
  NOR2_X1 U1022 ( .A1(n918), .A2(n917), .ZN(n921) );
  XOR2_X1 U1023 ( .A(G2084), .B(G34), .Z(n919) );
  XNOR2_X1 U1024 ( .A(KEYINPUT54), .B(n919), .ZN(n920) );
  NAND2_X1 U1025 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1026 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1027 ( .A1(G29), .A2(n924), .ZN(n1016) );
  INV_X1 U1028 ( .A(G16), .ZN(n978) );
  XOR2_X1 U1029 ( .A(n978), .B(KEYINPUT56), .Z(n953) );
  XNOR2_X1 U1030 ( .A(KEYINPUT121), .B(n925), .ZN(n927) );
  NAND2_X1 U1031 ( .A1(G1971), .A2(G303), .ZN(n926) );
  NAND2_X1 U1032 ( .A1(n927), .A2(n926), .ZN(n944) );
  XOR2_X1 U1033 ( .A(n928), .B(G1348), .Z(n930) );
  XNOR2_X1 U1034 ( .A(G299), .B(G1956), .ZN(n929) );
  NOR2_X1 U1035 ( .A1(n930), .A2(n929), .ZN(n942) );
  XOR2_X1 U1036 ( .A(n932), .B(n931), .Z(n934) );
  XOR2_X1 U1037 ( .A(G301), .B(G1961), .Z(n933) );
  NAND2_X1 U1038 ( .A1(n934), .A2(n933), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT122), .B(n945), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G168), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(n946), .B(KEYINPUT120), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(KEYINPUT57), .B(n949), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n980) );
  XOR2_X1 U1051 ( .A(G1986), .B(G24), .Z(n956) );
  XNOR2_X1 U1052 ( .A(G1976), .B(KEYINPUT125), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(n954), .B(G23), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(G22), .B(G1971), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1057 ( .A(KEYINPUT58), .B(n959), .Z(n975) );
  XOR2_X1 U1058 ( .A(G1961), .B(G5), .Z(n970) );
  XOR2_X1 U1059 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n968) );
  XOR2_X1 U1060 ( .A(G19), .B(G1341), .Z(n963) );
  XNOR2_X1 U1061 ( .A(G1956), .B(G20), .ZN(n961) );
  XNOR2_X1 U1062 ( .A(G1981), .B(G6), .ZN(n960) );
  NOR2_X1 U1063 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1064 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1065 ( .A(KEYINPUT59), .B(G1348), .Z(n964) );
  XNOR2_X1 U1066 ( .A(G4), .B(n964), .ZN(n965) );
  NOR2_X1 U1067 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1068 ( .A(n968), .B(n967), .ZN(n969) );
  NAND2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(G21), .B(G1966), .ZN(n971) );
  NOR2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1072 ( .A(KEYINPUT124), .B(n973), .Z(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(KEYINPUT61), .B(n976), .ZN(n977) );
  NAND2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n1013) );
  XNOR2_X1 U1077 ( .A(G164), .B(G2078), .ZN(n985) );
  XOR2_X1 U1078 ( .A(n982), .B(n981), .Z(n983) );
  XNOR2_X1 U1079 ( .A(n983), .B(KEYINPUT114), .ZN(n984) );
  NAND2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(n986), .B(KEYINPUT115), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(KEYINPUT50), .B(n987), .ZN(n1004) );
  XNOR2_X1 U1083 ( .A(G160), .B(G2084), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT112), .B(n996), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G2090), .B(G162), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(n997), .B(KEYINPUT113), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(KEYINPUT51), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(G29), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(KEYINPUT116), .B(n1011), .Z(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(G11), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(n1018), .B(n1017), .ZN(G311) );
  XNOR2_X1 U1104 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

