//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n203), .B1(new_n204), .B2(G13), .ZN(new_n205));
  INV_X1    g0005(.A(G13), .ZN(new_n206));
  NAND4_X1  g0006(.A1(new_n206), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n213), .B(new_n218), .C1(G107), .C2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G116), .A2(G270), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n204), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n227), .A2(new_n211), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n210), .B(new_n231), .C1(new_n234), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G226), .B(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G159), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT72), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT68), .B(G58), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(new_n211), .ZN(new_n261));
  OR2_X1    g0061(.A1(KEYINPUT68), .A2(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT68), .A2(G58), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n262), .A2(KEYINPUT72), .A3(G68), .A4(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n261), .A2(new_n235), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n258), .B1(new_n265), .B2(G20), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT7), .ZN(new_n269));
  NOR4_X1   g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .A4(G20), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n269), .B1(new_n271), .B2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n267), .A2(new_n268), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n233), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT71), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(new_n269), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n270), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n266), .B(KEYINPUT16), .C1(new_n278), .C2(new_n211), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n232), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT67), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(KEYINPUT67), .A3(new_n232), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT7), .B1(new_n274), .B2(new_n233), .ZN(new_n286));
  OAI21_X1  g0086(.A(G68), .B1(new_n286), .B2(new_n270), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n266), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n279), .B(new_n285), .C1(new_n288), .C2(KEYINPUT16), .ZN(new_n289));
  INV_X1    g0089(.A(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  OAI211_X1 g0091(.A(G1), .B(G13), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n223), .A2(G1698), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n271), .B(new_n293), .C1(G223), .C2(G1698), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G87), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G1), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G41), .B2(G45), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n292), .A2(new_n298), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n228), .ZN(new_n303));
  OAI21_X1  g0103(.A(G200), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n296), .A2(new_n303), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G190), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT8), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n227), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n260), .B2(new_n307), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n297), .A2(G13), .A3(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n285), .B1(new_n297), .B2(G20), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n309), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n289), .A2(new_n304), .A3(new_n306), .A4(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT17), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n289), .A2(new_n313), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n305), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(G179), .B2(new_n305), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT18), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n211), .A2(G20), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n233), .A2(G33), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n325), .B1(new_n326), .B2(new_n224), .C1(new_n256), .C2(new_n222), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n327), .A2(new_n285), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(KEYINPUT11), .ZN(new_n330));
  INV_X1    g0130(.A(new_n310), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n211), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT12), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n312), .A2(G68), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n329), .A2(new_n330), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n228), .A2(G1698), .ZN(new_n337));
  OAI221_X1 g0137(.A(new_n337), .B1(G226), .B2(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G33), .A2(G97), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(G33), .A2(G41), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n232), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n300), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n302), .A2(new_n212), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n336), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n292), .B1(new_n338), .B2(new_n339), .ZN(new_n347));
  NOR4_X1   g0147(.A1(new_n347), .A2(new_n344), .A3(KEYINPUT13), .A4(new_n300), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n335), .B1(new_n349), .B2(G190), .ZN(new_n350));
  OAI21_X1  g0150(.A(G200), .B1(new_n346), .B2(new_n348), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(G169), .B1(new_n346), .B2(new_n348), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT14), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n349), .A2(G179), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(G169), .C1(new_n346), .C2(new_n348), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n335), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n324), .A2(new_n353), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G1698), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G222), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G223), .A2(G1698), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n271), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n342), .C1(G77), .C2(new_n271), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n366), .B(new_n301), .C1(new_n302), .C2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(G179), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n235), .B2(G50), .ZN(new_n372));
  INV_X1    g0172(.A(G150), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n372), .B1(new_n373), .B2(new_n256), .C1(new_n309), .C2(new_n326), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n374), .A2(new_n285), .B1(new_n312), .B2(G50), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n331), .A2(new_n222), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI211_X1 g0178(.A(new_n371), .B(new_n378), .C1(new_n318), .C2(new_n370), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n370), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n378), .B2(KEYINPUT9), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n370), .A2(G200), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n378), .A2(KEYINPUT9), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT10), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n385), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT10), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(new_n383), .A4(new_n382), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n379), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT69), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G238), .A2(G1698), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n271), .B(new_n392), .C1(new_n228), .C2(G1698), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n393), .B(new_n342), .C1(G107), .C2(new_n271), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n301), .C1(new_n225), .C2(new_n302), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G200), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT8), .B(G58), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT15), .B(G87), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n326), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n285), .B1(new_n312), .B2(G77), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n331), .A2(new_n224), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n391), .B1(new_n397), .B2(new_n405), .ZN(new_n406));
  OR2_X1    g0206(.A1(new_n395), .A2(new_n380), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n396), .A2(KEYINPUT69), .A3(new_n404), .A4(new_n403), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n395), .A2(G179), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n395), .A2(new_n318), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n405), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n413), .A2(KEYINPUT70), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(KEYINPUT70), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n390), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n361), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G264), .A2(G1698), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n418), .B1(new_n217), .B2(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n419));
  INV_X1    g0219(.A(G303), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n274), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n421), .A3(new_n342), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT5), .B(G41), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n297), .A2(G45), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(G274), .A3(new_n425), .ZN(new_n426));
  XOR2_X1   g0226(.A(KEYINPUT5), .B(G41), .Z(new_n427));
  OAI211_X1 g0227(.A(G270), .B(new_n292), .C1(new_n427), .C2(new_n424), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n422), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G116), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n331), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n280), .A2(new_n232), .B1(G20), .B2(new_n430), .ZN(new_n432));
  AOI21_X1  g0232(.A(G20), .B1(G33), .B2(G283), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G33), .B2(new_n216), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n432), .A2(new_n434), .A3(KEYINPUT20), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT20), .B1(new_n432), .B2(new_n434), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n297), .A2(G33), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n283), .A2(new_n310), .A3(new_n438), .A4(new_n284), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(new_n430), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n429), .B(G169), .C1(new_n437), .C2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT21), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n432), .A2(new_n434), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT20), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n432), .A2(new_n434), .A3(KEYINPUT20), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n280), .A2(KEYINPUT67), .A3(new_n232), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT67), .B1(new_n280), .B2(new_n232), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(G116), .A3(new_n310), .A4(new_n438), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n452), .A3(new_n431), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n453), .A2(KEYINPUT21), .A3(G169), .A4(new_n429), .ZN(new_n454));
  INV_X1    g0254(.A(G179), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n429), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n453), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n443), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n429), .A2(new_n380), .ZN(new_n459));
  INV_X1    g0259(.A(new_n453), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n429), .A2(G200), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n458), .A2(KEYINPUT76), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n462), .A2(new_n443), .A3(new_n457), .A4(new_n454), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT76), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n233), .A2(G33), .A3(G116), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n233), .A2(G107), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT23), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT3), .A2(G33), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT3), .A2(G33), .ZN(new_n472));
  AOI21_X1  g0272(.A(G20), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT22), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n214), .A2(KEYINPUT77), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n474), .B1(new_n473), .B2(new_n475), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n468), .B(new_n470), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT24), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n475), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(KEYINPUT24), .A3(new_n468), .A4(new_n470), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(new_n485), .A3(new_n285), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n439), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n310), .A2(G107), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n489), .B(KEYINPUT25), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(G250), .B(new_n362), .C1(new_n267), .C2(new_n268), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT78), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT78), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n271), .A2(new_n494), .A3(G250), .A4(new_n362), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G294), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n493), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n342), .B1(new_n423), .B2(new_n425), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n498), .A2(new_n342), .B1(G264), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n426), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n318), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G179), .B2(new_n501), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(G190), .A3(new_n426), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n486), .A2(new_n488), .A3(new_n504), .A4(new_n490), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n500), .A2(new_n426), .ZN(new_n506));
  INV_X1    g0306(.A(G200), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n491), .A2(new_n503), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  AND2_X1   g0310(.A1(G97), .A2(G107), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n487), .A2(KEYINPUT6), .A3(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G20), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n255), .A2(G77), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n233), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n487), .B1(new_n272), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n285), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n310), .A2(G97), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n523), .C1(new_n216), .C2(new_n439), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n499), .A2(G257), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n215), .B1(new_n471), .B2(new_n472), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n362), .A2(G244), .ZN(new_n530));
  OAI211_X1 g0330(.A(KEYINPUT73), .B(new_n528), .C1(new_n274), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n271), .A2(G244), .A3(new_n362), .A4(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n527), .A2(new_n529), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n525), .B1(new_n534), .B2(new_n342), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(new_n455), .A3(new_n426), .ZN(new_n536));
  INV_X1    g0336(.A(new_n426), .ZN(new_n537));
  AOI211_X1 g0337(.A(new_n537), .B(new_n525), .C1(new_n534), .C2(new_n342), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n524), .B(new_n536), .C1(new_n538), .C2(G169), .ZN(new_n539));
  OAI21_X1  g0339(.A(G107), .B1(new_n286), .B2(new_n270), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n515), .A2(G20), .B1(G77), .B2(new_n255), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n451), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n439), .A2(new_n216), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n542), .A2(new_n543), .A3(new_n522), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n534), .A2(new_n342), .ZN(new_n545));
  INV_X1    g0345(.A(new_n525), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(G190), .A3(new_n426), .A4(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n544), .B(new_n547), .C1(new_n538), .C2(new_n507), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT75), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n212), .A2(new_n362), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n225), .A2(G1698), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n551), .C1(new_n267), .C2(new_n268), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G33), .A2(G116), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n292), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n425), .A2(KEYINPUT74), .A3(G274), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n424), .B(G250), .C1(new_n341), .C2(new_n232), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT74), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n424), .B2(new_n299), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(G169), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n554), .A2(new_n559), .A3(G179), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n549), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n455), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n564), .B(KEYINPUT75), .C1(G169), .C2(new_n560), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n512), .A2(new_n214), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n339), .A2(new_n233), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(KEYINPUT19), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n233), .B(G68), .C1(new_n267), .C2(new_n268), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n339), .B2(G20), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(new_n285), .B1(new_n331), .B2(new_n401), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n439), .B2(new_n401), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n563), .A2(new_n565), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n451), .A2(G87), .A3(new_n310), .A4(new_n438), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n572), .A2(new_n285), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n401), .A2(new_n331), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n560), .A2(G190), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n507), .C2(new_n560), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n539), .A2(new_n548), .A3(new_n575), .A4(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n509), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n417), .A2(new_n467), .A3(new_n584), .ZN(G372));
  OAI21_X1  g0385(.A(new_n360), .B1(new_n352), .B2(new_n412), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n315), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT18), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n322), .B(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n587), .A2(new_n589), .B1(new_n386), .B2(new_n389), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n379), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n591), .A2(KEYINPUT85), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(KEYINPUT85), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n539), .A2(new_n548), .ZN(new_n595));
  AOI21_X1  g0395(.A(G169), .B1(new_n500), .B2(new_n426), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(new_n455), .B2(new_n506), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n458), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT82), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n559), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT79), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n554), .A2(new_n604), .ZN(new_n605));
  AOI211_X1 g0405(.A(KEYINPUT79), .B(new_n292), .C1(new_n552), .C2(new_n553), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n318), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n608), .A2(new_n574), .A3(new_n564), .ZN(new_n609));
  INV_X1    g0409(.A(new_n581), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n579), .A2(KEYINPUT80), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT80), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n573), .A2(new_n612), .A3(new_n576), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n611), .A2(new_n613), .B1(G200), .B2(new_n607), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT81), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n613), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n612), .B1(new_n573), .B2(new_n576), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n607), .A2(G200), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT81), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n609), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n505), .ZN(new_n623));
  INV_X1    g0423(.A(new_n508), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT82), .B1(new_n599), .B2(new_n458), .ZN(new_n627));
  OR3_X1    g0427(.A1(new_n602), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g0428(.A(new_n609), .B(KEYINPUT83), .Z(new_n629));
  INV_X1    g0429(.A(new_n539), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n622), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g0433(.A(KEYINPUT84), .B(KEYINPUT26), .Z(new_n634));
  AND4_X1   g0434(.A1(new_n630), .A2(new_n575), .A3(new_n582), .A4(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n629), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n628), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n417), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n594), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT86), .ZN(G369));
  NOR2_X1   g0441(.A1(new_n206), .A2(G20), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OR3_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .A3(G1), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT27), .B1(new_n643), .B2(G1), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n491), .A2(new_n649), .ZN(new_n650));
  OR3_X1    g0450(.A1(new_n509), .A2(new_n650), .A3(KEYINPUT87), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT87), .B1(new_n509), .B2(new_n650), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n599), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n648), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n460), .A2(new_n649), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n463), .B2(new_n466), .ZN(new_n657));
  INV_X1    g0457(.A(new_n458), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n656), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G330), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n655), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n599), .A2(new_n648), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n458), .A2(new_n648), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n651), .B2(new_n652), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n665), .A2(new_n666), .A3(new_n669), .ZN(G399));
  NAND3_X1  g0470(.A1(new_n208), .A2(KEYINPUT88), .A3(new_n291), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT88), .B1(new_n208), .B2(new_n291), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G1), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n512), .A2(new_n214), .A3(new_n430), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n676), .A2(new_n677), .B1(new_n236), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n638), .A2(new_n649), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(KEYINPUT29), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n630), .A2(new_n575), .A3(new_n582), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n631), .A2(new_n632), .B1(new_n683), .B2(new_n634), .ZN(new_n684));
  INV_X1    g0484(.A(new_n629), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n622), .A2(new_n600), .A3(new_n625), .A4(new_n595), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n682), .B1(new_n687), .B2(new_n649), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT92), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n493), .A2(new_n495), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n497), .A2(new_n496), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n342), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n499), .A2(G264), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(KEYINPUT89), .A3(new_n694), .A4(new_n560), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n456), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT89), .B1(new_n500), .B2(new_n560), .ZN(new_n697));
  INV_X1    g0497(.A(new_n535), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT91), .B1(new_n699), .B2(KEYINPUT30), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT30), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT90), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n607), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n603), .B(KEYINPUT90), .C1(new_n605), .C2(new_n606), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(new_n429), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n538), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n705), .A2(new_n455), .A3(new_n501), .A4(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n693), .A2(new_n694), .A3(new_n560), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT89), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n456), .A3(new_n535), .A4(new_n695), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT91), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n700), .A2(new_n701), .A3(new_n707), .A4(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT31), .B1(new_n715), .B2(new_n648), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n713), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n701), .A2(new_n707), .A3(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n690), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n648), .ZN(new_n721));
  AND3_X1   g0521(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n712), .B1(new_n711), .B2(new_n713), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n703), .A2(new_n429), .A3(new_n704), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n725), .A2(G179), .A3(new_n538), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n726), .A2(new_n501), .B1(KEYINPUT30), .B2(new_n699), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n649), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT92), .B(new_n721), .C1(new_n728), .C2(KEYINPUT31), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n623), .A2(new_n624), .B1(new_n597), .B2(new_n598), .ZN(new_n730));
  AND4_X1   g0530(.A1(new_n539), .A2(new_n548), .A3(new_n575), .A4(new_n582), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n467), .A2(new_n730), .A3(new_n731), .A4(new_n649), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT93), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n584), .A2(KEYINPUT93), .A3(new_n467), .A4(new_n649), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n720), .A2(new_n729), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n689), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n679), .B1(new_n740), .B2(G1), .ZN(G364));
  INV_X1    g0541(.A(KEYINPUT94), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n663), .B(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n297), .B1(new_n642), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n674), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n661), .A2(new_n662), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n744), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n748), .B1(new_n661), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n380), .A2(new_n507), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n233), .A2(G179), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n271), .B1(new_n757), .B2(new_n214), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n233), .A2(new_n455), .A3(KEYINPUT96), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT96), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(G20), .B2(G179), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n507), .A2(G190), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n756), .A2(new_n766), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n765), .A2(new_n224), .B1(new_n487), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n380), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n455), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n758), .B(new_n768), .C1(G97), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n763), .A2(new_n769), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT97), .ZN(new_n774));
  INV_X1    g0574(.A(new_n260), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n763), .A2(new_n766), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n763), .A2(new_n755), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n778), .A2(G68), .B1(new_n780), .B2(G50), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n756), .A2(new_n764), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n257), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n772), .A2(new_n776), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n765), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n774), .A2(G322), .ZN(new_n788));
  INV_X1    g0588(.A(new_n767), .ZN(new_n789));
  INV_X1    g0589(.A(new_n782), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G283), .A2(new_n789), .B1(new_n790), .B2(G329), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT98), .ZN(new_n792));
  INV_X1    g0592(.A(new_n757), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n780), .A2(G326), .B1(G303), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n771), .ZN(new_n795));
  INV_X1    g0595(.A(G294), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n274), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(new_n778), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n788), .A2(new_n792), .A3(new_n794), .A4(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n785), .B1(new_n787), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n232), .B1(G20), .B2(new_n318), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n208), .A2(G355), .A3(new_n271), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n250), .A2(G45), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT95), .ZN(new_n806));
  INV_X1    g0606(.A(new_n208), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n271), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(G45), .B2(new_n236), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n804), .B1(G116), .B2(new_n208), .C1(new_n806), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n753), .A2(new_n802), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n754), .A2(new_n803), .A3(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n750), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n405), .A2(new_n648), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n409), .A2(new_n412), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT100), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n409), .A2(KEYINPUT100), .A3(new_n412), .A4(new_n816), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n602), .A2(new_n626), .A3(new_n627), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT26), .B1(new_n622), .B2(new_n630), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n685), .B1(new_n824), .B2(new_n635), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n822), .B(new_n649), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n680), .ZN(new_n827));
  INV_X1    g0627(.A(new_n412), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n648), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n821), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n826), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(new_n738), .Z(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n748), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n274), .B1(new_n786), .B2(new_n782), .C1(new_n765), .C2(new_n430), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n774), .A2(G294), .B1(G97), .B2(new_n771), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n778), .A2(G283), .B1(G87), .B2(new_n789), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(new_n487), .C2(new_n757), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n834), .B(new_n837), .C1(G303), .C2(new_n780), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT99), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n774), .A2(G143), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n778), .A2(G150), .B1(new_n780), .B2(G137), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n840), .B(new_n841), .C1(new_n257), .C2(new_n765), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT34), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n271), .B1(new_n260), .B2(new_n795), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n842), .A2(new_n843), .B1(G50), .B2(new_n793), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n211), .B2(new_n767), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n844), .B(new_n846), .C1(G132), .C2(new_n790), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n802), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n802), .A2(new_n751), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n224), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n819), .A2(new_n820), .B1(new_n828), .B2(new_n648), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n751), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n848), .A2(new_n747), .A3(new_n850), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n833), .A2(new_n853), .ZN(G384));
  AOI21_X1  g0654(.A(new_n430), .B1(new_n515), .B2(KEYINPUT35), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n855), .B(new_n234), .C1(KEYINPUT35), .C2(new_n515), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  NAND4_X1  g0657(.A1(new_n261), .A2(G77), .A3(new_n237), .A4(new_n264), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n222), .A2(G68), .ZN(new_n859));
  AOI21_X1  g0659(.A(G13), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n857), .B1(G1), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT101), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n412), .A2(new_n648), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n826), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n335), .A2(new_n648), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT102), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n359), .A2(new_n867), .A3(new_n335), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n359), .B2(new_n335), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n353), .B(new_n866), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n359), .A2(new_n335), .A3(new_n648), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n865), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n279), .A2(new_n285), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n276), .B1(new_n275), .B2(new_n269), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n519), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(G68), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT16), .B1(new_n878), .B2(new_n266), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n313), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT103), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n646), .ZN(new_n883));
  OAI211_X1 g0683(.A(KEYINPUT103), .B(new_n313), .C1(new_n874), .C2(new_n879), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n882), .A2(KEYINPUT104), .A3(new_n883), .A4(new_n884), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n882), .A2(new_n321), .A3(new_n884), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n887), .A2(new_n314), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT105), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n289), .A2(new_n313), .B1(new_n320), .B2(new_n646), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n314), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n895), .B2(KEYINPUT37), .ZN(new_n896));
  INV_X1    g0696(.A(new_n314), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(new_n893), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(KEYINPUT105), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n891), .A2(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n589), .A2(new_n315), .B1(new_n887), .B2(new_n888), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n890), .A2(KEYINPUT37), .B1(new_n896), .B2(new_n900), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n906), .B1(new_n907), .B2(new_n903), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n873), .A2(new_n909), .B1(new_n323), .B2(new_n646), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n907), .A2(new_n906), .A3(new_n903), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT105), .B1(new_n898), .B2(new_n899), .ZN(new_n914));
  NOR4_X1   g0714(.A1(new_n897), .A2(new_n893), .A3(new_n892), .A4(KEYINPUT37), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n317), .A2(new_n883), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n316), .B2(new_n323), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n911), .B1(new_n912), .B2(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n868), .A2(new_n869), .A3(new_n648), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT106), .Z(new_n923));
  NAND3_X1  g0723(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT39), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n910), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n417), .B1(new_n681), .B2(new_n688), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n594), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT108), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n870), .A2(new_n871), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n830), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n728), .A2(KEYINPUT31), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n716), .B1(new_n734), .B2(new_n735), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT107), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n716), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n736), .A2(new_n940), .A3(new_n934), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n872), .A2(new_n851), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT107), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n909), .A2(new_n939), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n903), .B1(new_n891), .B2(new_n901), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n920), .B1(new_n946), .B2(KEYINPUT38), .ZN(new_n947));
  OAI21_X1  g0747(.A(KEYINPUT40), .B1(new_n947), .B2(new_n943), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n949), .A2(new_n941), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(G330), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n662), .B1(new_n935), .B2(new_n934), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n417), .A2(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n950), .A2(new_n417), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n931), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n929), .A2(new_n930), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n955), .B(new_n956), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n642), .A2(new_n297), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n862), .B1(new_n957), .B2(new_n958), .ZN(G367));
  INV_X1    g0759(.A(new_n665), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n595), .B1(new_n544), .B2(new_n649), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n630), .A2(new_n648), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n653), .A2(new_n667), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n965), .A2(KEYINPUT42), .A3(new_n963), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n539), .B1(new_n961), .B2(new_n599), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n649), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT42), .B1(new_n965), .B2(new_n963), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n619), .A2(new_n648), .ZN(new_n971));
  MUX2_X1   g0771(.A(new_n629), .B(new_n622), .S(new_n971), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n970), .A2(KEYINPUT43), .A3(new_n972), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n964), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n974), .A2(new_n975), .ZN(new_n980));
  INV_X1    g0780(.A(new_n964), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n980), .A2(new_n981), .A3(new_n977), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n674), .B(KEYINPUT41), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n653), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(new_n668), .C1(new_n599), .C2(new_n649), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n743), .B1(new_n965), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n664), .B(new_n669), .C1(new_n655), .C2(new_n668), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(new_n689), .A3(new_n738), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n963), .B1(new_n669), .B2(new_n666), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT44), .Z(new_n994));
  NOR3_X1   g0794(.A1(new_n669), .A2(new_n666), .A3(new_n963), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT45), .ZN(new_n996));
  AOI211_X1 g0796(.A(KEYINPUT109), .B(new_n665), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT109), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n960), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n665), .A2(KEYINPUT109), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n994), .A2(new_n999), .A3(new_n1000), .A4(new_n996), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n992), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n985), .B1(new_n1003), .B2(new_n740), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n983), .B1(new_n1004), .B2(new_n746), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n808), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n811), .B1(new_n208), .B2(new_n401), .C1(new_n241), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n765), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1008), .A2(G50), .B1(new_n775), .B2(new_n793), .ZN(new_n1009));
  INV_X1    g0809(.A(G137), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1009), .B1(new_n224), .B2(new_n767), .C1(new_n1010), .C2(new_n782), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G159), .B2(new_n778), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n774), .A2(G150), .B1(G68), .B2(new_n771), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n780), .A2(G143), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1012), .A2(new_n271), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n757), .A2(new_n430), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT46), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n796), .A2(new_n777), .B1(new_n779), .B2(new_n786), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(G317), .C2(new_n790), .ZN(new_n1019));
  INV_X1    g0819(.A(G283), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n765), .A2(new_n1020), .B1(new_n487), .B2(new_n795), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT110), .Z(new_n1022));
  NAND2_X1  g0822(.A1(new_n789), .A2(G97), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n774), .A2(G303), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1015), .B1(new_n271), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT47), .Z(new_n1027));
  INV_X1    g0827(.A(new_n802), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n747), .B(new_n1007), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n972), .A2(G20), .A3(new_n752), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1005), .A2(new_n1032), .ZN(G387));
  OAI21_X1  g0833(.A(new_n739), .B1(new_n988), .B2(new_n989), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1034), .A2(new_n674), .A3(new_n991), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n655), .A2(new_n753), .ZN(new_n1036));
  INV_X1    g0836(.A(G45), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n246), .A2(new_n1037), .A3(new_n271), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n399), .A2(new_n222), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1039), .A2(KEYINPUT50), .B1(G68), .B2(G77), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n1037), .C1(KEYINPUT50), .C2(new_n1039), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n677), .B1(new_n1041), .B2(new_n274), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n208), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n811), .C1(new_n487), .C2(new_n208), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1036), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n795), .A2(new_n401), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n774), .B2(G50), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT111), .Z(new_n1048));
  NOR2_X1   g0848(.A1(new_n757), .A2(new_n224), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n271), .B1(new_n765), .B2(new_n211), .C1(new_n257), .C2(new_n779), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G150), .C2(new_n790), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n777), .A2(new_n309), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1048), .A2(new_n1023), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n774), .A2(G317), .B1(G303), .B2(new_n1008), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n778), .A2(G311), .ZN(new_n1055));
  XOR2_X1   g0855(.A(KEYINPUT112), .B(G322), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n780), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(KEYINPUT113), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(KEYINPUT113), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT48), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1061), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1063), .A2(new_n1064), .A3(new_n1059), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G283), .A2(new_n771), .B1(new_n793), .B2(G294), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(KEYINPUT49), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n789), .A2(G116), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n790), .A2(G326), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1068), .A2(new_n274), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(KEYINPUT49), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1053), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1045), .B1(new_n1073), .B2(new_n802), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n746), .A2(new_n990), .B1(new_n1074), .B2(new_n747), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1035), .A2(new_n1075), .ZN(G393));
  AOI22_X1  g0876(.A1(G107), .A2(new_n789), .B1(new_n790), .B2(new_n1056), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n274), .C1(new_n765), .C2(new_n796), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n774), .A2(G311), .B1(G317), .B2(new_n780), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT114), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT52), .Z(new_n1081));
  AOI211_X1 g0881(.A(new_n1078), .B(new_n1081), .C1(G283), .C2(new_n793), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n430), .B2(new_n795), .C1(new_n420), .C2(new_n777), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n774), .A2(G159), .B1(G150), .B2(new_n780), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT51), .Z(new_n1085));
  NOR2_X1   g0885(.A1(new_n795), .A2(new_n224), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n271), .B1(new_n777), .B2(new_n222), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(G68), .C2(new_n793), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1008), .A2(new_n399), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G87), .A2(new_n789), .B1(new_n790), .B2(G143), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1085), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1028), .B1(new_n1083), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n963), .A2(new_n753), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n811), .B1(new_n216), .B2(new_n208), .C1(new_n1006), .C2(new_n253), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1092), .A2(new_n748), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n994), .A2(new_n996), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n998), .A3(new_n960), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1001), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1096), .B1(new_n1099), .B2(new_n746), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n674), .B1(new_n1099), .B2(new_n992), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n991), .B1(new_n1098), .B2(new_n1001), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(G390));
  INV_X1    g0903(.A(KEYINPUT116), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n826), .A2(new_n864), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n872), .B1(new_n738), .B2(new_n851), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n952), .A2(new_n942), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n737), .A2(G330), .A3(new_n942), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT115), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n737), .A2(new_n942), .A3(KEYINPUT115), .A4(G330), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n687), .A2(new_n649), .A3(new_n822), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n864), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n941), .A2(G330), .A3(new_n830), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n872), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1105), .A2(new_n1108), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n927), .A2(new_n594), .A3(new_n953), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1104), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n927), .A2(new_n594), .A3(new_n953), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1116), .A2(new_n872), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1115), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n865), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1126));
  OAI211_X1 g0926(.A(KEYINPUT116), .B(new_n1121), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1120), .A2(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT39), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n920), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT39), .B1(new_n905), .B2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1129), .A2(new_n1131), .B1(new_n873), .B2(new_n923), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n872), .B1(new_n1114), .B2(new_n864), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n947), .A2(new_n1133), .A3(new_n923), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1113), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n923), .B1(new_n1105), .B2(new_n932), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n921), .B2(new_n924), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1107), .B1(new_n1139), .B2(new_n1134), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1128), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1120), .A2(new_n1127), .A3(new_n1140), .A4(new_n1137), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n674), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1132), .A2(new_n1135), .B1(new_n942), .B2(new_n952), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1139), .A2(new_n1113), .A3(new_n1134), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n746), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n752), .B1(new_n921), .B2(new_n924), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n309), .A2(new_n849), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT54), .B(G143), .Z(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1010), .A2(new_n777), .B1(new_n765), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n774), .B2(G132), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n771), .A2(G159), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n780), .A2(G128), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n757), .A2(new_n373), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT53), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G50), .A2(new_n789), .B1(new_n790), .B2(G125), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1158), .A2(new_n271), .A3(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1160), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n487), .A2(new_n777), .B1(new_n779), .B2(new_n1020), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n765), .A2(new_n216), .B1(new_n211), .B2(new_n767), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n757), .A2(new_n214), .B1(new_n782), .B2(new_n796), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1086), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n271), .B1(new_n774), .B2(G116), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1028), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1148), .A2(new_n748), .A3(new_n1150), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1147), .A2(KEYINPUT117), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT117), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n745), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n1169), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT118), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1171), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1144), .B1(new_n1176), .B2(new_n1177), .ZN(G378));
  XOR2_X1   g0978(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1179));
  XNOR2_X1  g0979(.A(new_n390), .B(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n377), .A2(new_n883), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n949), .B2(G330), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n662), .B(new_n1182), .C1(new_n945), .C2(new_n948), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n926), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n905), .A2(new_n908), .B1(new_n936), .B2(new_n938), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n936), .B1(new_n912), .B2(new_n920), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1187), .A2(new_n944), .B1(new_n1188), .B2(KEYINPUT40), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1182), .B1(new_n1189), .B2(new_n662), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n926), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n949), .A2(G330), .A3(new_n1183), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1186), .A2(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1120), .A2(new_n1127), .B1(new_n1140), .B2(new_n1137), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(KEYINPUT57), .C1(new_n1119), .C2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1119), .B1(new_n1128), .B2(new_n1141), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1186), .A2(new_n1193), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1196), .A2(new_n1200), .A3(new_n674), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1182), .A2(new_n752), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n765), .A2(new_n401), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G116), .B2(new_n780), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n211), .B2(new_n795), .C1(new_n216), .C2(new_n777), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G283), .B2(new_n790), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n774), .A2(G107), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n271), .B1(new_n789), .B2(new_n775), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1049), .A2(G41), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT58), .Z(new_n1211));
  NAND2_X1  g1011(.A1(new_n774), .A2(G128), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1008), .A2(G137), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G150), .A2(new_n771), .B1(new_n793), .B2(new_n1151), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n778), .A2(G132), .B1(new_n780), .B2(G125), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  XOR2_X1   g1016(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1217));
  OAI21_X1  g1017(.A(new_n291), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT120), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(G124), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1219), .A2(G124), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n782), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1218), .A2(G33), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n257), .C2(new_n767), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n222), .B1(new_n267), .B2(G41), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n802), .B1(new_n1211), .B2(new_n1227), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT121), .Z(new_n1229));
  AOI211_X1 g1029(.A(new_n1202), .B(new_n1229), .C1(new_n222), .C2(new_n849), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1194), .A2(new_n746), .B1(new_n747), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1201), .A2(new_n1231), .ZN(G375));
  NAND2_X1  g1032(.A1(new_n872), .A2(new_n751), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n849), .A2(new_n211), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n274), .B1(new_n779), .B2(new_n796), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1046), .B(new_n1235), .C1(G116), .C2(new_n778), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n774), .A2(G283), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n793), .A2(G97), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1008), .A2(G107), .B1(G77), .B2(new_n789), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n782), .A2(new_n420), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n271), .B1(new_n222), .B2(new_n795), .C1(new_n765), .C2(new_n373), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G132), .B2(new_n780), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n790), .A2(G128), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n774), .A2(G137), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n778), .A2(new_n1151), .B1(new_n775), .B2(new_n789), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n757), .A2(new_n257), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n1240), .A2(new_n1241), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n802), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1233), .A2(new_n747), .A3(new_n1234), .A4(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1118), .B2(new_n745), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n984), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1253), .B1(new_n1128), .B2(new_n1255), .ZN(G381));
  AND3_X1   g1056(.A1(new_n1144), .A2(new_n1174), .A3(new_n1171), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1201), .A2(new_n1231), .A3(new_n1257), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n979), .A2(new_n982), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n984), .B1(new_n1102), .B2(new_n739), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1260), .B2(new_n745), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(new_n1031), .ZN(new_n1262));
  INV_X1    g1062(.A(G384), .ZN(new_n1263));
  INV_X1    g1063(.A(G390), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1035), .A2(new_n814), .A3(new_n1075), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  OR3_X1    g1066(.A1(new_n1258), .A2(G381), .A3(new_n1266), .ZN(G407));
  NAND2_X1  g1067(.A1(new_n647), .A2(G213), .ZN(new_n1268));
  OR3_X1    g1068(.A1(new_n1258), .A2(KEYINPUT122), .A3(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT122), .B1(new_n1258), .B2(new_n1268), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(G407), .A2(new_n1269), .A3(G213), .A4(new_n1270), .ZN(G409));
  NAND3_X1  g1071(.A1(new_n1201), .A2(G378), .A3(new_n1231), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1194), .B1(new_n1119), .B2(new_n1195), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1231), .B1(new_n1273), .B2(new_n985), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1257), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1120), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1254), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT123), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n674), .B1(new_n1254), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1277), .A2(KEYINPUT123), .A3(new_n1254), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1280), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1285), .A2(G384), .A3(new_n1253), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G384), .B1(new_n1285), .B2(new_n1253), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1276), .A2(new_n1288), .A3(new_n1268), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n647), .A2(G213), .A3(G2897), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1277), .A2(KEYINPUT123), .A3(new_n1254), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT123), .B1(new_n1277), .B2(new_n1254), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1293), .A2(new_n1294), .A3(new_n1282), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1263), .B1(new_n1295), .B2(new_n1252), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1285), .A2(G384), .A3(new_n1253), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1291), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1292), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1276), .A2(new_n1268), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1276), .A2(new_n1288), .A3(new_n1304), .A4(new_n1268), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1290), .A2(new_n1302), .A3(new_n1303), .A4(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n814), .B1(new_n1035), .B2(new_n1075), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1265), .A2(new_n1307), .A3(KEYINPUT125), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(G387), .A2(new_n1309), .A3(new_n1264), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1265), .A2(new_n1307), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1264), .B(new_n1311), .C1(new_n1261), .C2(new_n1031), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G390), .B1(new_n1005), .B2(new_n1032), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1312), .B1(new_n1313), .B2(new_n1308), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1262), .A2(G390), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1310), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1306), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT124), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1286), .A2(new_n1287), .A3(new_n1291), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1298), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1318), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1292), .A2(KEYINPUT124), .A3(new_n1299), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(new_n1301), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT126), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1324), .B1(new_n1316), .B2(KEYINPUT61), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(G387), .A2(new_n1264), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1309), .B1(new_n1262), .B2(G390), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1326), .B1(new_n1327), .B2(new_n1312), .ZN(new_n1328));
  OAI211_X1 g1128(.A(KEYINPUT126), .B(new_n1303), .C1(new_n1328), .C2(new_n1310), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1325), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1289), .A2(new_n1331), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1276), .A2(new_n1288), .A3(KEYINPUT63), .A4(new_n1268), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1323), .A2(new_n1330), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1317), .A2(new_n1334), .ZN(G405));
  OAI21_X1  g1135(.A(new_n1316), .B1(new_n1287), .B2(new_n1286), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1288), .B1(new_n1328), .B2(new_n1310), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G375), .A2(new_n1257), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1339), .A2(KEYINPUT127), .A3(new_n1272), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1340), .B1(KEYINPUT127), .B2(new_n1339), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1338), .B(new_n1341), .ZN(G402));
endmodule


