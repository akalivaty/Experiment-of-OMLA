

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X2 U548 ( .A(n657), .Z(n513) );
  XNOR2_X1 U549 ( .A(n596), .B(KEYINPUT64), .ZN(n657) );
  XOR2_X1 U550 ( .A(n600), .B(KEYINPUT28), .Z(n514) );
  AND2_X1 U551 ( .A1(G160), .A2(G40), .ZN(n595) );
  OR2_X1 U552 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U553 ( .A1(G651), .A2(n568), .ZN(n774) );
  XOR2_X1 U554 ( .A(KEYINPUT1), .B(n544), .Z(n775) );
  NOR2_X2 U555 ( .A1(n537), .A2(n536), .ZN(G160) );
  AND2_X1 U556 ( .A1(G2104), .A2(G2105), .ZN(n863) );
  NAND2_X1 U557 ( .A1(G114), .A2(n863), .ZN(n515) );
  XNOR2_X1 U558 ( .A(n515), .B(KEYINPUT86), .ZN(n518) );
  INV_X1 U559 ( .A(G2104), .ZN(n516) );
  NOR2_X4 U560 ( .A1(G2105), .A2(n516), .ZN(n859) );
  NAND2_X1 U561 ( .A1(n859), .A2(G102), .ZN(n517) );
  NAND2_X1 U562 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n519), .Z(n860) );
  NAND2_X1 U565 ( .A1(G138), .A2(n860), .ZN(n523) );
  INV_X1 U566 ( .A(G2104), .ZN(n520) );
  NAND2_X1 U567 ( .A1(n520), .A2(G2105), .ZN(n521) );
  XNOR2_X1 U568 ( .A(n521), .B(KEYINPUT65), .ZN(n865) );
  NAND2_X1 U569 ( .A1(G126), .A2(n865), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U571 ( .A1(n525), .A2(n524), .ZN(G164) );
  NAND2_X1 U572 ( .A1(G101), .A2(n859), .ZN(n528) );
  XNOR2_X1 U573 ( .A(KEYINPUT66), .B(n528), .ZN(n527) );
  INV_X1 U574 ( .A(KEYINPUT23), .ZN(n526) );
  NAND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n531) );
  XOR2_X1 U576 ( .A(KEYINPUT66), .B(n528), .Z(n529) );
  NAND2_X1 U577 ( .A1(n529), .A2(KEYINPUT23), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n533) );
  NAND2_X1 U579 ( .A1(G137), .A2(n860), .ZN(n532) );
  NAND2_X1 U580 ( .A1(n533), .A2(n532), .ZN(n537) );
  NAND2_X1 U581 ( .A1(G113), .A2(n863), .ZN(n535) );
  NAND2_X1 U582 ( .A1(G125), .A2(n865), .ZN(n534) );
  NAND2_X1 U583 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .ZN(n538) );
  XNOR2_X1 U585 ( .A(n538), .B(KEYINPUT67), .ZN(n568) );
  NAND2_X1 U586 ( .A1(G52), .A2(n774), .ZN(n539) );
  XNOR2_X1 U587 ( .A(n539), .B(KEYINPUT69), .ZN(n548) );
  INV_X1 U588 ( .A(G651), .ZN(n543) );
  NOR2_X1 U589 ( .A1(n568), .A2(n543), .ZN(n778) );
  NAND2_X1 U590 ( .A1(G77), .A2(n778), .ZN(n541) );
  NOR2_X1 U591 ( .A1(G543), .A2(G651), .ZN(n779) );
  NAND2_X1 U592 ( .A1(G90), .A2(n779), .ZN(n540) );
  NAND2_X1 U593 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U594 ( .A(n542), .B(KEYINPUT9), .ZN(n546) );
  NOR2_X1 U595 ( .A1(G543), .A2(n543), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G64), .A2(n775), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U598 ( .A1(n548), .A2(n547), .ZN(G171) );
  NAND2_X1 U599 ( .A1(G51), .A2(n774), .ZN(n550) );
  NAND2_X1 U600 ( .A1(G63), .A2(n775), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U602 ( .A(KEYINPUT6), .B(n551), .ZN(n557) );
  NAND2_X1 U603 ( .A1(n779), .A2(G89), .ZN(n552) );
  XNOR2_X1 U604 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U605 ( .A1(G76), .A2(n778), .ZN(n553) );
  NAND2_X1 U606 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U607 ( .A(n555), .B(KEYINPUT5), .Z(n556) );
  NOR2_X1 U608 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U609 ( .A(KEYINPUT7), .B(n558), .Z(n559) );
  XOR2_X1 U610 ( .A(KEYINPUT77), .B(n559), .Z(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(n778), .A2(G75), .ZN(n560) );
  XOR2_X1 U613 ( .A(KEYINPUT81), .B(n560), .Z(n562) );
  NAND2_X1 U614 ( .A1(n779), .A2(G88), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U616 ( .A(KEYINPUT82), .B(n563), .Z(n567) );
  NAND2_X1 U617 ( .A1(G50), .A2(n774), .ZN(n565) );
  NAND2_X1 U618 ( .A1(G62), .A2(n775), .ZN(n564) );
  AND2_X1 U619 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U620 ( .A1(n567), .A2(n566), .ZN(G303) );
  NAND2_X1 U621 ( .A1(G49), .A2(n774), .ZN(n570) );
  NAND2_X1 U622 ( .A1(G87), .A2(n568), .ZN(n569) );
  NAND2_X1 U623 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U624 ( .A1(n775), .A2(n571), .ZN(n573) );
  NAND2_X1 U625 ( .A1(G651), .A2(G74), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n573), .A2(n572), .ZN(G288) );
  NAND2_X1 U627 ( .A1(G61), .A2(n775), .ZN(n574) );
  XNOR2_X1 U628 ( .A(n574), .B(KEYINPUT80), .ZN(n581) );
  NAND2_X1 U629 ( .A1(G86), .A2(n779), .ZN(n576) );
  NAND2_X1 U630 ( .A1(G48), .A2(n774), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U632 ( .A1(n778), .A2(G73), .ZN(n577) );
  XOR2_X1 U633 ( .A(KEYINPUT2), .B(n577), .Z(n578) );
  NOR2_X1 U634 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U635 ( .A1(n581), .A2(n580), .ZN(G305) );
  NAND2_X1 U636 ( .A1(G85), .A2(n779), .ZN(n583) );
  NAND2_X1 U637 ( .A1(G47), .A2(n774), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U639 ( .A1(G72), .A2(n778), .ZN(n584) );
  XOR2_X1 U640 ( .A(KEYINPUT68), .B(n584), .Z(n585) );
  NOR2_X1 U641 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U642 ( .A1(n775), .A2(G60), .ZN(n587) );
  NAND2_X1 U643 ( .A1(n588), .A2(n587), .ZN(G290) );
  NAND2_X1 U644 ( .A1(G53), .A2(n774), .ZN(n590) );
  NAND2_X1 U645 ( .A1(G65), .A2(n775), .ZN(n589) );
  NAND2_X1 U646 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U647 ( .A1(G78), .A2(n778), .ZN(n592) );
  NAND2_X1 U648 ( .A1(G91), .A2(n779), .ZN(n591) );
  NAND2_X1 U649 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U650 ( .A1(n594), .A2(n593), .ZN(n916) );
  NOR2_X1 U651 ( .A1(G164), .A2(G1384), .ZN(n684) );
  NAND2_X1 U652 ( .A1(n684), .A2(n595), .ZN(n596) );
  XNOR2_X1 U653 ( .A(n513), .B(KEYINPUT91), .ZN(n640) );
  NAND2_X1 U654 ( .A1(G2072), .A2(n640), .ZN(n597) );
  XNOR2_X1 U655 ( .A(n597), .B(KEYINPUT27), .ZN(n599) );
  INV_X1 U656 ( .A(G1956), .ZN(n995) );
  NOR2_X1 U657 ( .A1(n640), .A2(n995), .ZN(n598) );
  NOR2_X1 U658 ( .A1(n599), .A2(n598), .ZN(n601) );
  NOR2_X1 U659 ( .A1(n916), .A2(n601), .ZN(n600) );
  NAND2_X1 U660 ( .A1(n916), .A2(n601), .ZN(n636) );
  NAND2_X1 U661 ( .A1(G79), .A2(n778), .ZN(n603) );
  NAND2_X1 U662 ( .A1(G54), .A2(n774), .ZN(n602) );
  NAND2_X1 U663 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U664 ( .A(n604), .B(KEYINPUT75), .ZN(n606) );
  NAND2_X1 U665 ( .A1(G92), .A2(n779), .ZN(n605) );
  NAND2_X1 U666 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U667 ( .A1(n775), .A2(G66), .ZN(n607) );
  XOR2_X1 U668 ( .A(KEYINPUT74), .B(n607), .Z(n608) );
  NOR2_X1 U669 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U670 ( .A(KEYINPUT15), .B(n610), .Z(n882) );
  NAND2_X1 U671 ( .A1(n779), .A2(G81), .ZN(n611) );
  XNOR2_X1 U672 ( .A(n611), .B(KEYINPUT12), .ZN(n613) );
  NAND2_X1 U673 ( .A1(G68), .A2(n778), .ZN(n612) );
  NAND2_X1 U674 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U675 ( .A(n614), .B(KEYINPUT13), .ZN(n616) );
  NAND2_X1 U676 ( .A1(G43), .A2(n774), .ZN(n615) );
  NAND2_X1 U677 ( .A1(n616), .A2(n615), .ZN(n621) );
  XOR2_X1 U678 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n618) );
  NAND2_X1 U679 ( .A1(G56), .A2(n775), .ZN(n617) );
  XNOR2_X1 U680 ( .A(n618), .B(n617), .ZN(n619) );
  XOR2_X1 U681 ( .A(KEYINPUT71), .B(n619), .Z(n620) );
  NOR2_X1 U682 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U683 ( .A(KEYINPUT73), .B(n622), .ZN(n906) );
  INV_X1 U684 ( .A(G1996), .ZN(n623) );
  NOR2_X1 U685 ( .A1(n513), .A2(n623), .ZN(n624) );
  XOR2_X1 U686 ( .A(n624), .B(KEYINPUT26), .Z(n626) );
  NAND2_X1 U687 ( .A1(n513), .A2(G1341), .ZN(n625) );
  NAND2_X1 U688 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U689 ( .A1(n906), .A2(n627), .ZN(n628) );
  OR2_X1 U690 ( .A1(n882), .A2(n628), .ZN(n634) );
  NAND2_X1 U691 ( .A1(n882), .A2(n628), .ZN(n632) );
  NAND2_X1 U692 ( .A1(G2067), .A2(n640), .ZN(n630) );
  NAND2_X1 U693 ( .A1(n513), .A2(G1348), .ZN(n629) );
  NAND2_X1 U694 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U695 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U696 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U697 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U698 ( .A1(n514), .A2(n637), .ZN(n639) );
  XOR2_X1 U699 ( .A(KEYINPUT92), .B(KEYINPUT29), .Z(n638) );
  XNOR2_X1 U700 ( .A(n639), .B(n638), .ZN(n644) );
  XNOR2_X1 U701 ( .A(KEYINPUT25), .B(G2078), .ZN(n932) );
  NAND2_X1 U702 ( .A1(n932), .A2(n640), .ZN(n642) );
  INV_X1 U703 ( .A(G1961), .ZN(n991) );
  NAND2_X1 U704 ( .A1(n513), .A2(n991), .ZN(n641) );
  NAND2_X1 U705 ( .A1(n642), .A2(n641), .ZN(n650) );
  NAND2_X1 U706 ( .A1(n650), .A2(G171), .ZN(n643) );
  NAND2_X1 U707 ( .A1(n644), .A2(n643), .ZN(n655) );
  NAND2_X1 U708 ( .A1(n513), .A2(G8), .ZN(n656) );
  NOR2_X1 U709 ( .A1(G1966), .A2(n656), .ZN(n669) );
  NOR2_X1 U710 ( .A1(n513), .A2(G2084), .ZN(n666) );
  NOR2_X1 U711 ( .A1(n669), .A2(n666), .ZN(n645) );
  XOR2_X1 U712 ( .A(n645), .B(KEYINPUT93), .Z(n646) );
  NAND2_X1 U713 ( .A1(G8), .A2(n646), .ZN(n648) );
  XNOR2_X1 U714 ( .A(KEYINPUT30), .B(KEYINPUT94), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X1 U716 ( .A1(G168), .A2(n649), .ZN(n652) );
  NOR2_X1 U717 ( .A1(G171), .A2(n650), .ZN(n651) );
  NOR2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U719 ( .A(KEYINPUT31), .B(n653), .Z(n654) );
  NAND2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n667) );
  NAND2_X1 U721 ( .A1(n667), .A2(G286), .ZN(n663) );
  NOR2_X1 U722 ( .A1(G1971), .A2(n656), .ZN(n659) );
  NOR2_X1 U723 ( .A1(n513), .A2(G2090), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U725 ( .A1(n660), .A2(G303), .ZN(n661) );
  XOR2_X1 U726 ( .A(KEYINPUT95), .B(n661), .Z(n662) );
  NAND2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U728 ( .A1(n664), .A2(G8), .ZN(n665) );
  XNOR2_X1 U729 ( .A(KEYINPUT32), .B(n665), .ZN(n673) );
  NAND2_X1 U730 ( .A1(G8), .A2(n666), .ZN(n671) );
  INV_X1 U731 ( .A(n667), .ZN(n668) );
  NOR2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n720) );
  NOR2_X1 U735 ( .A1(G1976), .A2(G288), .ZN(n679) );
  NOR2_X1 U736 ( .A1(G1971), .A2(G303), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n679), .A2(n674), .ZN(n920) );
  XNOR2_X1 U738 ( .A(KEYINPUT96), .B(n920), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n720), .A2(n675), .ZN(n676) );
  NAND2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n919) );
  NAND2_X1 U741 ( .A1(n676), .A2(n919), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n677), .A2(n656), .ZN(n678) );
  NOR2_X1 U743 ( .A1(n678), .A2(KEYINPUT33), .ZN(n716) );
  XOR2_X1 U744 ( .A(G1981), .B(G305), .Z(n903) );
  INV_X1 U745 ( .A(n903), .ZN(n682) );
  NAND2_X1 U746 ( .A1(n679), .A2(KEYINPUT33), .ZN(n680) );
  NOR2_X1 U747 ( .A1(n656), .A2(n680), .ZN(n681) );
  OR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n714) );
  NAND2_X1 U749 ( .A1(G160), .A2(G40), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n744) );
  NAND2_X1 U751 ( .A1(G104), .A2(n859), .ZN(n686) );
  NAND2_X1 U752 ( .A1(G140), .A2(n860), .ZN(n685) );
  NAND2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U754 ( .A(KEYINPUT34), .B(n687), .ZN(n692) );
  NAND2_X1 U755 ( .A1(G116), .A2(n863), .ZN(n689) );
  NAND2_X1 U756 ( .A1(G128), .A2(n865), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U758 ( .A(KEYINPUT35), .B(n690), .Z(n691) );
  NOR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U760 ( .A(KEYINPUT36), .B(n693), .ZN(n855) );
  XNOR2_X1 U761 ( .A(G2067), .B(KEYINPUT37), .ZN(n741) );
  NOR2_X1 U762 ( .A1(n855), .A2(n741), .ZN(n963) );
  NAND2_X1 U763 ( .A1(n744), .A2(n963), .ZN(n739) );
  XOR2_X1 U764 ( .A(KEYINPUT88), .B(KEYINPUT38), .Z(n695) );
  NAND2_X1 U765 ( .A1(G105), .A2(n859), .ZN(n694) );
  XNOR2_X1 U766 ( .A(n695), .B(n694), .ZN(n699) );
  NAND2_X1 U767 ( .A1(G117), .A2(n863), .ZN(n697) );
  NAND2_X1 U768 ( .A1(G129), .A2(n865), .ZN(n696) );
  NAND2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U770 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U771 ( .A1(n860), .A2(G141), .ZN(n700) );
  NAND2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n877) );
  NAND2_X1 U773 ( .A1(G1996), .A2(n877), .ZN(n710) );
  NAND2_X1 U774 ( .A1(G95), .A2(n859), .ZN(n703) );
  NAND2_X1 U775 ( .A1(G107), .A2(n863), .ZN(n702) );
  NAND2_X1 U776 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U777 ( .A1(G119), .A2(n865), .ZN(n704) );
  XNOR2_X1 U778 ( .A(KEYINPUT87), .B(n704), .ZN(n705) );
  NOR2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U780 ( .A1(n860), .A2(G131), .ZN(n707) );
  NAND2_X1 U781 ( .A1(n708), .A2(n707), .ZN(n871) );
  NAND2_X1 U782 ( .A1(G1991), .A2(n871), .ZN(n709) );
  NAND2_X1 U783 ( .A1(n710), .A2(n709), .ZN(n955) );
  NAND2_X1 U784 ( .A1(n744), .A2(n955), .ZN(n732) );
  NAND2_X1 U785 ( .A1(n739), .A2(n732), .ZN(n711) );
  XNOR2_X1 U786 ( .A(n711), .B(KEYINPUT89), .ZN(n713) );
  XNOR2_X1 U787 ( .A(G1986), .B(G290), .ZN(n908) );
  NAND2_X1 U788 ( .A1(n744), .A2(n908), .ZN(n712) );
  NAND2_X1 U789 ( .A1(n713), .A2(n712), .ZN(n717) );
  OR2_X1 U790 ( .A1(n714), .A2(n717), .ZN(n715) );
  NOR2_X1 U791 ( .A1(n716), .A2(n715), .ZN(n730) );
  INV_X1 U792 ( .A(n717), .ZN(n728) );
  NOR2_X1 U793 ( .A1(G2090), .A2(G303), .ZN(n718) );
  NAND2_X1 U794 ( .A1(G8), .A2(n718), .ZN(n719) );
  NAND2_X1 U795 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U796 ( .A1(n721), .A2(n656), .ZN(n726) );
  NOR2_X1 U797 ( .A1(G1981), .A2(G305), .ZN(n722) );
  XOR2_X1 U798 ( .A(n722), .B(KEYINPUT24), .Z(n723) );
  NOR2_X1 U799 ( .A1(n656), .A2(n723), .ZN(n724) );
  XOR2_X1 U800 ( .A(n724), .B(KEYINPUT90), .Z(n725) );
  NAND2_X1 U801 ( .A1(n726), .A2(n725), .ZN(n727) );
  AND2_X1 U802 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U803 ( .A(n731), .B(KEYINPUT97), .ZN(n747) );
  NOR2_X1 U804 ( .A1(G1996), .A2(n877), .ZN(n959) );
  INV_X1 U805 ( .A(n732), .ZN(n736) );
  NOR2_X1 U806 ( .A1(n871), .A2(G1991), .ZN(n733) );
  XNOR2_X1 U807 ( .A(n733), .B(KEYINPUT98), .ZN(n967) );
  NOR2_X1 U808 ( .A1(G1986), .A2(G290), .ZN(n734) );
  NOR2_X1 U809 ( .A1(n967), .A2(n734), .ZN(n735) );
  NOR2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U811 ( .A1(n959), .A2(n737), .ZN(n738) );
  XNOR2_X1 U812 ( .A(n738), .B(KEYINPUT39), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U814 ( .A1(n855), .A2(n741), .ZN(n954) );
  NAND2_X1 U815 ( .A1(n742), .A2(n954), .ZN(n743) );
  XOR2_X1 U816 ( .A(KEYINPUT99), .B(n743), .Z(n745) );
  NAND2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U819 ( .A(n748), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U820 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U821 ( .A(G57), .ZN(G237) );
  INV_X1 U822 ( .A(G132), .ZN(G219) );
  INV_X1 U823 ( .A(G82), .ZN(G220) );
  NAND2_X1 U824 ( .A1(G7), .A2(G661), .ZN(n749) );
  XNOR2_X1 U825 ( .A(n749), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U826 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n751) );
  INV_X1 U827 ( .A(G223), .ZN(n811) );
  NAND2_X1 U828 ( .A1(G567), .A2(n811), .ZN(n750) );
  XNOR2_X1 U829 ( .A(n751), .B(n750), .ZN(G234) );
  INV_X1 U830 ( .A(G860), .ZN(n773) );
  OR2_X1 U831 ( .A1(n906), .A2(n773), .ZN(G153) );
  INV_X1 U832 ( .A(G171), .ZN(G301) );
  INV_X1 U833 ( .A(n882), .ZN(n911) );
  NOR2_X1 U834 ( .A1(G868), .A2(n911), .ZN(n753) );
  INV_X1 U835 ( .A(G868), .ZN(n795) );
  NOR2_X1 U836 ( .A1(n795), .A2(G301), .ZN(n752) );
  NOR2_X1 U837 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U838 ( .A(KEYINPUT76), .B(n754), .ZN(G284) );
  INV_X1 U839 ( .A(n916), .ZN(G299) );
  XNOR2_X1 U840 ( .A(KEYINPUT78), .B(n795), .ZN(n755) );
  NOR2_X1 U841 ( .A1(G286), .A2(n755), .ZN(n757) );
  NOR2_X1 U842 ( .A1(G868), .A2(G299), .ZN(n756) );
  NOR2_X1 U843 ( .A1(n757), .A2(n756), .ZN(G297) );
  NAND2_X1 U844 ( .A1(n773), .A2(G559), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n758), .A2(n882), .ZN(n759) );
  XNOR2_X1 U846 ( .A(n759), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 U847 ( .A1(G559), .A2(n911), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n760), .A2(G868), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n906), .A2(n795), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(G282) );
  NAND2_X1 U851 ( .A1(G99), .A2(n859), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G111), .A2(n863), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n865), .A2(G123), .ZN(n765) );
  XOR2_X1 U855 ( .A(KEYINPUT18), .B(n765), .Z(n766) );
  NOR2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n860), .A2(G135), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n964) );
  XOR2_X1 U859 ( .A(n964), .B(G2096), .Z(n771) );
  XNOR2_X1 U860 ( .A(G2100), .B(KEYINPUT79), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(G156) );
  NAND2_X1 U862 ( .A1(G559), .A2(n882), .ZN(n772) );
  XOR2_X1 U863 ( .A(n906), .B(n772), .Z(n791) );
  NAND2_X1 U864 ( .A1(n773), .A2(n791), .ZN(n784) );
  NAND2_X1 U865 ( .A1(G55), .A2(n774), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G67), .A2(n775), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n783) );
  NAND2_X1 U868 ( .A1(G80), .A2(n778), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G93), .A2(n779), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n794) );
  XOR2_X1 U872 ( .A(n784), .B(n794), .Z(G145) );
  INV_X1 U873 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U874 ( .A(n916), .B(n794), .ZN(n789) );
  XNOR2_X1 U875 ( .A(G166), .B(G290), .ZN(n787) );
  XNOR2_X1 U876 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n785) );
  XNOR2_X1 U877 ( .A(n785), .B(G288), .ZN(n786) );
  XNOR2_X1 U878 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n789), .B(n788), .ZN(n790) );
  XNOR2_X1 U880 ( .A(n790), .B(G305), .ZN(n881) );
  XNOR2_X1 U881 ( .A(n791), .B(n881), .ZN(n792) );
  XNOR2_X1 U882 ( .A(KEYINPUT84), .B(n792), .ZN(n793) );
  NOR2_X1 U883 ( .A1(n795), .A2(n793), .ZN(n797) );
  AND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(G295) );
  NAND2_X1 U886 ( .A1(G2078), .A2(G2084), .ZN(n798) );
  XOR2_X1 U887 ( .A(KEYINPUT20), .B(n798), .Z(n799) );
  NAND2_X1 U888 ( .A1(G2090), .A2(n799), .ZN(n800) );
  XNOR2_X1 U889 ( .A(KEYINPUT21), .B(n800), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n801), .A2(G2072), .ZN(G158) );
  XOR2_X1 U891 ( .A(KEYINPUT85), .B(G44), .Z(n802) );
  XNOR2_X1 U892 ( .A(KEYINPUT3), .B(n802), .ZN(G218) );
  NOR2_X1 U893 ( .A1(G220), .A2(G219), .ZN(n803) );
  XOR2_X1 U894 ( .A(KEYINPUT22), .B(n803), .Z(n804) );
  NOR2_X1 U895 ( .A1(G218), .A2(n804), .ZN(n805) );
  NAND2_X1 U896 ( .A1(G96), .A2(n805), .ZN(n816) );
  NAND2_X1 U897 ( .A1(n816), .A2(G2106), .ZN(n809) );
  NAND2_X1 U898 ( .A1(G69), .A2(G120), .ZN(n806) );
  NOR2_X1 U899 ( .A1(G237), .A2(n806), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G108), .A2(n807), .ZN(n817) );
  NAND2_X1 U901 ( .A1(n817), .A2(G567), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n818) );
  NAND2_X1 U903 ( .A1(G483), .A2(G661), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n818), .A2(n810), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n813), .A2(G36), .ZN(G176) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n811), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n812) );
  NAND2_X1 U908 ( .A1(G661), .A2(n812), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G1), .A2(G3), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U911 ( .A(n815), .B(KEYINPUT100), .ZN(G188) );
  XNOR2_X1 U912 ( .A(G96), .B(KEYINPUT101), .ZN(G221) );
  INV_X1 U914 ( .A(G120), .ZN(G236) );
  INV_X1 U915 ( .A(G69), .ZN(G235) );
  NOR2_X1 U916 ( .A1(n817), .A2(n816), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  INV_X1 U918 ( .A(n818), .ZN(G319) );
  XOR2_X1 U919 ( .A(G2474), .B(G1961), .Z(n820) );
  XNOR2_X1 U920 ( .A(G1996), .B(G1991), .ZN(n819) );
  XNOR2_X1 U921 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U922 ( .A(n821), .B(KEYINPUT104), .Z(n823) );
  XNOR2_X1 U923 ( .A(G1976), .B(G1971), .ZN(n822) );
  XNOR2_X1 U924 ( .A(n823), .B(n822), .ZN(n827) );
  XOR2_X1 U925 ( .A(G1956), .B(G1966), .Z(n825) );
  XNOR2_X1 U926 ( .A(G1986), .B(G1981), .ZN(n824) );
  XNOR2_X1 U927 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U928 ( .A(n827), .B(n826), .Z(n829) );
  XNOR2_X1 U929 ( .A(KEYINPUT105), .B(KEYINPUT41), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n829), .B(n828), .ZN(G229) );
  XOR2_X1 U931 ( .A(KEYINPUT102), .B(G2678), .Z(n831) );
  XNOR2_X1 U932 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U934 ( .A(KEYINPUT42), .B(G2090), .Z(n833) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2072), .ZN(n832) );
  XNOR2_X1 U936 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U937 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U938 ( .A(G2096), .B(G2100), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n839) );
  XOR2_X1 U940 ( .A(G2078), .B(G2084), .Z(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(G227) );
  NAND2_X1 U942 ( .A1(G100), .A2(n859), .ZN(n841) );
  NAND2_X1 U943 ( .A1(G112), .A2(n863), .ZN(n840) );
  NAND2_X1 U944 ( .A1(n841), .A2(n840), .ZN(n846) );
  NAND2_X1 U945 ( .A1(G124), .A2(n865), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n842), .B(KEYINPUT44), .ZN(n844) );
  NAND2_X1 U947 ( .A1(n860), .A2(G136), .ZN(n843) );
  NAND2_X1 U948 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U949 ( .A1(n846), .A2(n845), .ZN(G162) );
  NAND2_X1 U950 ( .A1(G118), .A2(n863), .ZN(n848) );
  NAND2_X1 U951 ( .A1(G130), .A2(n865), .ZN(n847) );
  NAND2_X1 U952 ( .A1(n848), .A2(n847), .ZN(n854) );
  NAND2_X1 U953 ( .A1(G106), .A2(n859), .ZN(n850) );
  NAND2_X1 U954 ( .A1(G142), .A2(n860), .ZN(n849) );
  NAND2_X1 U955 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U956 ( .A(KEYINPUT45), .B(n851), .Z(n852) );
  XNOR2_X1 U957 ( .A(KEYINPUT106), .B(n852), .ZN(n853) );
  NOR2_X1 U958 ( .A1(n854), .A2(n853), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n857), .B(n964), .ZN(n858) );
  XNOR2_X1 U961 ( .A(G162), .B(n858), .ZN(n873) );
  NAND2_X1 U962 ( .A1(G103), .A2(n859), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G139), .A2(n860), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n870) );
  NAND2_X1 U965 ( .A1(n863), .A2(G115), .ZN(n864) );
  XOR2_X1 U966 ( .A(KEYINPUT107), .B(n864), .Z(n867) );
  NAND2_X1 U967 ( .A1(n865), .A2(G127), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U969 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n971) );
  XNOR2_X1 U971 ( .A(n871), .B(n971), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n879) );
  XOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n875) );
  XNOR2_X1 U974 ( .A(G160), .B(G164), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n880) );
  NOR2_X1 U978 ( .A1(G37), .A2(n880), .ZN(G395) );
  XNOR2_X1 U979 ( .A(n906), .B(n881), .ZN(n884) );
  XNOR2_X1 U980 ( .A(G171), .B(n882), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n885), .B(G286), .ZN(n886) );
  NOR2_X1 U983 ( .A1(G37), .A2(n886), .ZN(G397) );
  XOR2_X1 U984 ( .A(G2451), .B(G2430), .Z(n888) );
  XNOR2_X1 U985 ( .A(G2438), .B(G2443), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n894) );
  XOR2_X1 U987 ( .A(G2435), .B(G2454), .Z(n890) );
  XNOR2_X1 U988 ( .A(G1341), .B(G1348), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n892) );
  XOR2_X1 U990 ( .A(G2446), .B(G2427), .Z(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U992 ( .A(n894), .B(n893), .Z(n895) );
  NAND2_X1 U993 ( .A1(G14), .A2(n895), .ZN(n901) );
  NAND2_X1 U994 ( .A1(G319), .A2(n901), .ZN(n898) );
  NOR2_X1 U995 ( .A1(G229), .A2(G227), .ZN(n896) );
  XNOR2_X1 U996 ( .A(KEYINPUT49), .B(n896), .ZN(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n900) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n899) );
  NAND2_X1 U999 ( .A1(n900), .A2(n899), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(G108), .ZN(G238) );
  INV_X1 U1002 ( .A(n901), .ZN(G401) );
  XOR2_X1 U1003 ( .A(G1966), .B(G168), .Z(n902) );
  XNOR2_X1 U1004 ( .A(KEYINPUT117), .B(n902), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n905), .B(KEYINPUT57), .ZN(n915) );
  XNOR2_X1 U1007 ( .A(G171), .B(G1961), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(G1341), .B(n906), .ZN(n907) );
  NOR2_X1 U1009 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(G1348), .B(n911), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n925) );
  XNOR2_X1 U1014 ( .A(n916), .B(G1956), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(G1971), .A2(G303), .ZN(n917) );
  NAND2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1019 ( .A(KEYINPUT118), .B(n923), .Z(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n927) );
  XOR2_X1 U1021 ( .A(KEYINPUT56), .B(G16), .Z(n926) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n953) );
  XOR2_X1 U1023 ( .A(G2090), .B(G35), .Z(n931) );
  XNOR2_X1 U1024 ( .A(KEYINPUT54), .B(G34), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(n928), .B(KEYINPUT115), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n929), .B(G2084), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n948) );
  XNOR2_X1 U1028 ( .A(G27), .B(n932), .ZN(n940) );
  XOR2_X1 U1029 ( .A(G2067), .B(G26), .Z(n935) );
  XOR2_X1 U1030 ( .A(G32), .B(KEYINPUT112), .Z(n933) );
  XNOR2_X1 U1031 ( .A(G1996), .B(n933), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT111), .B(G2072), .Z(n936) );
  XNOR2_X1 U1034 ( .A(G33), .B(n936), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1037 ( .A(KEYINPUT113), .B(n941), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n942), .A2(G28), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(G25), .B(G1991), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(KEYINPUT53), .B(n945), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT114), .B(n946), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(KEYINPUT116), .B(n949), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n950), .A2(G29), .ZN(n951) );
  XOR2_X1 U1046 ( .A(KEYINPUT55), .B(n951), .Z(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n982) );
  INV_X1 U1048 ( .A(n954), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n978) );
  XNOR2_X1 U1050 ( .A(G2090), .B(G162), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(KEYINPUT109), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(KEYINPUT51), .B(KEYINPUT110), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n961), .B(n960), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n970) );
  XNOR2_X1 U1056 ( .A(G160), .B(G2084), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(n968), .B(KEYINPUT108), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n976) );
  XOR2_X1 U1061 ( .A(G2072), .B(n971), .Z(n973) );
  XOR2_X1 U1062 ( .A(G164), .B(G2078), .Z(n972) );
  NOR2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1064 ( .A(KEYINPUT50), .B(n974), .Z(n975) );
  NOR2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1066 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(KEYINPUT52), .B(n979), .ZN(n980) );
  NAND2_X1 U1068 ( .A1(n980), .A2(G29), .ZN(n981) );
  NAND2_X1 U1069 ( .A1(n982), .A2(n981), .ZN(n1016) );
  XOR2_X1 U1070 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n989) );
  XNOR2_X1 U1071 ( .A(G1986), .B(G24), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G22), .B(G1971), .ZN(n983) );
  NOR2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(G1976), .B(KEYINPUT121), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(n985), .B(G23), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(n989), .B(n988), .ZN(n990) );
  XOR2_X1 U1078 ( .A(KEYINPUT58), .B(n990), .Z(n1008) );
  XOR2_X1 U1079 ( .A(G1966), .B(G21), .Z(n993) );
  XNOR2_X1 U1080 ( .A(n991), .B(G5), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n1005) );
  XNOR2_X1 U1082 ( .A(KEYINPUT59), .B(G1348), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(n994), .B(G4), .ZN(n1001) );
  XOR2_X1 U1084 ( .A(G1341), .B(G19), .Z(n997) );
  XNOR2_X1 U1085 ( .A(n995), .B(G20), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G6), .B(G1981), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(KEYINPUT119), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT120), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1009), .B(KEYINPUT61), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(n1011), .B(n1010), .Z(n1012) );
  NOR2_X1 U1098 ( .A1(G16), .A2(n1012), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT126), .B(n1013), .Z(n1014) );
  NAND2_X1 U1100 ( .A1(G11), .A2(n1014), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(n1017), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

