//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n559,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G567), .B1(new_n456), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G101), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n460), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n468), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n466), .B1(new_n477), .B2(G2105), .ZN(G160));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n473), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n460), .B1(new_n471), .B2(new_n472), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT70), .ZN(new_n490));
  AOI21_X1  g065(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n491));
  AOI211_X1 g066(.A(new_n481), .B(new_n490), .C1(G136), .C2(new_n491), .ZN(G162));
  OAI211_X1 g067(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n473), .A2(new_n495), .A3(G138), .A4(new_n460), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n460), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT71), .A4(G2104), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n501), .A2(new_n505), .B1(new_n485), .B2(G126), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT73), .B1(new_n509), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT5), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(new_n513), .B1(new_n509), .B2(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OR3_X1    g091(.A1(new_n515), .A2(KEYINPUT74), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT74), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT72), .A3(G50), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n514), .A2(new_n519), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n522), .A2(new_n525), .B1(new_n526), .B2(G88), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n517), .A2(new_n518), .A3(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  XOR2_X1   g104(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n521), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n526), .A2(G89), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(G168));
  AND2_X1   g112(.A1(new_n514), .A2(G64), .ZN(new_n538));
  AND2_X1   g113(.A1(G77), .A2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(G651), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g117(.A(KEYINPUT76), .B(G651), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n526), .A2(G90), .B1(G52), .B2(new_n521), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AND2_X1   g121(.A1(new_n514), .A2(G56), .ZN(new_n547));
  AND2_X1   g122(.A1(G68), .A2(G543), .ZN(new_n548));
  OAI21_X1  g123(.A(G651), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n526), .A2(G81), .B1(G43), .B2(new_n521), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G860), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT78), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g133(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n559));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  AND2_X1   g137(.A1(new_n526), .A2(G91), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  OAI21_X1  g139(.A(G53), .B1(new_n564), .B2(KEYINPUT80), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n520), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(KEYINPUT80), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NOR3_X1   g144(.A1(new_n563), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n514), .A2(G65), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT81), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n516), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  NAND2_X1  g152(.A1(new_n521), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n514), .A2(G87), .A3(new_n519), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n510), .A2(new_n513), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n509), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(G48), .B2(new_n521), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n526), .A2(G86), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n516), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n514), .A2(new_n519), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n593), .A2(new_n594), .B1(new_n595), .B2(new_n520), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n592), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n526), .A2(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT10), .Z(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n585), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n521), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G321));
  MUX2_X1   g183(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g184(.A(G280), .B(KEYINPUT82), .ZN(G297));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n606), .B1(new_n611), .B2(G860), .ZN(G148));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n611), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(new_n615));
  INV_X1    g190(.A(new_n554), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(G868), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n614), .A2(new_n613), .A3(G868), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g195(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n621));
  NOR3_X1   g196(.A1(new_n469), .A2(new_n470), .A3(G2105), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G2100), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT85), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n624), .A2(G2100), .ZN(new_n627));
  INV_X1    g202(.A(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n488), .A2(G123), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT86), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G111), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n630), .A2(new_n631), .B1(new_n633), .B2(G2105), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n632), .A2(new_n634), .B1(new_n491), .B2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n627), .B1(new_n628), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n626), .B(new_n638), .C1(new_n628), .C2(new_n637), .ZN(G156));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n643), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT87), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  NOR2_X1   g233(.A1(G2072), .A2(G2078), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n442), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n657), .A2(new_n660), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(KEYINPUT17), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n664), .B(new_n658), .C1(new_n657), .C2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT89), .ZN(new_n667));
  INV_X1    g242(.A(new_n657), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n658), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT90), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT20), .Z(new_n682));
  OR2_X1    g257(.A1(new_n675), .A2(new_n677), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(new_n680), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n680), .A3(new_n678), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT91), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n692), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  OR3_X1    g271(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n693), .B2(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  MUX2_X1   g274(.A(G6), .B(G305), .S(G16), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT94), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(G288), .A2(KEYINPUT95), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n578), .A2(new_n579), .A3(new_n705), .A4(new_n580), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G23), .B(new_n707), .S(G16), .Z(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G22), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G166), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1971), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n703), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n491), .A2(G131), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n460), .A2(G107), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n721));
  INV_X1    g296(.A(G119), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n719), .B1(new_n720), .B2(new_n721), .C1(new_n487), .C2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT92), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(new_n717), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT93), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n727), .A2(new_n729), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G24), .ZN(new_n733));
  INV_X1    g308(.A(G290), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1986), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n730), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n716), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT36), .ZN(new_n740));
  NAND2_X1  g315(.A1(G299), .A2(G16), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n732), .A2(G20), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT102), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT23), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n717), .A2(G35), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G162), .B2(new_n717), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n746), .B1(new_n749), .B2(G2090), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT103), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G19), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n616), .B2(G16), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(G1341), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n717), .A2(G32), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n488), .A2(G129), .ZN(new_n756));
  INV_X1    g331(.A(G105), .ZN(new_n757));
  OR3_X1    g332(.A1(new_n465), .A2(KEYINPUT100), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(KEYINPUT100), .B1(new_n465), .B2(new_n757), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT26), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n758), .A2(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n756), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n491), .A2(G141), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT99), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n755), .B1(new_n769), .B2(new_n717), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT101), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT27), .B(G1996), .Z(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G1961), .ZN(new_n774));
  NOR2_X1   g349(.A1(G171), .A2(new_n732), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G5), .B2(new_n732), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n754), .B(new_n773), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n749), .A2(G2090), .ZN(new_n778));
  OAI22_X1  g353(.A1(new_n776), .A2(new_n774), .B1(G1341), .B2(new_n753), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n717), .A2(G26), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT28), .Z(new_n781));
  OR2_X1    g356(.A1(G104), .A2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n782), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT96), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G140), .B2(new_n491), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n488), .A2(G128), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n781), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT97), .B(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G160), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT24), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n792), .A2(G34), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n717), .B1(new_n792), .B2(G34), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n791), .A2(new_n717), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2084), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n717), .A2(G33), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n473), .A2(G127), .ZN(new_n798));
  NAND2_X1  g373(.A1(G115), .A2(G2104), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n460), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n491), .A2(G139), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT25), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n800), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT98), .Z(new_n806));
  AOI21_X1  g381(.A(new_n797), .B1(new_n806), .B2(G29), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n790), .B(new_n796), .C1(G2072), .C2(new_n808), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n779), .B(new_n809), .C1(new_n772), .C2(new_n771), .ZN(new_n810));
  NOR2_X1   g385(.A1(G4), .A2(G16), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n606), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1348), .ZN(new_n813));
  NOR2_X1   g388(.A1(G164), .A2(new_n717), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G27), .B2(new_n717), .ZN(new_n815));
  INV_X1    g390(.A(G2078), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT31), .B(G11), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT30), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(G28), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n717), .B1(new_n819), .B2(G28), .ZN(new_n821));
  OAI221_X1 g396(.A(new_n818), .B1(new_n820), .B2(new_n821), .C1(new_n636), .C2(new_n717), .ZN(new_n822));
  NOR2_X1   g397(.A1(G168), .A2(new_n732), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n732), .B2(G21), .ZN(new_n824));
  INV_X1    g399(.A(G1966), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G2072), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n807), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n815), .A2(new_n816), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n824), .B2(new_n825), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n813), .A2(new_n817), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n777), .A2(new_n778), .A3(new_n810), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n751), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n740), .A2(new_n833), .ZN(G150));
  INV_X1    g409(.A(G150), .ZN(G311));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n593), .A2(new_n836), .B1(new_n837), .B2(new_n520), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT104), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(new_n516), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n843), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n616), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n843), .B(KEYINPUT105), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n554), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n605), .A2(new_n611), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n851), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n555), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n636), .B(new_n791), .ZN(new_n859));
  XOR2_X1   g434(.A(G162), .B(new_n859), .Z(new_n860));
  XOR2_X1   g435(.A(new_n806), .B(new_n768), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n723), .B(KEYINPUT106), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n491), .A2(G142), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  INV_X1    g440(.A(G118), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n865), .B1(new_n866), .B2(G2105), .ZN(new_n867));
  AOI211_X1 g442(.A(new_n864), .B(new_n867), .C1(new_n488), .C2(G130), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n862), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n861), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n787), .B(new_n507), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n623), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n870), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n860), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n875), .ZN(new_n877));
  INV_X1    g452(.A(new_n860), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n878), .A3(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g457(.A(new_n734), .B(new_n707), .ZN(new_n883));
  XNOR2_X1  g458(.A(G303), .B(G305), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(KEYINPUT107), .B2(KEYINPUT42), .ZN(new_n887));
  NAND2_X1  g462(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n887), .B(new_n888), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n851), .B(new_n614), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n605), .B(G299), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n891), .B(KEYINPUT41), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n889), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n889), .B1(new_n893), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(G868), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n843), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n899), .B1(G868), .B2(new_n900), .ZN(G295));
  OAI21_X1  g476(.A(new_n899), .B1(G868), .B2(new_n900), .ZN(G331));
  AOI21_X1  g477(.A(G301), .B1(KEYINPUT108), .B2(G168), .ZN(new_n903));
  OR2_X1    g478(.A1(G168), .A2(KEYINPUT108), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n851), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n903), .B(new_n904), .Z(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n848), .A3(new_n850), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n892), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n894), .A2(new_n906), .A3(new_n908), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n912), .B2(new_n885), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n886), .A3(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT44), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n885), .ZN(new_n921));
  AND4_X1   g496(.A1(new_n917), .A2(new_n921), .A3(new_n880), .A4(new_n914), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n917), .B1(new_n913), .B2(new_n914), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n924), .ZN(G397));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n507), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT45), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n928), .B2(new_n927), .ZN(new_n930));
  NAND2_X1  g505(.A1(G160), .A2(G40), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G1996), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n768), .B(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G2067), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n787), .B(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n723), .B(new_n728), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(G290), .B(G1986), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n932), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G8), .ZN(new_n942));
  INV_X1    g517(.A(G40), .ZN(new_n943));
  AOI211_X1 g518(.A(new_n943), .B(new_n466), .C1(new_n477), .C2(G2105), .ZN(new_n944));
  AOI21_X1  g519(.A(G1384), .B1(new_n497), .B2(new_n506), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G288), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(G1976), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n704), .A2(G1976), .A3(new_n706), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n946), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n946), .A2(new_n952), .A3(new_n953), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n950), .A3(new_n949), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n587), .A2(G651), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n521), .A2(G48), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT113), .B(G86), .Z(new_n961));
  OR2_X1    g536(.A1(new_n593), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(G1981), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n588), .A2(new_n687), .A3(new_n589), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n965), .A3(KEYINPUT49), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n966), .A2(new_n946), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n965), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT114), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n971), .B(KEYINPUT49), .C1(new_n964), .C2(new_n965), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n967), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n958), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n927), .A2(KEYINPUT110), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n945), .B2(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n945), .A2(KEYINPUT45), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n976), .A2(new_n978), .A3(new_n944), .A4(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n979), .A2(new_n944), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n983), .A2(KEYINPUT111), .A3(new_n976), .A4(new_n978), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n984), .A3(new_n713), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n945), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n988), .B2(new_n931), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n944), .B(KEYINPUT116), .C1(new_n987), .C2(new_n945), .ZN(new_n990));
  INV_X1    g565(.A(G2090), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n945), .A2(new_n987), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n985), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G8), .ZN(new_n995));
  AND3_X1   g570(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n974), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n979), .A2(new_n944), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n945), .A2(KEYINPUT45), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n825), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n927), .A2(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(G2084), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n944), .A4(new_n992), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(G168), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  AOI21_X1  g582(.A(G168), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT51), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1010), .A3(G8), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1003), .A2(new_n991), .A3(new_n944), .A4(new_n992), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n942), .B1(new_n985), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n998), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1009), .A2(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n1016));
  OAI211_X1 g591(.A(G40), .B(G160), .C1(new_n945), .C2(new_n987), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n945), .A2(new_n987), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1003), .A2(KEYINPUT119), .A3(new_n944), .A4(new_n992), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT123), .B(G1961), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT124), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1019), .A2(KEYINPUT124), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n930), .A2(KEYINPUT53), .A3(new_n816), .A4(new_n983), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n982), .A2(new_n984), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n816), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G301), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1001), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n983), .A2(KEYINPUT53), .A3(new_n816), .A4(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1022), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(G2078), .B1(new_n982), .B2(new_n984), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1036), .B(G301), .C1(KEYINPUT53), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT54), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n999), .B(new_n1015), .C1(new_n1033), .C2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT53), .B1(new_n1029), .B2(new_n816), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1027), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G301), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1036), .ZN(new_n1044));
  OAI21_X1  g619(.A(G171), .B1(new_n1044), .B2(new_n1041), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT54), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT125), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n999), .A2(new_n1015), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1027), .A2(new_n1041), .A3(G171), .ZN(new_n1050));
  AOI21_X1  g625(.A(G301), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT125), .ZN(new_n1053));
  OAI211_X1 g628(.A(KEYINPUT54), .B(new_n1038), .C1(new_n1042), .C2(G301), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1048), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1047), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT56), .B(G2072), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n980), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1956), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n992), .B1(new_n1017), .B2(new_n986), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT116), .B1(new_n1003), .B2(new_n944), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT117), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n989), .A2(new_n992), .A3(new_n990), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n1060), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1059), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(G299), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n570), .A2(new_n1070), .A3(new_n1071), .A4(new_n575), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1068), .A2(new_n1076), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1059), .B(new_n1075), .C1(new_n1064), .C2(new_n1067), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n931), .A2(new_n927), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT58), .B(G1341), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n980), .A2(G1996), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n616), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(KEYINPUT120), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1084), .B(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1019), .A2(new_n1088), .A3(new_n1020), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1081), .A2(new_n935), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n606), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n605), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT60), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n605), .A2(KEYINPUT60), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1087), .B(new_n1094), .C1(new_n1091), .C2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1080), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1078), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1068), .A2(KEYINPUT121), .A3(new_n1076), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1059), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1065), .A2(new_n1066), .A3(new_n1060), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1066), .B1(new_n1065), .B2(new_n1060), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1100), .B1(new_n1104), .B2(new_n1075), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1098), .B1(new_n1099), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT122), .B1(new_n1106), .B2(new_n1079), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT121), .B1(new_n1068), .B2(new_n1076), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1100), .A3(new_n1075), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1078), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1110), .A2(new_n1111), .A3(KEYINPUT61), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1097), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1077), .B1(new_n1098), .B2(new_n1093), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1056), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(G8), .A3(G168), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n974), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1119));
  INV_X1    g694(.A(G1976), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n973), .A2(new_n1120), .A3(new_n947), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n965), .B(KEYINPUT115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1119), .A2(KEYINPUT63), .B1(new_n946), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(KEYINPUT63), .B2(new_n1117), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1045), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n999), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n941), .B1(new_n1115), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n932), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n769), .B2(new_n936), .ZN(new_n1136));
  OR3_X1    g711(.A1(new_n1135), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT46), .B1(new_n1135), .B2(G1996), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n1139), .B(KEYINPUT47), .Z(new_n1140));
  NAND3_X1  g715(.A1(new_n937), .A2(new_n728), .A3(new_n725), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n785), .A2(new_n935), .A3(new_n786), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n932), .A2(new_n689), .A3(new_n734), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1145), .A2(KEYINPUT48), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n939), .A2(new_n932), .B1(KEYINPUT48), .B2(new_n1145), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1143), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1140), .A2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT126), .Z(new_n1150));
  NAND2_X1  g725(.A1(new_n1134), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g726(.A(G319), .B1(new_n653), .B2(new_n654), .ZN(new_n1153));
  NOR2_X1   g727(.A1(G227), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g728(.A1(new_n697), .A2(new_n881), .A3(new_n698), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g729(.A(new_n1155), .B1(new_n916), .B2(new_n918), .ZN(G308));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1157));
  OAI21_X1  g731(.A(new_n1157), .B1(new_n923), .B2(new_n922), .ZN(G225));
endmodule


