//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n752, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  XOR2_X1   g002(.A(KEYINPUT84), .B(G36gat), .Z(new_n204));
  AOI22_X1  g003(.A1(new_n202), .A2(new_n203), .B1(new_n204), .B2(G29gat), .ZN(new_n205));
  OR3_X1    g004(.A1(KEYINPUT83), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT83), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(KEYINPUT14), .A3(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n208), .C1(KEYINPUT14), .C2(new_n207), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n203), .A2(new_n202), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT17), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT85), .ZN(new_n217));
  INV_X1    g016(.A(G1gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n213), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n215), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n214), .A2(new_n223), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT18), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n214), .B(new_n223), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n227), .B(KEYINPUT13), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n229), .A2(new_n230), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G169gat), .B(G197gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT82), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G113gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n240));
  INV_X1    g039(.A(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n239), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT12), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n231), .A2(new_n234), .A3(new_n235), .A4(new_n244), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT76), .B(KEYINPUT31), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT70), .B(G197gat), .ZN(new_n253));
  INV_X1    g052(.A(G204gat), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n254), .ZN(new_n256));
  XOR2_X1   g055(.A(KEYINPUT71), .B(G218gat), .Z(new_n257));
  INV_X1    g056(.A(G211gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n255), .B(new_n256), .C1(new_n259), .C2(KEYINPUT22), .ZN(new_n260));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n252), .B1(new_n262), .B2(KEYINPUT29), .ZN(new_n263));
  XOR2_X1   g062(.A(G141gat), .B(G148gat), .Z(new_n264));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265));
  INV_X1    g064(.A(G155gat), .ZN(new_n266));
  INV_X1    g065(.A(G162gat), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT2), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G155gat), .B(G162gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n262), .B(KEYINPUT72), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(KEYINPUT29), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n273), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G22gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G228gat), .A2(G233gat), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n281), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT78), .ZN(new_n286));
  XNOR2_X1  g085(.A(G78gat), .B(G106gat), .ZN(new_n287));
  INV_X1    g086(.A(G50gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT78), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n282), .A2(new_n283), .A3(new_n291), .A4(new_n284), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n286), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n290), .B1(new_n286), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n251), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n286), .A2(new_n292), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n289), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n286), .A2(new_n290), .A3(new_n292), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n250), .A3(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G127gat), .B(G134gat), .Z(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(KEYINPUT1), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(G113gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(G120gat), .ZN(new_n304));
  INV_X1    g103(.A(G120gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n304), .B(new_n306), .C1(G113gat), .C2(new_n305), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G113gat), .B(G120gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n300), .B1(new_n309), .B2(KEYINPUT1), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n271), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT4), .ZN(new_n313));
  INV_X1    g112(.A(new_n311), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n271), .B2(new_n252), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n276), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT5), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n272), .A2(new_n314), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n322), .A2(new_n312), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT5), .B1(new_n323), .B2(new_n317), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n321), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G1gat), .B(G29gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT0), .ZN(new_n327));
  XOR2_X1   g126(.A(G57gat), .B(G85gat), .Z(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n325), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n325), .A2(new_n330), .ZN(new_n333));
  INV_X1    g132(.A(new_n331), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n325), .A2(new_n330), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(KEYINPUT29), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT65), .B(G190gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT27), .B(G183gat), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(KEYINPUT67), .Z(new_n345));
  AND2_X1   g144(.A1(new_n342), .A2(KEYINPUT28), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G169gat), .ZN(new_n348));
  INV_X1    g147(.A(G176gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT26), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT26), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI221_X1 g155(.A(new_n350), .B1(new_n351), .B2(new_n352), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT24), .B1(new_n351), .B2(new_n352), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(G183gat), .A3(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(G183gat), .B2(G190gat), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT23), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT23), .B1(new_n348), .B2(new_n349), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n364), .A2(new_n365), .A3(new_n356), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT25), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n362), .B1(G183gat), .B2(new_n341), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n366), .A2(KEYINPUT25), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n340), .B1(new_n358), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT66), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n370), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n358), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n339), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n275), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n374), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n358), .A2(new_n370), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n377), .A2(new_n340), .B1(new_n339), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n376), .B1(new_n379), .B2(new_n275), .ZN(new_n380));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  OR2_X1    g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n384), .B(KEYINPUT73), .Z(new_n385));
  NAND2_X1  g184(.A1(new_n380), .A2(new_n383), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT30), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n338), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n377), .B(new_n311), .ZN(new_n390));
  NAND2_X1  g189(.A1(G227gat), .A2(G233gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n391), .B(KEYINPUT64), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n394), .A2(KEYINPUT34), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(KEYINPUT34), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n377), .B(new_n314), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT33), .B1(new_n397), .B2(new_n392), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT69), .B(G71gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(G99gat), .ZN(new_n400));
  XOR2_X1   g199(.A(G15gat), .B(G43gat), .Z(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n395), .B(new_n396), .C1(new_n398), .C2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n398), .A2(new_n403), .ZN(new_n405));
  INV_X1    g204(.A(new_n396), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n394), .A2(KEYINPUT34), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n397), .A2(new_n392), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT32), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n404), .B2(new_n408), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n295), .A2(new_n299), .A3(new_n389), .A4(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT35), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT37), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n383), .B1(new_n380), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n379), .B2(new_n275), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n375), .A2(new_n371), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n274), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT38), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n386), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n337), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n419), .B1(new_n418), .B2(new_n380), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT38), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n316), .A2(new_n318), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT79), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT39), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n330), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n323), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT39), .B1(new_n433), .B2(new_n318), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(KEYINPUT80), .A2(KEYINPUT40), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n333), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n435), .A2(new_n436), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n426), .A2(new_n428), .B1(new_n440), .B2(new_n388), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n299), .A3(new_n295), .ZN(new_n442));
  INV_X1    g241(.A(new_n414), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT36), .B1(new_n443), .B2(new_n412), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n413), .A2(new_n414), .A3(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n295), .A2(new_n299), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n442), .B(new_n447), .C1(new_n448), .C2(new_n389), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n249), .B1(new_n417), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT7), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT87), .ZN(new_n454));
  AND2_X1   g253(.A1(G85gat), .A2(G92gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n457));
  INV_X1    g256(.A(G92gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G85gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(KEYINPUT88), .A2(G92gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G99gat), .ZN(new_n463));
  INV_X1    g262(.A(G106gat), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT8), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(KEYINPUT87), .A3(new_n453), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n456), .A2(new_n462), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G99gat), .B(G106gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n465), .A2(new_n467), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n472), .A2(new_n469), .A3(new_n456), .A4(new_n462), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n215), .A2(new_n225), .A3(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(G190gat), .B(G218gat), .Z(new_n476));
  INV_X1    g275(.A(KEYINPUT41), .ZN(new_n477));
  NAND2_X1  g276(.A1(G232gat), .A2(G233gat), .ZN(new_n478));
  OAI22_X1  g277(.A1(new_n476), .A2(KEYINPUT89), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n474), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n213), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(KEYINPUT89), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n482), .B(new_n483), .Z(new_n484));
  XOR2_X1   g283(.A(G134gat), .B(G162gat), .Z(new_n485));
  NAND2_X1  g284(.A1(new_n478), .A2(new_n477), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n488), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT21), .ZN(new_n492));
  AND2_X1   g291(.A1(G71gat), .A2(G78gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(G71gat), .A2(G78gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G57gat), .B(G64gat), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G57gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G64gat), .ZN(new_n500));
  INV_X1    g299(.A(G64gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(G57gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G71gat), .B(G78gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n497), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n223), .B1(new_n492), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n492), .ZN(new_n511));
  NAND2_X1  g310(.A1(G231gat), .A2(G233gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(G127gat), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n510), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G155gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(G183gat), .B(G211gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n515), .B(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n491), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G230gat), .A2(G233gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT10), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n507), .A2(new_n471), .A3(new_n473), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n471), .A2(new_n473), .B1(new_n498), .B2(new_n506), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT90), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT90), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n474), .A2(new_n508), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n523), .B(new_n524), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(KEYINPUT10), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n474), .A2(new_n508), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n507), .A2(new_n471), .A3(new_n473), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n480), .A2(KEYINPUT90), .A3(new_n507), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT10), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(new_n523), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n522), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n536), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(new_n522), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT92), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G120gat), .B(G148gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G176gat), .B(G204gat), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  XOR2_X1   g346(.A(new_n547), .B(KEYINPUT93), .Z(new_n548));
  NOR2_X1   g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT94), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n547), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n540), .A2(new_n543), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n549), .A2(new_n550), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n450), .A2(new_n521), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(new_n337), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(new_n218), .ZN(G1324gat));
  INV_X1    g359(.A(new_n388), .ZN(new_n561));
  OR3_X1    g360(.A1(new_n558), .A2(KEYINPUT96), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT96), .B1(new_n558), .B2(new_n561), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(G8gat), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n558), .A2(new_n561), .ZN(new_n565));
  XOR2_X1   g364(.A(KEYINPUT16), .B(G8gat), .Z(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(KEYINPUT42), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n562), .B2(new_n563), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT95), .B(KEYINPUT42), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n564), .B(new_n567), .C1(new_n569), .C2(new_n570), .ZN(G1325gat));
  OAI21_X1  g370(.A(G15gat), .B1(new_n558), .B2(new_n447), .ZN(new_n572));
  INV_X1    g371(.A(new_n415), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n573), .A2(G15gat), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n572), .B1(new_n558), .B2(new_n574), .ZN(G1326gat));
  NAND2_X1  g374(.A1(new_n295), .A2(new_n299), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n450), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n521), .A2(new_n557), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT43), .B(G22gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(G1327gat));
  INV_X1    g380(.A(new_n491), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n417), .B2(new_n449), .ZN(new_n583));
  INV_X1    g382(.A(new_n557), .ZN(new_n584));
  INV_X1    g383(.A(new_n520), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(new_n249), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n589), .A2(G29gat), .A3(new_n337), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT45), .Z(new_n591));
  INV_X1    g390(.A(new_n588), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n416), .A2(KEYINPUT35), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n416), .A2(KEYINPUT35), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n449), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT97), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n417), .A2(new_n597), .A3(new_n449), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n582), .A2(KEYINPUT44), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n491), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT44), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n592), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(G29gat), .B1(new_n604), .B2(new_n337), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n591), .A2(new_n605), .ZN(G1328gat));
  NOR3_X1   g405(.A1(new_n589), .A2(new_n204), .A3(new_n561), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT46), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n204), .B1(new_n604), .B2(new_n561), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(G1329gat));
  INV_X1    g409(.A(G43gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n589), .B2(new_n573), .ZN(new_n612));
  INV_X1    g411(.A(new_n447), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(G43gat), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n612), .B1(new_n604), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT47), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT47), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n617), .B(new_n612), .C1(new_n604), .C2(new_n614), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(G1330gat));
  INV_X1    g418(.A(KEYINPUT48), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n288), .B1(new_n603), .B2(new_n576), .ZN(new_n621));
  NOR4_X1   g420(.A1(new_n577), .A2(G50gat), .A3(new_n582), .A4(new_n587), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  AOI211_X1 g423(.A(new_n448), .B(new_n592), .C1(new_n600), .C2(new_n602), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n624), .B(KEYINPUT48), .C1(new_n625), .C2(new_n288), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(G1331gat));
  NAND3_X1  g426(.A1(new_n521), .A2(new_n249), .A3(new_n584), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT98), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n596), .A2(new_n598), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(new_n337), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT99), .B(G57gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(G1332gat));
  AOI21_X1  g432(.A(new_n561), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n596), .A2(new_n598), .A3(new_n629), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT100), .ZN(new_n636));
  OR2_X1    g435(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1333gat));
  OAI21_X1  g437(.A(G71gat), .B1(new_n630), .B2(new_n447), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n573), .A2(G71gat), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n630), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT50), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1334gat));
  NOR2_X1   g442(.A1(new_n630), .A2(new_n448), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(G78gat), .Z(G1335gat));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n585), .A2(new_n248), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n584), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n648), .B1(new_n600), .B2(new_n602), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n460), .B1(new_n649), .B2(new_n338), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n595), .A2(new_n491), .A3(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(KEYINPUT101), .A2(KEYINPUT51), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT51), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n583), .A2(new_n653), .A3(new_n654), .A4(new_n647), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n337), .A2(new_n557), .A3(G85gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT102), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n646), .B1(new_n650), .B2(new_n661), .ZN(new_n662));
  AOI211_X1 g461(.A(new_n337), .B(new_n648), .C1(new_n600), .C2(new_n602), .ZN(new_n663));
  OAI211_X1 g462(.A(KEYINPUT103), .B(new_n660), .C1(new_n663), .C2(new_n460), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(G1336gat));
  AND2_X1   g464(.A1(new_n459), .A2(new_n461), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n649), .B2(new_n388), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n651), .A2(new_n668), .A3(KEYINPUT51), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT51), .B1(new_n651), .B2(new_n668), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n561), .A2(G92gat), .A3(new_n557), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT52), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT52), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n657), .A3(new_n671), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n561), .B(new_n648), .C1(new_n600), .C2(new_n602), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n675), .B(new_n676), .C1(new_n677), .C2(new_n666), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n678), .ZN(G1337gat));
  NOR2_X1   g478(.A1(new_n573), .A2(G99gat), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n656), .A2(new_n657), .A3(new_n584), .A4(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n649), .A2(new_n613), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n463), .ZN(G1338gat));
  XOR2_X1   g482(.A(KEYINPUT105), .B(G106gat), .Z(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n649), .B2(new_n576), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n448), .A2(G106gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n584), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n669), .A2(new_n670), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT53), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT53), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n656), .A2(new_n657), .A3(new_n584), .A4(new_n686), .ZN(new_n691));
  AOI211_X1 g490(.A(new_n448), .B(new_n648), .C1(new_n600), .C2(new_n602), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n684), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n693), .ZN(G1339gat));
  AOI22_X1  g493(.A1(new_n537), .A2(new_n523), .B1(KEYINPUT10), .B2(new_n525), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n541), .A2(new_n524), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT91), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT54), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n699), .A3(new_n522), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(KEYINPUT55), .A3(new_n552), .ZN(new_n701));
  INV_X1    g500(.A(new_n522), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n695), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n539), .A2(KEYINPUT54), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT106), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n539), .A2(new_n703), .A3(new_n706), .A4(KEYINPUT54), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n701), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT107), .B1(new_n708), .B2(new_n553), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n700), .A2(KEYINPUT55), .A3(new_n552), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n699), .B1(new_n698), .B2(new_n522), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n706), .B1(new_n711), .B2(new_n703), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n706), .A2(new_n539), .A3(KEYINPUT54), .A4(new_n703), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n554), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n709), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n552), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n705), .B2(new_n707), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT108), .B1(new_n719), .B2(KEYINPUT55), .ZN(new_n720));
  OR3_X1    g519(.A1(new_n719), .A2(KEYINPUT108), .A3(KEYINPUT55), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n717), .A2(new_n248), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n232), .A2(new_n233), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n227), .B1(new_n226), .B2(new_n228), .ZN(new_n724));
  OAI211_X1 g523(.A(KEYINPUT109), .B(new_n243), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n243), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n247), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n555), .B2(new_n556), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n722), .A2(KEYINPUT110), .A3(new_n730), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n582), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n721), .A2(new_n720), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n736), .A2(new_n491), .A3(new_n717), .A4(new_n729), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n585), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n578), .A2(new_n248), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n740), .A2(new_n576), .A3(new_n573), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n388), .A2(new_n337), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(G113gat), .A3(new_n248), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n303), .B1(new_n743), .B2(new_n249), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1340gat));
  NOR2_X1   g548(.A1(new_n743), .A2(new_n557), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n305), .ZN(G1341gat));
  NAND2_X1  g550(.A1(new_n744), .A2(new_n585), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G127gat), .ZN(G1342gat));
  AOI211_X1 g552(.A(new_n582), .B(new_n743), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1343gat));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n448), .B2(new_n613), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n576), .A2(KEYINPUT115), .A3(new_n447), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n561), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n740), .B2(new_n337), .ZN(new_n762));
  OAI211_X1 g561(.A(KEYINPUT114), .B(new_n338), .C1(new_n738), .C2(new_n739), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n249), .A2(G141gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n768), .B(new_n576), .C1(new_n738), .C2(new_n739), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n742), .B1(new_n444), .B2(new_n446), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT112), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n772), .B(new_n742), .C1(new_n444), .C2(new_n446), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n248), .B1(KEYINPUT55), .B2(new_n719), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n714), .A2(new_n554), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n730), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n582), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n585), .B1(new_n778), .B2(new_n737), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n576), .B1(new_n779), .B2(new_n739), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n774), .B1(KEYINPUT57), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n769), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G141gat), .B1(new_n782), .B2(new_n249), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n781), .A3(KEYINPUT113), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n248), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G141gat), .ZN(new_n790));
  AOI211_X1 g589(.A(new_n785), .B(new_n767), .C1(new_n790), .C2(new_n766), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n769), .A2(KEYINPUT113), .A3(new_n781), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT113), .B1(new_n769), .B2(new_n781), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(new_n249), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n766), .B1(new_n794), .B2(new_n241), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT116), .B1(new_n795), .B2(KEYINPUT58), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n784), .B1(new_n791), .B2(new_n796), .ZN(G1344gat));
  INV_X1    g596(.A(G148gat), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n792), .A2(new_n793), .ZN(new_n799));
  AOI211_X1 g598(.A(KEYINPUT59), .B(new_n798), .C1(new_n799), .C2(new_n584), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n764), .A2(new_n798), .A3(new_n584), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n739), .B(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n779), .ZN(new_n806));
  AOI211_X1 g605(.A(KEYINPUT57), .B(new_n448), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n738), .A2(new_n739), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n576), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(KEYINPUT57), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n774), .A2(new_n557), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n798), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT117), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n802), .B(new_n803), .C1(new_n800), .C2(new_n814), .ZN(G1345gat));
  NAND2_X1  g614(.A1(new_n787), .A2(new_n788), .ZN(new_n816));
  OAI21_X1  g615(.A(G155gat), .B1(new_n816), .B2(new_n520), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n764), .A2(new_n266), .A3(new_n585), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1346gat));
  OAI21_X1  g618(.A(G162gat), .B1(new_n816), .B2(new_n582), .ZN(new_n820));
  INV_X1    g619(.A(new_n764), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n582), .A2(G162gat), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n820), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT119), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n820), .B(new_n826), .C1(new_n821), .C2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1347gat));
  NOR2_X1   g627(.A1(new_n561), .A2(new_n338), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n741), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n249), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(new_n348), .ZN(G1348gat));
  NOR2_X1   g631(.A1(new_n830), .A2(new_n557), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(new_n349), .ZN(G1349gat));
  OAI21_X1  g633(.A(new_n351), .B1(new_n830), .B2(new_n520), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n741), .A2(new_n585), .A3(new_n829), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n345), .ZN(new_n837));
  XNOR2_X1  g636(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n837), .B(new_n838), .ZN(G1350gat));
  NOR2_X1   g638(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n576), .A2(new_n573), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n808), .A2(new_n841), .A3(new_n491), .A4(new_n829), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n842), .A2(new_n843), .A3(G190gat), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n842), .B2(G190gat), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n840), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(G190gat), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT121), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n842), .A2(new_n843), .A3(G190gat), .ZN(new_n849));
  XOR2_X1   g648(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n842), .A2(new_n341), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n846), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT123), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n846), .A2(new_n851), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1351gat));
  NAND4_X1  g656(.A1(new_n808), .A2(new_n576), .A3(new_n447), .A4(new_n829), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(G197gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n248), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n447), .A2(new_n829), .ZN(new_n862));
  XOR2_X1   g661(.A(new_n862), .B(KEYINPUT124), .Z(new_n863));
  NAND2_X1  g662(.A1(new_n810), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n249), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n861), .B1(new_n865), .B2(new_n860), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT125), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n868), .B(new_n861), .C1(new_n865), .C2(new_n860), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1352gat));
  OAI21_X1  g669(.A(G204gat), .B1(new_n864), .B2(new_n557), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n557), .A2(G204gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n859), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT62), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n871), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n871), .A2(KEYINPUT126), .A3(new_n874), .A4(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1353gat));
  NAND3_X1  g680(.A1(new_n859), .A2(new_n258), .A3(new_n585), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n810), .A2(new_n585), .A3(new_n863), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n883), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT63), .B1(new_n883), .B2(G211gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1354gat));
  NOR3_X1   g685(.A1(new_n864), .A2(new_n257), .A3(new_n582), .ZN(new_n887));
  AOI21_X1  g686(.A(G218gat), .B1(new_n859), .B2(new_n491), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(G1355gat));
endmodule


