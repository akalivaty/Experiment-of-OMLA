//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT65), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n202), .C2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n214), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n220), .A2(new_n215), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n208), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n231), .B(new_n234), .C1(new_n223), .C2(new_n224), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n226), .A2(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n256), .A3(G274), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  AND2_X1   g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(new_n255), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT67), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(new_n254), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G226), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n254), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n264), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n277), .A2(G223), .B1(new_n280), .B2(G77), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1698), .B1(new_n275), .B2(new_n276), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G222), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n266), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n271), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n269), .A2(new_n270), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G200), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(G190), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n229), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G150), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT8), .B(G58), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n274), .A2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(G58), .A2(G68), .ZN(new_n300));
  INV_X1    g0100(.A(G50), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n207), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n293), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n206), .A2(G20), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G50), .ZN(new_n306));
  XOR2_X1   g0106(.A(new_n306), .B(KEYINPUT69), .Z(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n229), .A3(new_n292), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n303), .B1(G50), .B2(new_n304), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT9), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n290), .A2(new_n291), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(G169), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n289), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n288), .A2(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n314), .A2(new_n309), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n275), .A2(new_n276), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(G232), .A3(G1698), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(G226), .A3(new_n272), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n266), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n258), .A2(new_n263), .B1(G238), .B2(new_n267), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n324), .B2(new_n325), .ZN(new_n328));
  OAI21_X1  g0128(.A(G200), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n304), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n210), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT12), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n294), .A2(G50), .B1(G20), .B2(new_n210), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n298), .B2(new_n212), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n335));
  INV_X1    g0135(.A(new_n308), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G68), .A3(new_n305), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT11), .B1(new_n334), .B2(new_n293), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n267), .A2(G238), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n264), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n282), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n256), .B1(new_n343), .B2(new_n320), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT13), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(G190), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n329), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT14), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n345), .A2(G179), .A3(new_n346), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT14), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(G169), .C1(new_n327), .C2(new_n328), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n340), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n349), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n293), .ZN(new_n358));
  INV_X1    g0158(.A(new_n296), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n297), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n358), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n336), .A2(G77), .A3(new_n305), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT70), .B1(new_n330), .B2(new_n212), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n330), .A2(KEYINPUT70), .A3(new_n212), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n277), .A2(G238), .B1(new_n280), .B2(G107), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n319), .A2(G232), .A3(new_n272), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n266), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n258), .A2(new_n263), .B1(G244), .B2(new_n267), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n369), .B1(new_n375), .B2(new_n313), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n315), .A3(new_n374), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(G200), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n379), .B(new_n369), .C1(new_n380), .C2(new_n375), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n312), .A2(new_n318), .A3(new_n357), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G58), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n210), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n300), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n294), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT71), .B(G33), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n279), .B1(new_n392), .B2(KEYINPUT3), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n391), .B1(new_n393), .B2(new_n207), .ZN(new_n394));
  AND2_X1   g0194(.A1(KEYINPUT71), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT71), .A2(G33), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT3), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n397), .A2(new_n391), .A3(new_n207), .A4(new_n275), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G68), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n390), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n392), .B2(KEYINPUT3), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n276), .A2(new_n207), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n391), .B1(new_n403), .B2(new_n279), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n210), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n389), .B1(new_n405), .B2(new_n388), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n400), .A2(new_n406), .A3(new_n293), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n296), .B1(new_n206), .B2(G20), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n336), .B1(new_n330), .B2(new_n296), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n265), .A2(G1698), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G223), .B2(G1698), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n275), .B2(new_n397), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n274), .A2(new_n217), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n266), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n256), .A2(G232), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n258), .B2(new_n263), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n417), .A3(new_n380), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(G200), .B1(new_n414), .B2(new_n417), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n407), .B(new_n409), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT17), .ZN(new_n422));
  INV_X1    g0222(.A(new_n409), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n397), .A2(new_n207), .A3(new_n275), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT7), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(G68), .A3(new_n398), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n358), .B1(new_n426), .B2(new_n390), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n423), .B1(new_n427), .B2(new_n406), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n414), .A2(new_n417), .A3(G179), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n313), .B1(new_n414), .B2(new_n417), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT18), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT72), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n407), .A2(new_n409), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n414), .A2(new_n417), .A3(G179), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n414), .A2(new_n417), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(new_n313), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n432), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n433), .B1(new_n432), .B2(new_n439), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n422), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n383), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT77), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n294), .A2(G77), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G97), .A2(G107), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT6), .B1(new_n204), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT6), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n448), .A2(new_n202), .A3(G107), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n445), .B1(new_n450), .B2(new_n207), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n203), .B1(new_n402), .B2(new_n404), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n293), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n304), .A2(G97), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT73), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n274), .B2(G1), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n206), .A2(KEYINPUT73), .A3(G33), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n308), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n454), .B1(new_n459), .B2(G97), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g0261(.A(KEYINPUT74), .B(KEYINPUT4), .Z(new_n462));
  NAND2_X1  g0262(.A1(new_n397), .A2(new_n275), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n213), .A2(G1698), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT4), .A2(G244), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n319), .A2(new_n272), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(G250), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n266), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n206), .A2(G45), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G257), .A3(new_n256), .ZN(new_n476));
  OR2_X1    g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n261), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n471), .A2(new_n380), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(G200), .B1(new_n471), .B2(new_n482), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n461), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n471), .A2(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n313), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n453), .A2(new_n460), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n471), .A2(new_n315), .A3(new_n482), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(KEYINPUT71), .A2(G33), .ZN(new_n492));
  NAND2_X1  g0292(.A1(KEYINPUT71), .A2(G33), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n273), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n207), .B(G68), .C1(new_n494), .C2(new_n279), .ZN(new_n495));
  NOR3_X1   g0295(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n496));
  AOI21_X1  g0296(.A(G20), .B1(G33), .B2(G97), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT19), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT19), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n297), .A2(new_n499), .A3(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n358), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g0302(.A1(new_n308), .A2(new_n458), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n217), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n362), .A2(new_n304), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n266), .A2(new_n259), .A3(new_n473), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT75), .B1(new_n253), .B2(G1), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT75), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(new_n206), .A3(G45), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n256), .A2(new_n508), .A3(new_n510), .A4(G250), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT76), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n218), .B1(new_n260), .B2(new_n255), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n514), .A2(KEYINPUT76), .A3(new_n510), .A4(new_n508), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n507), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n211), .A2(new_n272), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n213), .A2(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n397), .B2(new_n275), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n395), .A2(new_n396), .ZN(new_n521));
  INV_X1    g0321(.A(G116), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n266), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G200), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n516), .A2(new_n524), .A3(G190), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n506), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(new_n313), .ZN(new_n529));
  INV_X1    g0329(.A(new_n505), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n459), .A2(new_n362), .ZN(new_n531));
  AOI21_X1  g0331(.A(G20), .B1(new_n397), .B2(new_n275), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(G68), .B1(new_n498), .B2(new_n500), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n530), .B(new_n531), .C1(new_n533), .C2(new_n358), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n516), .A2(new_n524), .A3(new_n315), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n529), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n444), .B1(new_n491), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n471), .A2(new_n380), .A3(new_n482), .ZN(new_n539));
  INV_X1    g0339(.A(new_n469), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n277), .B2(G250), .ZN(new_n541));
  INV_X1    g0341(.A(new_n464), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n397), .B2(new_n275), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n541), .B(new_n467), .C1(new_n543), .C2(new_n462), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n481), .B1(new_n544), .B2(new_n266), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n539), .B1(new_n545), .B2(G200), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n545), .A2(new_n315), .B1(new_n453), .B2(new_n460), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n461), .A2(new_n546), .B1(new_n547), .B2(new_n487), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n528), .A2(new_n536), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(KEYINPUT77), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n538), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n218), .A2(new_n272), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n219), .A2(G1698), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n397), .B2(new_n275), .ZN(new_n555));
  INV_X1    g0355(.A(G294), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n521), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n266), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n472), .A2(new_n474), .B1(new_n260), .B2(new_n255), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G264), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n480), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n313), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n558), .A2(new_n315), .A3(new_n480), .A4(new_n560), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n203), .A2(G20), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT23), .ZN(new_n567));
  XNOR2_X1  g0367(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n392), .A2(new_n207), .A3(G116), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT22), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n532), .B2(G87), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n207), .A3(G87), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n280), .B2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n217), .A2(KEYINPUT22), .A3(G20), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n319), .A2(KEYINPUT82), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n571), .B1(new_n573), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT24), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n207), .B(G87), .C1(new_n494), .C2(new_n279), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT22), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n576), .A2(new_n578), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n571), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n358), .B1(new_n581), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n503), .A2(new_n203), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n304), .A2(G107), .ZN(new_n590));
  XNOR2_X1  g0390(.A(KEYINPUT83), .B(KEYINPUT25), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n565), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n586), .B1(new_n585), .B2(new_n571), .ZN(new_n596));
  AOI211_X1 g0396(.A(KEYINPUT24), .B(new_n570), .C1(new_n583), .C2(new_n584), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n293), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(G200), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n561), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(G190), .B2(new_n561), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n593), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n219), .A2(new_n272), .ZN(new_n604));
  INV_X1    g0404(.A(G264), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G1698), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n607), .B1(new_n397), .B2(new_n275), .ZN(new_n608));
  XNOR2_X1  g0408(.A(KEYINPUT78), .B(G303), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n319), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n266), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n559), .A2(G270), .B1(new_n261), .B2(new_n479), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n611), .A2(new_n612), .A3(G179), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n330), .A2(new_n522), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n469), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT20), .ZN(new_n616));
  AOI22_X1  g0416(.A1(KEYINPUT80), .A2(new_n616), .B1(new_n522), .B2(G20), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n617), .A3(new_n293), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n616), .A2(KEYINPUT80), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n615), .A2(new_n617), .A3(new_n293), .A4(new_n619), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT79), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n459), .B2(G116), .ZN(new_n625));
  NOR4_X1   g0425(.A1(new_n308), .A2(new_n458), .A3(KEYINPUT79), .A4(new_n522), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n614), .B(new_n623), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n613), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT81), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT81), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n613), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n313), .B1(new_n611), .B2(new_n612), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n627), .A2(KEYINPUT21), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT21), .B1(new_n627), .B2(new_n633), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n611), .A2(new_n612), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n627), .B1(G200), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n611), .A2(new_n612), .A3(G190), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n632), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n603), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n443), .A2(new_n551), .A3(new_n642), .ZN(G372));
  INV_X1    g0443(.A(KEYINPUT84), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n537), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n528), .A2(new_n536), .A3(KEYINPUT84), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n548), .A3(new_n602), .A4(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n635), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n627), .A2(new_n633), .A3(KEYINPUT21), .ZN(new_n649));
  INV_X1    g0449(.A(new_n631), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n630), .B1(new_n613), .B2(new_n627), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n564), .B1(new_n598), .B2(new_n593), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n490), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n645), .A2(new_n656), .A3(new_n657), .A4(new_n646), .ZN(new_n658));
  INV_X1    g0458(.A(new_n536), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n528), .A2(new_n536), .A3(new_n547), .A4(new_n487), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n443), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT85), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n434), .A2(new_n665), .A3(new_n438), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n434), .B2(new_n438), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n435), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT85), .B1(new_n428), .B2(new_n431), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(KEYINPUT18), .A3(new_n666), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n378), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n355), .A2(new_n356), .B1(new_n673), .B2(new_n348), .ZN(new_n674));
  INV_X1    g0474(.A(new_n422), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n317), .B1(new_n312), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n664), .A2(new_n677), .ZN(G369));
  NAND3_X1  g0478(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n595), .A2(new_n652), .A3(new_n602), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n653), .A2(new_n685), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT87), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(KEYINPUT87), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n627), .A2(new_n684), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT86), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n641), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n652), .A2(new_n694), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n595), .A2(new_n602), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n684), .B1(new_n588), .B2(new_n594), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n653), .A2(new_n684), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n691), .A2(new_n703), .ZN(G399));
  NAND2_X1  g0504(.A1(new_n496), .A2(new_n522), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n232), .A2(new_n252), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(G1), .ZN(new_n708));
  INV_X1    g0508(.A(new_n228), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  AOI21_X1  g0511(.A(G179), .B1(new_n516), .B2(new_n524), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n486), .A2(new_n712), .A3(new_n561), .A4(new_n637), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n516), .A2(new_n524), .A3(new_n558), .A4(new_n560), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n611), .A2(new_n612), .A3(G179), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n486), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n713), .B1(new_n716), .B2(KEYINPUT30), .ZN(new_n717));
  INV_X1    g0517(.A(new_n714), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n545), .A4(new_n613), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n684), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n516), .A2(new_n524), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n558), .A2(new_n560), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n545), .A2(new_n724), .A3(new_n613), .A4(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n719), .A3(new_n713), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n684), .B1(new_n538), .B2(new_n550), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(new_n642), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT88), .B1(new_n733), .B2(new_n692), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n551), .A2(new_n642), .A3(new_n685), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n729), .B2(new_n684), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT88), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(new_n740), .A3(G330), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n663), .A2(new_n685), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n536), .A2(KEYINPUT89), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT89), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n529), .A2(new_n747), .A3(new_n534), .A4(new_n535), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n660), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(new_n750), .B2(new_n657), .ZN(new_n751));
  INV_X1    g0551(.A(new_n646), .ZN(new_n752));
  AOI21_X1  g0552(.A(KEYINPUT84), .B1(new_n528), .B2(new_n536), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n752), .A2(new_n753), .A3(new_n490), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n751), .B1(new_n754), .B2(new_n657), .ZN(new_n755));
  OAI211_X1 g0555(.A(KEYINPUT29), .B(new_n685), .C1(new_n755), .C2(new_n655), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n742), .B1(new_n745), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n711), .B1(new_n757), .B2(G1), .ZN(G364));
  INV_X1    g0558(.A(new_n707), .ZN(new_n759));
  INV_X1    g0559(.A(G13), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n206), .B1(new_n761), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n319), .A2(new_n232), .ZN(new_n765));
  INV_X1    g0565(.A(G355), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n765), .A2(new_n766), .B1(G116), .B2(new_n232), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n247), .A2(new_n253), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n393), .A2(new_n232), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n253), .B2(new_n228), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n229), .B1(G20), .B2(new_n313), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n764), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n207), .A2(new_n315), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n207), .A2(G179), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(new_n380), .A3(G200), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n782), .A2(new_n210), .B1(new_n784), .B2(new_n203), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n779), .A2(G190), .A3(new_n599), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n319), .B1(new_n786), .B2(new_n384), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n780), .A2(new_n380), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n301), .B1(new_n790), .B2(new_n217), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n779), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n787), .B(new_n791), .C1(G77), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n783), .A2(new_n792), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT32), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n380), .A2(G179), .A3(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n207), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n785), .B(new_n800), .C1(G97), .C2(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT90), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT90), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  INV_X1    g0607(.A(G329), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n784), .A2(new_n807), .B1(new_n796), .B2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT91), .Z(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n280), .B1(new_n793), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n786), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G322), .B2(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G294), .A2(new_n803), .B1(new_n788), .B2(G326), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  INV_X1    g0616(.A(new_n790), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n781), .A2(new_n816), .B1(new_n817), .B2(G303), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n810), .A2(new_n814), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n805), .A2(new_n806), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n778), .B1(new_n820), .B2(new_n775), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n695), .A2(new_n696), .ZN(new_n822));
  INV_X1    g0622(.A(new_n774), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(G330), .ZN(new_n825));
  INV_X1    g0625(.A(new_n697), .ZN(new_n826));
  INV_X1    g0626(.A(new_n764), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n824), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT92), .Z(G396));
  INV_X1    g0630(.A(new_n742), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n381), .B1(new_n369), .B2(new_n685), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n378), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n378), .A2(new_n684), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n743), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n836), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n838), .B(new_n685), .C1(new_n655), .C2(new_n662), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n827), .B1(new_n831), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n831), .A2(new_n840), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(KEYINPUT96), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(KEYINPUT96), .B2(new_n842), .ZN(new_n844));
  INV_X1    g0644(.A(new_n775), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n802), .A2(new_n202), .B1(new_n786), .B2(new_n556), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT93), .Z(new_n847));
  OAI221_X1 g0647(.A(new_n280), .B1(new_n796), .B2(new_n811), .C1(new_n522), .C2(new_n793), .ZN(new_n848));
  INV_X1    g0648(.A(G303), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n789), .A2(new_n849), .B1(new_n784), .B2(new_n217), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n782), .A2(new_n807), .B1(new_n790), .B2(new_n203), .ZN(new_n851));
  OR4_X1    g0651(.A1(new_n847), .A2(new_n848), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n813), .A2(G143), .B1(new_n794), .B2(G159), .ZN(new_n853));
  INV_X1    g0653(.A(G150), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n782), .B2(new_n854), .C1(new_n855), .C2(new_n789), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT94), .Z(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n802), .A2(new_n384), .B1(new_n784), .B2(new_n210), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n463), .B1(new_n860), .B2(new_n796), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n859), .B(new_n861), .C1(G50), .C2(new_n817), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n852), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT95), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n845), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n866), .B2(new_n865), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n775), .A2(new_n772), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n827), .B1(new_n212), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n868), .B(new_n870), .C1(new_n773), .C2(new_n838), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n844), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  NOR2_X1   g0673(.A1(new_n761), .A2(new_n206), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n356), .A2(new_n684), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT97), .B1(new_n357), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n354), .A2(new_n352), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n345), .A2(new_n346), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n353), .B1(new_n878), .B2(G169), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n356), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AND4_X1   g0680(.A1(KEYINPUT97), .A2(new_n880), .A3(new_n348), .A4(new_n875), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n355), .A2(new_n349), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n876), .A2(new_n881), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(KEYINPUT100), .A2(KEYINPUT31), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n721), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n729), .A2(new_n684), .A3(new_n884), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n735), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n883), .A2(new_n838), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  INV_X1    g0694(.A(new_n682), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n434), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n672), .B2(new_n422), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT98), .B1(new_n428), .B2(new_n431), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT98), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n434), .A2(new_n899), .A3(new_n438), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n896), .A2(new_n902), .A3(new_n421), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n682), .B1(new_n407), .B2(new_n409), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n418), .B1(new_n437), .B2(G200), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n428), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n667), .B2(new_n668), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n904), .B1(KEYINPUT37), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n894), .B1(new_n897), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT99), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n400), .A2(new_n293), .ZN(new_n912));
  INV_X1    g0712(.A(new_n388), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT16), .B1(new_n426), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n409), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n915), .A2(new_n895), .B1(new_n428), .B2(new_n906), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n438), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n902), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n911), .B1(new_n904), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n907), .A2(new_n902), .A3(new_n898), .A4(new_n900), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n426), .A2(new_n913), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n389), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n423), .B1(new_n922), .B2(new_n427), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n421), .B1(new_n923), .B2(new_n682), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n431), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT37), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n920), .A2(new_n926), .A3(KEYINPUT99), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n923), .A2(new_n682), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n442), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(KEYINPUT38), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n910), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n893), .B(new_n932), .C1(KEYINPUT101), .C2(new_n890), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT40), .ZN(new_n934));
  INV_X1    g0734(.A(new_n893), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n904), .A2(new_n918), .A3(new_n911), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT99), .B1(new_n920), .B2(new_n926), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n930), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n894), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n931), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n443), .A2(new_n889), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n692), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n932), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n939), .A2(KEYINPUT39), .A3(new_n931), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n355), .A2(new_n356), .A3(new_n685), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n839), .A2(new_n835), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n940), .A2(new_n952), .A3(new_n883), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n672), .B2(new_n895), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n745), .A2(new_n756), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n383), .A2(new_n442), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n677), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n955), .B(new_n958), .Z(new_n959));
  AOI21_X1  g0759(.A(new_n874), .B1(new_n945), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n959), .B2(new_n945), .ZN(new_n961));
  INV_X1    g0761(.A(new_n450), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(KEYINPUT35), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(KEYINPUT35), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n963), .A2(G116), .A3(new_n230), .A4(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT36), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n709), .A2(new_n212), .A3(new_n385), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n210), .A2(G50), .ZN(new_n968));
  OAI211_X1 g0768(.A(G1), .B(new_n760), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n961), .A2(new_n966), .A3(new_n969), .ZN(G367));
  INV_X1    g0770(.A(KEYINPUT109), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n548), .B1(new_n461), .B2(new_n685), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n656), .A2(new_n684), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT105), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT44), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n691), .A2(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n974), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n975), .A2(new_n976), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n689), .A2(new_n690), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n977), .B(new_n980), .C1(KEYINPUT105), .C2(KEYINPUT44), .ZN(new_n981));
  INV_X1    g0781(.A(new_n690), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n974), .B1(new_n982), .B2(new_n688), .ZN(new_n983));
  XNOR2_X1  g0783(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n986), .A2(KEYINPUT106), .A3(new_n697), .A4(new_n702), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n697), .A2(KEYINPUT108), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n686), .A2(KEYINPUT107), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT108), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n989), .B1(new_n826), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n686), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n652), .A2(new_n685), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n700), .A2(new_n993), .A3(new_n701), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT107), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n988), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n988), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n697), .A2(KEYINPUT108), .B1(KEYINPUT107), .B2(new_n686), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n999), .A2(new_n1000), .A3(new_n996), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n956), .A2(new_n741), .A3(new_n734), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n981), .A2(new_n703), .A3(new_n985), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n987), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n703), .B1(new_n981), .B2(new_n985), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(KEYINPUT106), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n757), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n707), .B(KEYINPUT41), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n763), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n992), .A2(new_n974), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT42), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n490), .B1(new_n972), .B2(new_n595), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n685), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n645), .A2(new_n646), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n506), .A2(new_n685), .ZN(new_n1018));
  MUX2_X1   g0818(.A(new_n1017), .B(new_n536), .S(new_n1018), .Z(new_n1019));
  INV_X1    g0819(.A(KEYINPUT102), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT43), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n703), .A2(new_n978), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1016), .A2(new_n1024), .B1(KEYINPUT103), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n1016), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1025), .A2(KEYINPUT103), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n971), .B1(new_n1012), .B2(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1007), .A2(KEYINPUT106), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1034), .A2(new_n987), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1010), .B1(new_n1035), .B2(new_n757), .ZN(new_n1036));
  OAI211_X1 g0836(.A(KEYINPUT109), .B(new_n1031), .C1(new_n1036), .C2(new_n763), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n776), .B1(new_n232), .B2(new_n361), .C1(new_n243), .C2(new_n769), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n786), .A2(new_n854), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n802), .A2(new_n210), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G143), .C2(new_n788), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1042), .A2(KEYINPUT111), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1042), .A2(KEYINPUT111), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n319), .B1(new_n796), .B2(new_n855), .C1(new_n301), .C2(new_n793), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n784), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(G77), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n384), .B2(new_n790), .C1(new_n782), .C2(new_n797), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT112), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT110), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n796), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G283), .A2(new_n794), .B1(new_n1053), .B2(G317), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n609), .B2(new_n786), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n463), .B(new_n1055), .C1(G97), .C2(new_n1046), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n789), .A2(new_n811), .B1(new_n203), .B2(new_n802), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G294), .B2(new_n781), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n790), .A2(new_n522), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1056), .B(new_n1058), .C1(KEYINPUT46), .C2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1050), .B1(new_n1052), .B2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT47), .Z(new_n1062));
  OAI211_X1 g0862(.A(new_n764), .B(new_n1039), .C1(new_n1062), .C2(new_n845), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1019), .A2(new_n774), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1038), .A2(new_n1066), .ZN(G387));
  OR2_X1    g0867(.A1(new_n998), .A2(new_n1001), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n700), .A2(new_n701), .A3(new_n774), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n706), .A2(new_n765), .B1(G107), .B2(new_n232), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n240), .A2(new_n253), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n296), .A2(G50), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT50), .ZN(new_n1073));
  AOI211_X1 g0873(.A(G45), .B(new_n705), .C1(G68), .C2(G77), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n769), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1070), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n764), .B1(new_n1076), .B2(new_n777), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n790), .A2(new_n212), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT113), .B(G150), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n463), .B1(new_n796), .B2(new_n1079), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(G97), .C2(new_n1046), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT114), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n781), .A2(new_n359), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n813), .A2(G50), .B1(new_n794), .B2(G68), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n362), .A2(new_n803), .B1(new_n788), .B2(G159), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n463), .B1(G326), .B2(new_n1053), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n802), .A2(new_n807), .B1(new_n790), .B2(new_n556), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n609), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n813), .A2(G317), .B1(new_n794), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n788), .A2(G322), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n811), .C2(new_n782), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1088), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1093), .B2(new_n1092), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT49), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1087), .B1(new_n522), .B2(new_n784), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1086), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT115), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n845), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1077), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1068), .A2(new_n763), .B1(new_n1069), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1068), .A2(new_n757), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n759), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1068), .A2(new_n757), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT116), .Z(G393));
  INV_X1    g0909(.A(new_n1007), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1005), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n707), .B1(new_n1111), .B2(new_n1105), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1112), .A2(new_n1035), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n776), .B1(new_n202), .B2(new_n232), .C1(new_n250), .C2(new_n769), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n764), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n802), .A2(new_n212), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n782), .A2(new_n301), .B1(new_n784), .B2(new_n217), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(G68), .C2(new_n817), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n789), .A2(new_n854), .B1(new_n797), .B2(new_n786), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT51), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n359), .A2(new_n794), .B1(new_n1053), .B2(G143), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n463), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G317), .A2(new_n788), .B1(new_n813), .B2(G311), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT52), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n803), .A2(G116), .B1(new_n817), .B2(G283), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n781), .A2(new_n1089), .B1(new_n1046), .B2(G107), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n794), .A2(G294), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n319), .B1(new_n1053), .B2(G322), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1122), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1115), .B1(new_n1130), .B2(new_n775), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n974), .B2(new_n823), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1111), .B2(new_n762), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1113), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(G390));
  NAND2_X1  g0935(.A1(new_n949), .A2(new_n772), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n869), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n764), .B1(new_n359), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT119), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1116), .B1(G283), .B2(new_n788), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n203), .B2(new_n782), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n817), .A2(G87), .B1(new_n1046), .B2(G68), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n319), .B1(new_n813), .B2(G116), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G97), .A2(new_n794), .B1(new_n1053), .B2(G294), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G159), .A2(new_n803), .B1(new_n788), .B2(G128), .ZN(new_n1146));
  INV_X1    g0946(.A(G125), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n786), .A2(new_n860), .B1(new_n796), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n319), .B1(new_n793), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n781), .A2(G137), .B1(new_n1046), .B2(G50), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1146), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n790), .A2(new_n1079), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT53), .Z(new_n1155));
  OAI22_X1  g0955(.A1(new_n1141), .A2(new_n1145), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT120), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n775), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1136), .B(new_n1139), .C1(new_n1158), .C2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT117), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n692), .B1(new_n735), .B2(new_n888), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n838), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n883), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1162), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n692), .B(new_n836), .C1(new_n735), .C2(new_n888), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(KEYINPUT117), .A3(new_n883), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n950), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n952), .B2(new_n883), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n947), .B2(new_n948), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1170), .B1(new_n910), .B2(new_n931), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n685), .B(new_n833), .C1(new_n755), .C2(new_n655), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n835), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n883), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1169), .B1(new_n1172), .B2(new_n1177), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n839), .A2(new_n835), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n950), .B1(new_n1179), .B2(new_n1165), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n928), .A2(KEYINPUT38), .A3(new_n930), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT38), .B1(new_n928), .B2(new_n930), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1181), .A2(new_n1182), .A3(new_n946), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT39), .B1(new_n910), .B2(new_n931), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n740), .B1(new_n739), .B2(G330), .ZN(new_n1187));
  AOI211_X1 g0987(.A(KEYINPUT88), .B(new_n692), .C1(new_n735), .C2(new_n738), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n838), .B(new_n883), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1178), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1161), .B1(new_n1191), .B2(new_n762), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT121), .Z(new_n1193));
  AND2_X1   g0993(.A1(new_n1178), .A2(new_n1190), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n443), .A2(new_n1163), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1195), .B(new_n677), .C1(new_n956), .C2(new_n957), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n883), .B1(new_n742), .B2(new_n838), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n952), .B1(new_n1197), .B2(new_n1169), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1175), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1189), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1196), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT118), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1194), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1196), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT117), .B1(new_n1167), .B2(new_n883), .ZN(new_n1205));
  AND4_X1   g1005(.A1(KEYINPUT117), .A2(new_n1163), .A3(new_n883), .A4(new_n838), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n838), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1165), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1179), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1200), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1204), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(KEYINPUT118), .B1(new_n1212), .B2(new_n1191), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1203), .A2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1214), .B(new_n759), .C1(new_n1194), .C2(new_n1201), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1193), .A2(new_n1215), .ZN(G378));
  NAND2_X1  g1016(.A1(new_n312), .A2(new_n318), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n309), .A2(new_n895), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1217), .B(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1219), .B(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n942), .A2(G330), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1221), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n933), .A2(KEYINPUT40), .B1(new_n940), .B2(new_n935), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n1224), .B2(new_n692), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n955), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1222), .A2(new_n1225), .A3(new_n955), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1223), .A2(new_n772), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n764), .B1(G50), .B2(new_n1137), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1147), .A2(new_n789), .B1(new_n782), .B2(new_n860), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n813), .A2(G128), .B1(new_n794), .B2(G137), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n790), .B2(new_n1149), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(G150), .C2(new_n803), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1239));
  XOR2_X1   g1039(.A(KEYINPUT122), .B(G124), .Z(new_n1240));
  OAI211_X1 g1040(.A(new_n274), .B(new_n252), .C1(new_n1240), .C2(new_n796), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(G159), .B2(new_n1046), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1238), .A2(new_n1239), .A3(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n813), .A2(G107), .B1(new_n1053), .B2(G283), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n361), .B2(new_n793), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n393), .A2(new_n252), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n1041), .A4(new_n1078), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n788), .A2(G116), .B1(new_n1046), .B2(G58), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n202), .C2(new_n782), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT58), .ZN(new_n1250));
  OR2_X1    g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1246), .B(new_n301), .C1(G33), .C2(G41), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1243), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1232), .B1(new_n1254), .B2(new_n775), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1230), .A2(new_n763), .B1(new_n1231), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1202), .B1(new_n1194), .B2(new_n1201), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1212), .A2(new_n1191), .A3(KEYINPUT118), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1204), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT123), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1214), .A2(KEYINPUT123), .A3(new_n1204), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT57), .B1(new_n1263), .B2(new_n1230), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT57), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT123), .B1(new_n1214), .B2(new_n1204), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1260), .B(new_n1196), .C1(new_n1203), .C2(new_n1213), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n759), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1256), .B1(new_n1264), .B2(new_n1270), .ZN(G375));
  OAI22_X1  g1071(.A1(new_n782), .A2(new_n1149), .B1(new_n855), .B2(new_n786), .ZN(new_n1272));
  INV_X1    g1072(.A(G128), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n793), .A2(new_n854), .B1(new_n796), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G50), .B2(new_n803), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1046), .A2(G58), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT125), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n463), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(new_n1276), .B2(new_n463), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1275), .B1(new_n797), .B2(new_n790), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT126), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n1272), .B(new_n1282), .C1(G132), .C2(new_n788), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n788), .A2(G294), .B1(new_n794), .B2(G107), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n522), .B2(new_n782), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT124), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n280), .B1(new_n796), .B2(new_n849), .C1(new_n786), .C2(new_n807), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1047), .B1(new_n202), .B2(new_n790), .C1(new_n361), .C2(new_n802), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n775), .B1(new_n1283), .B2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1290), .B(new_n764), .C1(G68), .C2(new_n1137), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1165), .B2(new_n772), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n763), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1212), .A2(new_n1011), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1293), .A2(new_n1204), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(G381));
  INV_X1    g1097(.A(new_n1256), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n707), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1230), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1265), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1298), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  OR2_X1    g1102(.A1(G393), .A2(G396), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1134), .A2(new_n872), .ZN(new_n1304));
  NOR4_X1   g1104(.A1(new_n1303), .A2(G378), .A3(new_n1304), .A4(G381), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1302), .A2(new_n1038), .A3(new_n1305), .A4(new_n1066), .ZN(G407));
  INV_X1    g1106(.A(G378), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n683), .A2(G213), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1302), .A2(new_n1307), .A3(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(G407), .A2(G213), .A3(new_n1310), .ZN(G409));
  OAI211_X1 g1111(.A(G378), .B(new_n1256), .C1(new_n1264), .C2(new_n1270), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1256), .B1(new_n1300), .B2(new_n1010), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1307), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT60), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1201), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1296), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n759), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1317), .A2(new_n1296), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1294), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1321), .A2(new_n872), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n872), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1315), .A2(new_n1308), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(KEYINPUT62), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT61), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1309), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1325), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1309), .A2(G2897), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1324), .B(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1263), .A2(new_n1011), .A3(new_n1230), .ZN(new_n1334));
  AOI21_X1  g1134(.A(G378), .B1(new_n1334), .B2(new_n1256), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1335), .B1(new_n1302), .B2(G378), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1333), .B1(new_n1336), .B2(new_n1309), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1327), .A2(new_n1328), .A3(new_n1331), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G387), .A2(new_n1134), .ZN(new_n1339));
  XOR2_X1   g1139(.A(G393), .B(G396), .Z(new_n1340));
  NAND3_X1  g1140(.A1(new_n1038), .A2(new_n1066), .A3(G390), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1339), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(G393), .B(G396), .ZN(new_n1343));
  AOI21_X1  g1143(.A(G390), .B1(new_n1038), .B2(new_n1066), .ZN(new_n1344));
  AOI211_X1 g1144(.A(new_n1065), .B(new_n1134), .C1(new_n1033), .C2(new_n1037), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1343), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1342), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1338), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1332), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1324), .B(new_n1350), .ZN(new_n1351));
  OAI211_X1 g1151(.A(new_n1347), .B(new_n1328), .C1(new_n1329), .C2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT63), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1326), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT127), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1356), .B1(new_n1326), .B2(new_n1354), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1329), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1325), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1353), .A2(new_n1355), .A3(new_n1357), .A4(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1349), .A2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(G375), .A2(new_n1307), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1312), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(new_n1325), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1361), .A2(new_n1312), .A3(new_n1324), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  XNOR2_X1  g1165(.A(new_n1365), .B(new_n1348), .ZN(G402));
endmodule


