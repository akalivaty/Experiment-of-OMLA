//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G58), .A3(G68), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OR3_X1    g0007(.A1(new_n207), .A2(KEYINPUT65), .A3(G13), .ZN(new_n208));
  OAI21_X1  g0008(.A(KEYINPUT65), .B1(new_n207), .B2(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n206), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n214), .A2(KEYINPUT0), .ZN(new_n215));
  NOR2_X1   g0015(.A1(G58), .A2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT66), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(new_n217), .B2(new_n216), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT67), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n214), .A2(KEYINPUT0), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n215), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT68), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  INV_X1    g0028(.A(G68), .ZN(new_n229));
  INV_X1    g0029(.A(G238), .ZN(new_n230));
  INV_X1    g0030(.A(G87), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n206), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n233));
  INV_X1    g0033(.A(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G107), .ZN(new_n235));
  OAI221_X1 g0035(.A(new_n233), .B1(new_n203), .B2(new_n234), .C1(new_n235), .C2(new_n213), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n207), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n227), .A2(new_n238), .ZN(G361));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  INV_X1    g0045(.A(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(KEYINPUT2), .B(G226), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n244), .B(new_n249), .Z(G358));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT71), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(G68), .B(G77), .Z(new_n255));
  XOR2_X1   g0055(.A(G50), .B(G58), .Z(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n254), .B(new_n257), .Z(G351));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n260), .A2(new_n261), .A3(G274), .A4(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT72), .B(G226), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT73), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT73), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G1698), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(G222), .B2(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n260), .B1(new_n279), .B2(new_n203), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n269), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G179), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n221), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n261), .A2(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G50), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n297), .A2(new_n299), .B1(G50), .B2(new_n292), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT74), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n274), .B2(G20), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n222), .A2(KEYINPUT74), .A3(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G20), .A2(G33), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n302), .A2(new_n306), .B1(G150), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n202), .B2(new_n222), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n300), .B1(new_n309), .B2(new_n295), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n289), .A2(new_n291), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT75), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n312), .B(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n310), .A2(KEYINPUT9), .B1(new_n286), .B2(G190), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n310), .A2(KEYINPUT9), .B1(new_n317), .B2(new_n286), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT10), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n318), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT10), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n315), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n260), .B1(new_n279), .B2(new_n235), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G232), .A2(G1698), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n230), .B2(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n279), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n265), .ZN(new_n328));
  INV_X1    g0128(.A(new_n267), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(G244), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT76), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT76), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n327), .A2(new_n333), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G190), .ZN(new_n336));
  INV_X1    g0136(.A(new_n295), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT15), .B(G87), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n306), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n340), .A2(KEYINPUT77), .ZN(new_n341));
  INV_X1    g0141(.A(new_n307), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n301), .A2(new_n342), .B1(new_n222), .B2(new_n203), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n340), .B2(KEYINPUT77), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n337), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n296), .A2(G77), .A3(new_n298), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(G77), .B2(new_n292), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT78), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n332), .A2(new_n334), .A3(G200), .ZN(new_n350));
  OR3_X1    g0150(.A1(new_n345), .A2(KEYINPUT78), .A3(new_n347), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n336), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n335), .A2(new_n290), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n332), .A2(new_n334), .A3(new_n288), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n314), .A2(new_n323), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT18), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(KEYINPUT83), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n302), .A2(new_n298), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n297), .A2(new_n359), .B1(new_n292), .B2(new_n302), .ZN(new_n360));
  INV_X1    g0160(.A(G58), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(new_n229), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n362), .B2(new_n216), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n307), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n275), .A2(new_n222), .A3(new_n277), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT73), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n276), .B1(new_n275), .B2(new_n277), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n222), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n369), .B1(new_n372), .B2(new_n368), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n366), .B1(new_n373), .B2(new_n229), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n270), .A2(new_n271), .A3(G20), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT7), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT81), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n367), .A2(new_n379), .A3(new_n368), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n367), .B2(new_n368), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G68), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n365), .A2(new_n375), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n337), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n360), .B1(new_n376), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT82), .ZN(new_n387));
  INV_X1    g0187(.A(G1698), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n281), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G226), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G1698), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n389), .B(new_n391), .C1(new_n270), .C2(new_n271), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n260), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n260), .A2(G232), .A3(new_n266), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n265), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n288), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n260), .B1(new_n392), .B2(new_n393), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n265), .A2(new_n397), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n400), .A2(new_n401), .A3(new_n290), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n387), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(G169), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n396), .A2(new_n398), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT82), .B(new_n404), .C1(new_n405), .C2(new_n290), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n358), .B1(new_n386), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT81), .B1(new_n377), .B2(KEYINPUT7), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n367), .A2(new_n379), .A3(new_n368), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n369), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n384), .B1(new_n411), .B2(new_n229), .ZN(new_n412));
  AOI21_X1  g0212(.A(G20), .B1(new_n272), .B2(new_n278), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n378), .B1(new_n413), .B2(KEYINPUT7), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n365), .B1(new_n414), .B2(G68), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n412), .B(new_n295), .C1(new_n415), .C2(KEYINPUT16), .ZN(new_n416));
  INV_X1    g0216(.A(new_n360), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n405), .A2(new_n317), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n405), .B2(G190), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n416), .A2(new_n417), .ZN(new_n423));
  INV_X1    g0223(.A(new_n407), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n416), .A2(KEYINPUT17), .A3(new_n417), .A4(new_n419), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n408), .A2(new_n422), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n356), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT84), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT80), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G226), .A2(G1698), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n246), .B2(G1698), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n272), .A2(new_n433), .A3(new_n278), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT79), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT79), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n439), .A3(new_n395), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n265), .B1(new_n230), .B2(new_n267), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n431), .B1(new_n443), .B2(KEYINPUT13), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT13), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n440), .B2(new_n442), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n440), .A2(KEYINPUT80), .A3(new_n445), .A4(new_n442), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n444), .A2(new_n447), .A3(G190), .A4(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n260), .B1(new_n436), .B2(KEYINPUT79), .ZN(new_n450));
  AOI211_X1 g0250(.A(KEYINPUT13), .B(new_n441), .C1(new_n450), .C2(new_n439), .ZN(new_n451));
  OAI21_X1  g0251(.A(G200), .B1(new_n451), .B2(new_n446), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n293), .A2(new_n229), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT12), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n296), .A2(G68), .A3(new_n298), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT11), .ZN(new_n456));
  INV_X1    g0256(.A(G50), .ZN(new_n457));
  OAI22_X1  g0257(.A1(new_n342), .A2(new_n457), .B1(new_n222), .B2(G68), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n203), .B1(new_n304), .B2(new_n305), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n295), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n454), .B(new_n455), .C1(new_n456), .C2(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n460), .A2(new_n456), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n449), .A2(new_n452), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n463), .ZN(new_n465));
  OAI21_X1  g0265(.A(G169), .B1(new_n451), .B2(new_n446), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT14), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT14), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(G169), .C1(new_n451), .C2(new_n446), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n444), .A2(new_n447), .A3(G179), .A4(new_n448), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n464), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n429), .A2(new_n430), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n430), .B1(new_n429), .B2(new_n472), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n477), .A2(new_n234), .A3(G1698), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n272), .A2(new_n278), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT85), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT85), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n272), .A2(new_n278), .A3(new_n481), .A4(new_n478), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n272), .A2(new_n278), .A3(G250), .A4(G1698), .ZN(new_n483));
  OAI211_X1 g0283(.A(G244), .B(new_n388), .C1(new_n270), .C2(new_n271), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(new_n477), .B1(G33), .B2(G283), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n480), .A2(new_n482), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n395), .ZN(new_n487));
  INV_X1    g0287(.A(G274), .ZN(new_n488));
  INV_X1    g0288(.A(new_n221), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n259), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n263), .A2(G1), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n262), .A2(KEYINPUT86), .A3(KEYINPUT5), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT86), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(G41), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n491), .A3(new_n492), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n260), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n496), .B1(new_n498), .B2(new_n212), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n487), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n288), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n292), .A2(G97), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n261), .A2(G33), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n292), .A2(new_n505), .A3(new_n221), .A4(new_n294), .ZN(new_n506));
  INV_X1    g0306(.A(G97), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n510), .A2(new_n507), .A3(G107), .ZN(new_n511));
  XNOR2_X1  g0311(.A(G97), .B(G107), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n513), .A2(new_n222), .B1(new_n203), .B2(new_n342), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n414), .B2(G107), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n509), .B1(new_n515), .B2(new_n337), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n499), .B1(new_n486), .B2(new_n395), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n290), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n502), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n514), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n373), .B2(new_n235), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n508), .B1(new_n521), .B2(new_n295), .ZN(new_n522));
  AOI21_X1  g0322(.A(G200), .B1(new_n487), .B2(new_n500), .ZN(new_n523));
  AOI211_X1 g0323(.A(G190), .B(new_n499), .C1(new_n486), .C2(new_n395), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n206), .B1(new_n261), .B2(G45), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n490), .A2(new_n491), .B1(new_n260), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G238), .A2(G1698), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n234), .B2(G1698), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n275), .A2(new_n277), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n529), .A2(new_n530), .B1(G33), .B2(G116), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n527), .B(G190), .C1(new_n531), .C2(new_n260), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n230), .A2(new_n388), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n234), .A2(G1698), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(new_n270), .C2(new_n271), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n260), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n260), .A2(G274), .A3(new_n491), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n526), .A2(new_n260), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(G200), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n339), .A2(new_n292), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n506), .A2(new_n231), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n222), .B(G68), .C1(new_n270), .C2(new_n271), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n222), .B1(new_n435), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n231), .A2(new_n507), .A3(new_n235), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n507), .B1(new_n304), .B2(new_n305), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n545), .B(new_n549), .C1(new_n550), .C2(KEYINPUT19), .ZN(new_n551));
  AOI211_X1 g0351(.A(new_n543), .B(new_n544), .C1(new_n551), .C2(new_n295), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n295), .ZN(new_n553));
  INV_X1    g0353(.A(new_n543), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n506), .A2(new_n338), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n527), .B(G179), .C1(new_n531), .C2(new_n260), .ZN(new_n557));
  OAI21_X1  g0357(.A(G169), .B1(new_n537), .B2(new_n540), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n542), .A2(new_n552), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n519), .A2(new_n525), .A3(KEYINPUT87), .A4(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n519), .A2(new_n525), .A3(new_n560), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n222), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT22), .ZN(new_n566));
  OR3_X1    g0366(.A1(new_n231), .A2(KEYINPUT22), .A3(G20), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n279), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(G116), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n274), .A2(new_n569), .A3(G20), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT89), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n222), .B2(G107), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n572), .A2(KEYINPUT23), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(KEYINPUT23), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT24), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n568), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n337), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT25), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n292), .B2(G107), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n292), .A2(new_n581), .A3(G107), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n583), .A2(new_n584), .B1(new_n235), .B2(new_n506), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n497), .A2(G264), .A3(new_n260), .ZN(new_n586));
  INV_X1    g0386(.A(G294), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n274), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(G250), .A2(G1698), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n212), .B2(G1698), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n590), .B2(new_n530), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n496), .B(new_n586), .C1(new_n591), .C2(new_n260), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n206), .A2(new_n388), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n212), .A2(G1698), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n594), .B(new_n595), .C1(new_n270), .C2(new_n271), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n395), .B1(new_n597), .B2(new_n588), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(G190), .A3(new_n496), .A4(new_n586), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n580), .A2(new_n585), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n592), .A2(new_n288), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n598), .A2(new_n290), .A3(new_n496), .A4(new_n586), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n568), .A2(new_n578), .A3(new_n575), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n578), .B1(new_n568), .B2(new_n575), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n295), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n585), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(G303), .B1(new_n370), .B2(new_n371), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n212), .A2(new_n388), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n213), .A2(G1698), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n612), .B(new_n613), .C1(new_n270), .C2(new_n271), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT88), .B1(new_n615), .B2(new_n395), .ZN(new_n616));
  INV_X1    g0416(.A(G303), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n272), .B2(new_n278), .ZN(new_n618));
  INV_X1    g0418(.A(new_n614), .ZN(new_n619));
  OAI211_X1 g0419(.A(KEYINPUT88), .B(new_n395), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  MUX2_X1   g0422(.A(new_n292), .B(new_n506), .S(G116), .Z(new_n623));
  AOI22_X1  g0423(.A1(new_n294), .A2(new_n221), .B1(G20), .B2(new_n569), .ZN(new_n624));
  AOI21_X1  g0424(.A(G20), .B1(G33), .B2(G283), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(G33), .B2(new_n507), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT20), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n624), .A2(new_n626), .A3(KEYINPUT20), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G270), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n496), .B1(new_n498), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(G179), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n622), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n616), .B2(new_n621), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n629), .A2(G169), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT21), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n395), .B1(new_n618), .B2(new_n619), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT88), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n631), .B1(new_n642), .B2(new_n620), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT21), .B1(new_n643), .B2(new_n636), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n634), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n629), .B1(new_n635), .B2(G200), .ZN(new_n646));
  INV_X1    g0446(.A(G190), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(new_n635), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n610), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n476), .A2(new_n561), .A3(new_n564), .A4(new_n649), .ZN(G372));
  NAND2_X1  g0450(.A1(new_n518), .A2(new_n516), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n517), .A2(G169), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT92), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT26), .A4(new_n560), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n502), .A2(new_n560), .A3(new_n516), .A4(new_n518), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT92), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT90), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n557), .A2(new_n558), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n557), .B2(new_n558), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n556), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n544), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n553), .A2(new_n554), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n532), .A2(new_n541), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n657), .B1(new_n519), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n655), .A2(new_n658), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n535), .A2(new_n536), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n395), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n288), .B1(new_n673), .B2(new_n527), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n537), .A2(new_n540), .A3(new_n290), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT90), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n660), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n667), .B1(new_n677), .B2(new_n556), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n607), .A2(new_n608), .A3(new_n599), .A4(new_n593), .ZN(new_n679));
  AND4_X1   g0479(.A1(new_n519), .A2(new_n525), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT91), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n607), .A2(new_n608), .ZN(new_n682));
  INV_X1    g0482(.A(new_n604), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI211_X1 g0484(.A(KEYINPUT91), .B(new_n604), .C1(new_n607), .C2(new_n608), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n645), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n671), .A2(new_n687), .A3(new_n663), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n476), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n422), .A2(new_n427), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n449), .A2(new_n452), .A3(new_n463), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n348), .A3(new_n354), .A4(new_n353), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n471), .A2(new_n465), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n399), .A2(new_n402), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n357), .B1(new_n423), .B2(new_n696), .ZN(new_n697));
  AOI211_X1 g0497(.A(KEYINPUT18), .B(new_n695), .C1(new_n416), .C2(new_n417), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n323), .B1(new_n694), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(new_n314), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n689), .A2(new_n702), .ZN(G369));
  NAND2_X1  g0503(.A1(new_n639), .A2(new_n644), .ZN(new_n704));
  INV_X1    g0504(.A(new_n634), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n261), .A2(new_n222), .A3(G13), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G213), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G343), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n706), .A2(new_n629), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n629), .A2(new_n712), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n645), .A2(new_n648), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n682), .A2(new_n712), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n610), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n609), .A2(new_n712), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n684), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n609), .A2(new_n681), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n712), .B(KEYINPUT93), .Z(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n712), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n706), .A2(new_n610), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n723), .A2(new_n727), .A3(new_n729), .ZN(G399));
  NOR2_X1   g0530(.A1(new_n211), .A2(G41), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n548), .A2(G116), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n731), .A2(new_n261), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n219), .B2(new_n731), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT28), .Z(new_n736));
  INV_X1    g0536(.A(new_n609), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n645), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n680), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n519), .B2(new_n669), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n740), .B(new_n663), .C1(KEYINPUT26), .C2(new_n656), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT29), .B(new_n728), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n726), .ZN(new_n743));
  INV_X1    g0543(.A(new_n663), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(new_n680), .B2(new_n686), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n743), .B1(new_n745), .B2(new_n671), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n742), .B1(new_n746), .B2(KEYINPUT29), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n649), .A2(new_n561), .A3(new_n564), .A4(new_n726), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n598), .A2(new_n586), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n673), .A2(new_n527), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n749), .A2(new_n750), .A3(new_n631), .A4(new_n290), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n642), .A2(new_n620), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n751), .A2(new_n517), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n751), .A2(KEYINPUT30), .A3(new_n517), .A4(new_n752), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT94), .ZN(new_n757));
  INV_X1    g0557(.A(new_n592), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n517), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(new_n290), .A3(new_n750), .A4(new_n635), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n517), .A2(new_n757), .A3(new_n758), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n755), .B(new_n756), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n712), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT31), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n748), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n743), .A2(KEYINPUT31), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n755), .B1(new_n760), .B2(new_n761), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT95), .ZN(new_n769));
  INV_X1    g0569(.A(new_n756), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(new_n768), .B2(KEYINPUT95), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n767), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(G330), .B1(new_n766), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n747), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n736), .B1(new_n775), .B2(G1), .ZN(G364));
  AND2_X1   g0576(.A1(new_n222), .A2(G13), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n261), .B1(new_n777), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n731), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n718), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G330), .B2(new_n716), .ZN(new_n782));
  OAI21_X1  g0582(.A(G20), .B1(KEYINPUT97), .B2(G169), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(KEYINPUT97), .A2(G169), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n221), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n647), .A2(new_n317), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n222), .A2(new_n290), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G326), .A2(new_n791), .B1(new_n794), .B2(G311), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n222), .A2(G179), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n317), .A2(G190), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n789), .A2(new_n798), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  OAI221_X1 g0601(.A(new_n795), .B1(new_n796), .B2(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n647), .A2(G179), .A3(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n222), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n280), .B(new_n802), .C1(G294), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n789), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n807), .A2(new_n647), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G322), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n788), .A2(new_n797), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n617), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n797), .A2(new_n792), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(G329), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT98), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n799), .A2(new_n235), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n790), .A2(new_n457), .B1(new_n800), .B2(new_n229), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(G77), .C2(new_n794), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n805), .A2(G97), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n811), .A2(new_n231), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n279), .B(new_n821), .C1(G58), .C2(new_n808), .ZN(new_n822));
  INV_X1    g0622(.A(G159), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n813), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT32), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n819), .A2(new_n820), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n806), .A2(new_n815), .B1(new_n816), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n826), .A2(new_n816), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n787), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(G13), .A2(G33), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(G20), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n786), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n220), .A2(new_n263), .ZN(new_n835));
  INV_X1    g0635(.A(new_n530), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n210), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n257), .A2(G45), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT96), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n835), .B(new_n840), .C1(new_n839), .C2(new_n838), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n211), .A2(new_n279), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n842), .A2(G355), .B1(new_n569), .B2(new_n211), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n834), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n780), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n829), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n832), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n716), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n782), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  NOR2_X1   g0650(.A1(new_n355), .A2(new_n712), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n348), .A2(new_n712), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n352), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n851), .B1(new_n853), .B2(new_n355), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n746), .B(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n780), .B1(new_n855), .B2(new_n773), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n773), .B2(new_n855), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n280), .B1(G97), .B2(new_n805), .ZN(new_n858));
  INV_X1    g0658(.A(G311), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n811), .A2(new_n235), .B1(new_n813), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G303), .B2(new_n791), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n808), .A2(G294), .B1(G116), .B2(new_n794), .ZN(new_n862));
  INV_X1    g0662(.A(new_n800), .ZN(new_n863));
  INV_X1    g0663(.A(new_n799), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G283), .A2(new_n863), .B1(new_n864), .B2(G87), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n858), .A2(new_n861), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G150), .A2(new_n863), .B1(new_n794), .B2(G159), .ZN(new_n867));
  INV_X1    g0667(.A(G137), .ZN(new_n868));
  INV_X1    g0668(.A(G143), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n867), .B1(new_n868), .B2(new_n790), .C1(new_n869), .C2(new_n809), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT100), .Z(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT34), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n530), .B1(new_n811), .B2(new_n457), .ZN(new_n873));
  INV_X1    g0673(.A(G132), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n799), .A2(new_n229), .B1(new_n813), .B2(new_n874), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n873), .B(new_n875), .C1(G58), .C2(new_n805), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n871), .A2(KEYINPUT34), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n866), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n786), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n787), .A2(new_n831), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT99), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n845), .B1(new_n883), .B2(new_n203), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n880), .B(new_n884), .C1(new_n854), .C2(new_n831), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n857), .A2(new_n885), .ZN(G384));
  INV_X1    g0686(.A(new_n513), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n887), .A2(KEYINPUT35), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(KEYINPUT35), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(G116), .A3(new_n223), .A4(new_n889), .ZN(new_n890));
  XOR2_X1   g0690(.A(KEYINPUT101), .B(KEYINPUT36), .Z(new_n891));
  XNOR2_X1  g0691(.A(new_n890), .B(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n219), .B(G77), .C1(new_n361), .C2(new_n229), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n201), .A2(new_n229), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n261), .B(G13), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT104), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n411), .A2(new_n229), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n375), .B1(new_n898), .B2(new_n365), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n360), .B1(new_n899), .B2(new_n385), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n420), .B1(new_n900), .B2(new_n710), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n695), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n420), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n407), .A2(new_n710), .B1(new_n416), .B2(new_n417), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n900), .A2(new_n710), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n428), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT39), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT103), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  INV_X1    g0715(.A(new_n710), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n423), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n690), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n918), .B2(new_n699), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n905), .A2(new_n906), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n423), .B1(new_n696), .B2(new_n916), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT102), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n420), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n386), .A2(KEYINPUT102), .A3(new_n419), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n920), .B1(new_n925), .B2(KEYINPUT37), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n915), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n908), .A2(new_n910), .A3(KEYINPUT38), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n913), .A2(new_n914), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n914), .B1(new_n913), .B2(new_n930), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n471), .A2(new_n465), .A3(new_n728), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n688), .A2(new_n726), .A3(new_n854), .ZN(new_n935));
  INV_X1    g0735(.A(new_n851), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n465), .A2(new_n712), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n693), .A2(new_n691), .A3(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n465), .B(new_n712), .C1(new_n464), .C2(new_n471), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n935), .A2(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n911), .B2(new_n912), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n700), .A2(new_n710), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n897), .B1(new_n934), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n428), .A2(new_n909), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n412), .A2(new_n295), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT16), .B1(new_n383), .B2(new_n366), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n417), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n696), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n420), .C1(new_n710), .C2(new_n900), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n920), .B1(new_n951), .B2(KEYINPUT37), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n915), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n928), .B1(new_n953), .B2(new_n929), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT103), .B1(new_n945), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n933), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n913), .A2(new_n930), .A3(new_n914), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n958), .A2(KEYINPUT104), .A3(new_n942), .A4(new_n941), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n944), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n702), .B1(new_n475), .B2(new_n747), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n960), .B(new_n961), .Z(new_n962));
  NAND3_X1  g0762(.A1(new_n762), .A2(KEYINPUT31), .A3(new_n712), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n748), .A2(new_n765), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n938), .A2(new_n939), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n964), .A2(new_n965), .A3(KEYINPUT106), .A4(new_n854), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT40), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n927), .B2(new_n929), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n964), .A2(new_n965), .A3(new_n854), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT106), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n911), .A2(new_n912), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n967), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT105), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n969), .A2(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(KEYINPUT105), .B(new_n967), .C1(new_n970), .C2(new_n973), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n476), .A2(new_n964), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(G330), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n962), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n261), .B2(new_n777), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n962), .A2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n896), .B1(new_n984), .B2(new_n985), .ZN(G367));
  OAI211_X1 g0786(.A(new_n519), .B(new_n525), .C1(new_n522), .C2(new_n726), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n653), .A2(new_n743), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n645), .A2(new_n712), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n610), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n519), .B1(new_n987), .B2(new_n737), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n991), .A2(KEYINPUT42), .B1(new_n726), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(KEYINPUT42), .B2(new_n991), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n678), .B1(new_n552), .B2(new_n728), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n744), .A2(new_n665), .A3(new_n712), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n994), .A2(KEYINPUT43), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n987), .A2(new_n988), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n723), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n997), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n994), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n998), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1000), .B1(new_n998), .B2(new_n1005), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n731), .B(KEYINPUT41), .Z(new_n1009));
  NAND2_X1  g0809(.A1(new_n729), .A2(new_n727), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n999), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n999), .A3(KEYINPUT44), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT45), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1010), .B2(new_n999), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n989), .A2(new_n729), .A3(new_n727), .A4(KEYINPUT45), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1013), .A2(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(new_n723), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT107), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n729), .B1(new_n722), .B2(new_n990), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(new_n717), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n774), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1018), .A2(new_n723), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT107), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n1018), .B2(new_n723), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1020), .A2(new_n1023), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1009), .B1(new_n1027), .B2(new_n775), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1008), .B1(new_n1028), .B2(new_n779), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n244), .A2(new_n210), .A3(new_n836), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n833), .B1(new_n210), .B2(new_n338), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n780), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n793), .A2(new_n796), .B1(new_n799), .B2(new_n507), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n530), .B(new_n1033), .C1(G303), .C2(new_n808), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n811), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT46), .B1(new_n1035), .B2(G116), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G107), .B2(new_n805), .ZN(new_n1038));
  INV_X1    g0838(.A(G317), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n800), .A2(new_n587), .B1(new_n813), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G311), .B2(new_n791), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .A4(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G143), .A2(new_n791), .B1(new_n794), .B2(new_n201), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n805), .A2(G68), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n280), .A3(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G58), .A2(new_n1035), .B1(new_n814), .B2(G137), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT108), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(KEYINPUT108), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n800), .A2(new_n823), .B1(new_n799), .B2(new_n203), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G150), .B2(new_n808), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1042), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT47), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1032), .B1(new_n1053), .B2(new_n786), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n997), .B2(new_n847), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT109), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1029), .A2(new_n1056), .ZN(G387));
  INV_X1    g0857(.A(new_n1022), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n720), .A2(new_n721), .A3(new_n832), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n842), .A2(new_n733), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n249), .A2(new_n263), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n837), .ZN(new_n1062));
  OR3_X1    g0862(.A1(new_n301), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT50), .B1(new_n301), .B2(G50), .ZN(new_n1064));
  AOI21_X1  g0864(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1063), .A2(new_n732), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1062), .A2(new_n1066), .B1(new_n235), .B2(new_n211), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n780), .B1(new_n1067), .B2(new_n834), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n790), .A2(new_n823), .B1(new_n800), .B2(new_n301), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n836), .B(new_n1069), .C1(G97), .C2(new_n864), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n811), .A2(new_n203), .ZN(new_n1071));
  INV_X1    g0871(.A(G150), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n793), .A2(new_n229), .B1(new_n813), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(G50), .C2(new_n808), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n805), .A2(new_n339), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1070), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n790), .A2(new_n810), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n617), .A2(new_n793), .B1(new_n800), .B2(new_n859), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G317), .C2(new_n808), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1079), .A2(KEYINPUT48), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(KEYINPUT48), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n804), .A2(new_n796), .B1(new_n811), .B2(new_n587), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT49), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n530), .B1(new_n814), .B2(G326), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n569), .B2(new_n799), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT110), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1083), .A2(KEYINPUT49), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1076), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1068), .B1(new_n1090), .B2(new_n786), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1058), .A2(new_n779), .B1(new_n1059), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1023), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n731), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n775), .A2(new_n1058), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .ZN(G393));
  AND2_X1   g0896(.A1(new_n1018), .A2(new_n723), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1097), .A2(new_n1019), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n999), .A2(new_n832), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n254), .A2(new_n837), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n833), .B1(new_n507), .B2(new_n210), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n780), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n808), .A2(G159), .B1(new_n791), .B2(G150), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT112), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G68), .A2(new_n1035), .B1(new_n863), .B2(new_n201), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1108), .B1(new_n869), .B2(new_n813), .C1(new_n301), .C2(new_n793), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n530), .B1(new_n799), .B2(new_n231), .C1(new_n804), .C2(new_n203), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G294), .A2(new_n794), .B1(new_n863), .B2(G303), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n569), .B2(new_n804), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n808), .A2(G311), .B1(new_n791), .B2(G317), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT52), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n817), .B1(G283), .B2(new_n1035), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n810), .B2(new_n813), .ZN(new_n1118));
  NOR4_X1   g0918(.A1(new_n1114), .A2(new_n280), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1103), .B1(new_n1120), .B2(new_n786), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1099), .A2(new_n779), .B1(new_n1100), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1098), .A2(new_n1093), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n731), .A3(new_n1027), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(G390));
  INV_X1    g0925(.A(KEYINPUT114), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n940), .B2(new_n956), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n851), .B1(new_n746), .B2(new_n854), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n965), .ZN(new_n1129));
  OAI211_X1 g0929(.A(KEYINPUT114), .B(new_n933), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1127), .B(new_n1130), .C1(new_n931), .C2(new_n932), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n766), .A2(new_n772), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1132), .A2(G330), .A3(new_n854), .A4(new_n965), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n853), .A2(new_n355), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n728), .B(new_n1134), .C1(new_n739), .C2(new_n741), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n936), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n965), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n927), .A2(new_n929), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1137), .A2(new_n933), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1131), .A2(new_n1133), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n935), .A2(new_n936), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n956), .B1(new_n1142), .B2(new_n965), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n955), .A2(new_n957), .B1(new_n1143), .B2(KEYINPUT114), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1139), .B1(new_n1144), .B2(new_n1127), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n964), .A2(new_n965), .A3(G330), .A4(new_n854), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1141), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(G330), .B(new_n964), .C1(new_n473), .C2(new_n474), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(new_n702), .C1(new_n475), .C2(new_n747), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n854), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1129), .B1(new_n773), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1146), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1142), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n964), .A2(G330), .A3(new_n854), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1136), .B1(new_n1154), .B2(new_n1129), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1133), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1149), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1147), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1141), .B(new_n1157), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n731), .A3(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n779), .B(new_n1141), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n831), .B1(new_n955), .B2(new_n957), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n790), .A2(new_n796), .B1(new_n800), .B2(new_n235), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G294), .B2(new_n814), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n280), .B1(G77), .B2(new_n805), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n821), .B1(G68), .B2(new_n864), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n808), .A2(G116), .B1(G97), .B2(new_n794), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(G125), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n809), .A2(new_n874), .B1(new_n813), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G128), .B2(new_n791), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n811), .A2(new_n1072), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT115), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1172), .B(new_n1175), .C1(new_n793), .C2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G137), .A2(new_n863), .B1(new_n864), .B2(new_n201), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1179), .B(new_n280), .C1(new_n823), .C2(new_n804), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1169), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n786), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n780), .C1(new_n302), .C2(new_n882), .ZN(new_n1183));
  OR3_X1    g0983(.A1(new_n1163), .A2(KEYINPUT117), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT117), .B1(new_n1163), .B2(new_n1183), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1162), .A2(new_n1186), .A3(KEYINPUT118), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT118), .B1(new_n1162), .B2(new_n1186), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1161), .B1(new_n1188), .B2(new_n1189), .ZN(G378));
  NAND2_X1  g0990(.A1(new_n323), .A2(new_n312), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n311), .A2(new_n916), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1193), .B(new_n1194), .Z(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n976), .A2(G330), .A3(new_n977), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n974), .A2(new_n975), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n972), .A2(new_n966), .A3(new_n968), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1198), .A2(new_n1199), .A3(G330), .A4(new_n977), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1195), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1197), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n960), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n944), .A2(new_n1197), .A3(new_n1201), .A4(new_n959), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n779), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n780), .B1(new_n882), .B2(new_n201), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(G33), .A2(G41), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G50), .B(new_n1207), .C1(new_n836), .C2(new_n262), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n813), .A2(new_n796), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n790), .A2(new_n569), .B1(new_n800), .B2(new_n507), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G107), .C2(new_n808), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1071), .A2(G41), .A3(new_n530), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n794), .A2(new_n339), .B1(new_n864), .B2(G58), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(new_n1044), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT58), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1208), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n793), .A2(new_n868), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n790), .A2(new_n1170), .B1(new_n800), .B2(new_n874), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(G128), .C2(new_n808), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n1072), .B2(new_n804), .C1(new_n811), .C2(new_n1177), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT59), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n864), .A2(G159), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT119), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(G124), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(G124), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n814), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1221), .A2(new_n1222), .A3(new_n1226), .A4(new_n1207), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1220), .A2(KEYINPUT59), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1216), .B1(new_n1215), .B2(new_n1214), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1206), .B1(new_n1229), .B2(new_n786), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1196), .B2(new_n831), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1205), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1149), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1160), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1235), .A2(KEYINPUT57), .A3(new_n1204), .A4(new_n1203), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n731), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n944), .A2(new_n1197), .A3(new_n1201), .A4(new_n959), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1197), .A2(new_n1201), .B1(new_n944), .B2(new_n959), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1235), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1233), .B1(new_n1237), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT120), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT120), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n1233), .C1(new_n1237), .C2(new_n1241), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(G375));
  INV_X1    g1047(.A(new_n1009), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1152), .A2(new_n1142), .B1(new_n1155), .B2(new_n1133), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1149), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1158), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1129), .A2(new_n830), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n780), .B1(new_n882), .B2(G68), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n809), .A2(new_n796), .B1(new_n569), .B2(new_n800), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G107), .B2(new_n794), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n791), .A2(G294), .B1(new_n864), .B2(G77), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1255), .A2(new_n279), .A3(new_n1075), .A4(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n811), .A2(new_n507), .B1(new_n813), .B2(new_n617), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT121), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n808), .A2(G137), .B1(G128), .B2(new_n814), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n836), .B1(new_n864), .B2(G58), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1260), .B(new_n1261), .C1(new_n457), .C2(new_n804), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G132), .A2(new_n791), .B1(new_n1035), .B2(G159), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1263), .B1(new_n1072), .B2(new_n793), .C1(new_n800), .C2(new_n1177), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1257), .A2(new_n1259), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1253), .B1(new_n1265), .B2(new_n786), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT122), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1252), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1249), .B2(new_n778), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1251), .A2(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT123), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(G381));
  NAND2_X1  g1073(.A1(new_n1162), .A2(new_n1186), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT118), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n731), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1147), .B2(new_n1158), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1276), .A2(new_n1187), .B1(new_n1160), .B2(new_n1278), .ZN(new_n1279));
  OR4_X1    g1079(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(G381), .A2(G387), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1246), .A2(new_n1279), .A3(new_n1281), .ZN(G407));
  AOI21_X1  g1082(.A(G378), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n711), .A2(G213), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(KEYINPUT124), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(G213), .A3(G407), .ZN(G409));
  NAND3_X1  g1087(.A1(G387), .A2(new_n1124), .A3(new_n1122), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(G393), .B(new_n849), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1029), .A2(G390), .A3(new_n1056), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1289), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1029), .A2(G390), .A3(new_n1056), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G390), .B1(new_n1029), .B2(new_n1056), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1291), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT60), .B1(new_n1249), .B2(new_n1149), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1250), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1153), .A2(KEYINPUT60), .A3(new_n1149), .A4(new_n1156), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1299), .A2(new_n731), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G384), .B1(new_n1301), .B2(new_n1270), .ZN(new_n1302));
  INV_X1    g1102(.A(G384), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1303), .B(new_n1269), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT61), .B1(new_n1306), .B2(KEYINPUT62), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1299), .A2(new_n731), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n1250), .B2(new_n1297), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1303), .B1(new_n1309), .B2(new_n1269), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1301), .A2(G384), .A3(new_n1270), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1284), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(G2897), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1310), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1285), .A2(G2897), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT126), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1315), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1318), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT126), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1310), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1319), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT62), .B1(new_n1317), .B2(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(G378), .B(new_n1233), .C1(new_n1237), .C2(new_n1241), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1240), .A2(new_n1248), .A3(new_n1235), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1279), .B1(new_n1325), .B2(new_n1232), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1285), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1307), .B1(new_n1323), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1330));
  AND4_X1   g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1284), .A4(new_n1305), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1296), .B1(new_n1328), .B2(new_n1331), .ZN(new_n1332));
  OR2_X1    g1132(.A1(new_n1296), .A2(KEYINPUT61), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1305), .A2(KEYINPUT63), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1333), .B1(new_n1327), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1330), .A2(new_n1284), .ZN(new_n1336));
  NOR3_X1   g1136(.A1(new_n1314), .A2(new_n1316), .A3(KEYINPUT126), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1320), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1312), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1341));
  AOI21_X1  g1141(.A(KEYINPUT63), .B1(new_n1341), .B2(new_n1305), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1335), .B(new_n1340), .C1(new_n1342), .C2(KEYINPUT125), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1342), .A2(KEYINPUT125), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1332), .B1(new_n1343), .B2(new_n1344), .ZN(G405));
  AND2_X1   g1145(.A1(new_n1242), .A2(G378), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1283), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1305), .B1(new_n1291), .B2(new_n1295), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT127), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1291), .A2(new_n1305), .A3(new_n1295), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1349), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1351), .ZN(new_n1353));
  OAI21_X1  g1153(.A(KEYINPUT127), .B1(new_n1353), .B2(new_n1348), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1352), .A2(new_n1354), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1347), .B(new_n1355), .ZN(G402));
endmodule


