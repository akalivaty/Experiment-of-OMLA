

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592;

  XOR2_X1 U325 ( .A(G183GAT), .B(KEYINPUT18), .Z(n293) );
  XOR2_X1 U326 ( .A(KEYINPUT25), .B(n398), .Z(n294) );
  XNOR2_X1 U327 ( .A(n428), .B(KEYINPUT74), .ZN(n429) );
  XNOR2_X1 U328 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n384) );
  XNOR2_X1 U329 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U330 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U331 ( .A(n450), .B(n449), .ZN(n483) );
  NOR2_X1 U332 ( .A1(n502), .A2(n517), .ZN(n452) );
  INV_X1 U333 ( .A(G190GAT), .ZN(n480) );
  XNOR2_X1 U334 ( .A(n480), .B(KEYINPUT58), .ZN(n481) );
  XNOR2_X1 U335 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U336 ( .A(n482), .B(n481), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(G211GAT), .B(G155GAT), .Z(n296) );
  XNOR2_X1 U338 ( .A(G183GAT), .B(G127GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n298) );
  XOR2_X1 U340 ( .A(G22GAT), .B(G78GAT), .Z(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n315) );
  XOR2_X1 U342 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n300) );
  XNOR2_X1 U343 ( .A(G57GAT), .B(KEYINPUT15), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U345 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n302) );
  XNOR2_X1 U346 ( .A(KEYINPUT85), .B(KEYINPUT12), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U349 ( .A(G64GAT), .B(G15GAT), .Z(n306) );
  XNOR2_X1 U350 ( .A(G8GAT), .B(G1GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U353 ( .A(n309), .B(KEYINPUT83), .Z(n313) );
  XOR2_X1 U354 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n311) );
  XNOR2_X1 U355 ( .A(G71GAT), .B(KEYINPUT73), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n444) );
  XNOR2_X1 U357 ( .A(n444), .B(KEYINPUT82), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U359 ( .A(n315), .B(n314), .ZN(n317) );
  NAND2_X1 U360 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U361 ( .A(n317), .B(n316), .ZN(n586) );
  INV_X1 U362 ( .A(n586), .ZN(n570) );
  XOR2_X1 U363 ( .A(G162GAT), .B(G134GAT), .Z(n319) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(G29GAT), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n334) );
  XOR2_X1 U366 ( .A(G190GAT), .B(KEYINPUT80), .Z(n387) );
  XOR2_X1 U367 ( .A(G92GAT), .B(G106GAT), .Z(n321) );
  XNOR2_X1 U368 ( .A(G36GAT), .B(G218GAT), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U370 ( .A(n387), .B(n322), .Z(n324) );
  NAND2_X1 U371 ( .A1(G232GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U373 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n326) );
  XNOR2_X1 U374 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U376 ( .A(n328), .B(n327), .Z(n332) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n329), .B(KEYINPUT8), .ZN(n421) );
  XNOR2_X1 U379 ( .A(G99GAT), .B(G85GAT), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n330), .B(KEYINPUT75), .ZN(n430) );
  XNOR2_X1 U381 ( .A(n421), .B(n430), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n334), .B(n333), .ZN(n485) );
  INV_X1 U384 ( .A(n485), .ZN(n560) );
  XNOR2_X1 U385 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n560), .B(n335), .ZN(n590) );
  XOR2_X1 U387 ( .A(G120GAT), .B(G57GAT), .Z(n431) );
  XOR2_X1 U388 ( .A(n431), .B(G85GAT), .Z(n338) );
  XNOR2_X1 U389 ( .A(G29GAT), .B(G113GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n336), .B(G1GAT), .ZN(n413) );
  XNOR2_X1 U391 ( .A(G141GAT), .B(n413), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n343) );
  XNOR2_X1 U393 ( .A(G134GAT), .B(G127GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n339), .B(KEYINPUT0), .ZN(n368) );
  XOR2_X1 U395 ( .A(n368), .B(KEYINPUT6), .Z(n341) );
  NAND2_X1 U396 ( .A1(G225GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U398 ( .A(n343), .B(n342), .Z(n352) );
  XOR2_X1 U399 ( .A(KEYINPUT2), .B(G162GAT), .Z(n345) );
  XNOR2_X1 U400 ( .A(G155GAT), .B(G148GAT), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U402 ( .A(KEYINPUT3), .B(n346), .ZN(n366) );
  INV_X1 U403 ( .A(n366), .ZN(n350) );
  XOR2_X1 U404 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n348) );
  XNOR2_X1 U405 ( .A(KEYINPUT1), .B(KEYINPUT93), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n404) );
  XOR2_X1 U409 ( .A(KEYINPUT91), .B(KEYINPUT23), .Z(n355) );
  XNOR2_X1 U410 ( .A(G50GAT), .B(G22GAT), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n353), .B(G141GAT), .ZN(n416) );
  XOR2_X1 U412 ( .A(G106GAT), .B(G78GAT), .Z(n432) );
  XNOR2_X1 U413 ( .A(n416), .B(n432), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U415 ( .A(KEYINPUT92), .B(KEYINPUT22), .Z(n357) );
  NAND2_X1 U416 ( .A1(G228GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n359), .B(n358), .Z(n365) );
  XNOR2_X1 U419 ( .A(G211GAT), .B(G218GAT), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n360), .B(KEYINPUT21), .ZN(n361) );
  XOR2_X1 U421 ( .A(n361), .B(KEYINPUT90), .Z(n363) );
  XNOR2_X1 U422 ( .A(G197GAT), .B(G204GAT), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n393) );
  XNOR2_X1 U424 ( .A(n393), .B(KEYINPUT24), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n477) );
  XOR2_X1 U427 ( .A(n368), .B(G190GAT), .Z(n370) );
  NAND2_X1 U428 ( .A1(G227GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U430 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n372) );
  XNOR2_X1 U431 ( .A(G113GAT), .B(G71GAT), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U433 ( .A(n374), .B(n373), .Z(n379) );
  XOR2_X1 U434 ( .A(G120GAT), .B(G176GAT), .Z(n376) );
  XNOR2_X1 U435 ( .A(G169GAT), .B(G99GAT), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U437 ( .A(G43GAT), .B(n377), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U439 ( .A(n380), .B(KEYINPUT20), .Z(n383) );
  XNOR2_X1 U440 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n293), .B(n381), .ZN(n385) );
  XNOR2_X1 U442 ( .A(G15GAT), .B(n385), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n399) );
  XOR2_X1 U444 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U445 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n389), .B(n388), .ZN(n391) );
  XNOR2_X1 U447 ( .A(G176GAT), .B(G92GAT), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n390), .B(G64GAT), .ZN(n443) );
  XOR2_X1 U449 ( .A(n391), .B(n443), .Z(n395) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(G36GAT), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n392), .B(G8GAT), .ZN(n415) );
  XNOR2_X1 U452 ( .A(n415), .B(n393), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n507) );
  NAND2_X1 U454 ( .A1(n399), .A2(n507), .ZN(n396) );
  XOR2_X1 U455 ( .A(KEYINPUT97), .B(n396), .Z(n397) );
  NAND2_X1 U456 ( .A1(n477), .A2(n397), .ZN(n398) );
  BUF_X1 U457 ( .A(n399), .Z(n537) );
  NOR2_X1 U458 ( .A1(n477), .A2(n537), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n400), .B(KEYINPUT26), .ZN(n577) );
  XNOR2_X1 U460 ( .A(n507), .B(KEYINPUT27), .ZN(n405) );
  NAND2_X1 U461 ( .A1(n577), .A2(n405), .ZN(n401) );
  NAND2_X1 U462 ( .A1(n294), .A2(n401), .ZN(n402) );
  XOR2_X1 U463 ( .A(KEYINPUT98), .B(n402), .Z(n403) );
  NOR2_X1 U464 ( .A1(n404), .A2(n403), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n477), .B(KEYINPUT28), .ZN(n536) );
  INV_X1 U466 ( .A(n536), .ZN(n523) );
  OR2_X1 U467 ( .A1(n537), .A2(n523), .ZN(n406) );
  XNOR2_X1 U468 ( .A(KEYINPUT94), .B(n404), .ZN(n527) );
  NAND2_X1 U469 ( .A1(n527), .A2(n405), .ZN(n533) );
  NOR2_X1 U470 ( .A1(n406), .A2(n533), .ZN(n407) );
  NOR2_X1 U471 ( .A1(n408), .A2(n407), .ZN(n489) );
  NOR2_X1 U472 ( .A1(n590), .A2(n489), .ZN(n409) );
  NAND2_X1 U473 ( .A1(n570), .A2(n409), .ZN(n410) );
  XOR2_X1 U474 ( .A(KEYINPUT37), .B(n410), .Z(n502) );
  XOR2_X1 U475 ( .A(G15GAT), .B(G197GAT), .Z(n412) );
  XNOR2_X1 U476 ( .A(KEYINPUT70), .B(KEYINPUT66), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U478 ( .A(n414), .B(n413), .Z(n418) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n427) );
  XOR2_X1 U481 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n420) );
  XNOR2_X1 U482 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n425) );
  XOR2_X1 U484 ( .A(n421), .B(KEYINPUT69), .Z(n423) );
  NAND2_X1 U485 ( .A1(G229GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U487 ( .A(n425), .B(n424), .Z(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n579) );
  INV_X1 U489 ( .A(KEYINPUT41), .ZN(n451) );
  AND2_X1 U490 ( .A1(G230GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n438) );
  INV_X1 U492 ( .A(n438), .ZN(n436) );
  XOR2_X1 U493 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n434) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n437) );
  INV_X1 U496 ( .A(n437), .ZN(n435) );
  NAND2_X1 U497 ( .A1(n436), .A2(n435), .ZN(n440) );
  NAND2_X1 U498 ( .A1(n438), .A2(n437), .ZN(n439) );
  NAND2_X1 U499 ( .A1(n440), .A2(n439), .ZN(n442) );
  XOR2_X1 U500 ( .A(G148GAT), .B(G204GAT), .Z(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n450) );
  XOR2_X1 U502 ( .A(n444), .B(n443), .Z(n448) );
  XOR2_X1 U503 ( .A(KEYINPUT78), .B(KEYINPUT33), .Z(n446) );
  XNOR2_X1 U504 ( .A(KEYINPUT31), .B(KEYINPUT76), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n451), .B(n483), .ZN(n457) );
  OR2_X1 U507 ( .A1(n579), .A2(n457), .ZN(n517) );
  XOR2_X1 U508 ( .A(KEYINPUT109), .B(n452), .Z(n530) );
  NAND2_X1 U509 ( .A1(n530), .A2(n523), .ZN(n456) );
  XOR2_X1 U510 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n454) );
  XNOR2_X1 U511 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n453) );
  XNOR2_X1 U512 ( .A(n456), .B(n455), .ZN(G1339GAT) );
  XOR2_X1 U513 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n460) );
  INV_X1 U514 ( .A(n457), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n458), .A2(n579), .ZN(n459) );
  XOR2_X1 U516 ( .A(n460), .B(n459), .Z(n461) );
  NOR2_X1 U517 ( .A1(n586), .A2(n461), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT114), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n463), .A2(n485), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n464), .B(KEYINPUT115), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT47), .ZN(n471) );
  XOR2_X1 U522 ( .A(KEYINPUT71), .B(n579), .Z(n539) );
  NOR2_X1 U523 ( .A1(n590), .A2(n570), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT45), .ZN(n467) );
  XNOR2_X1 U525 ( .A(KEYINPUT65), .B(n467), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n539), .A2(n468), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n469), .A2(n483), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n473) );
  INV_X1 U529 ( .A(KEYINPUT48), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n473), .B(n472), .ZN(n534) );
  XOR2_X1 U531 ( .A(KEYINPUT122), .B(n507), .Z(n474) );
  NOR2_X1 U532 ( .A1(n534), .A2(n474), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT54), .B(n475), .Z(n476) );
  NOR2_X1 U534 ( .A1(n527), .A2(n476), .ZN(n578) );
  NAND2_X1 U535 ( .A1(n477), .A2(n578), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT55), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n479), .A2(n537), .ZN(n569) );
  NOR2_X1 U538 ( .A1(n485), .A2(n569), .ZN(n482) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n491) );
  INV_X1 U540 ( .A(n483), .ZN(n582) );
  INV_X1 U541 ( .A(n539), .ZN(n563) );
  NOR2_X1 U542 ( .A1(n582), .A2(n563), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(KEYINPUT79), .ZN(n501) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(KEYINPUT87), .Z(n487) );
  NAND2_X1 U545 ( .A1(n586), .A2(n485), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  OR2_X1 U547 ( .A1(n489), .A2(n488), .ZN(n516) );
  NOR2_X1 U548 ( .A1(n501), .A2(n516), .ZN(n497) );
  NAND2_X1 U549 ( .A1(n497), .A2(n527), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n497), .A2(n507), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U554 ( .A1(n497), .A2(n537), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n496) );
  XOR2_X1 U556 ( .A(G15GAT), .B(KEYINPUT99), .Z(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n499) );
  NAND2_X1 U559 ( .A1(n497), .A2(n523), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(n500), .ZN(G1327GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT39), .B(KEYINPUT104), .Z(n505) );
  NOR2_X1 U563 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U564 ( .A(KEYINPUT38), .B(n503), .ZN(n513) );
  NAND2_X1 U565 ( .A1(n513), .A2(n527), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(n506), .ZN(G1328GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n509) );
  NAND2_X1 U569 ( .A1(n507), .A2(n513), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U571 ( .A(G36GAT), .B(n510), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n513), .A2(n537), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(KEYINPUT40), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G43GAT), .B(n512), .ZN(G1330GAT) );
  XOR2_X1 U575 ( .A(G50GAT), .B(KEYINPUT107), .Z(n515) );
  NAND2_X1 U576 ( .A1(n523), .A2(n513), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n515), .B(n514), .ZN(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n519) );
  NOR2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n524), .A2(n527), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U582 ( .A(G57GAT), .B(n520), .Z(G1332GAT) );
  NAND2_X1 U583 ( .A1(n524), .A2(n507), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n521), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U585 ( .A1(n524), .A2(n537), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .Z(n526) );
  NAND2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NAND2_X1 U590 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n530), .A2(n507), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n530), .A2(n537), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(KEYINPUT110), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G99GAT), .B(n532), .ZN(G1338GAT) );
  XOR2_X1 U597 ( .A(G113GAT), .B(KEYINPUT117), .Z(n541) );
  NOR2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(n535), .Z(n551) );
  NAND2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U601 ( .A1(n551), .A2(n538), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n548), .A2(n539), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n543) );
  NAND2_X1 U605 ( .A1(n548), .A2(n458), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n546) );
  NAND2_X1 U609 ( .A1(n548), .A2(n586), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U613 ( .A1(n548), .A2(n560), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT120), .ZN(n554) );
  INV_X1 U616 ( .A(n577), .ZN(n552) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n561), .A2(n579), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U621 ( .A1(n561), .A2(n458), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U625 ( .A1(n561), .A2(n586), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n569), .ZN(n564) );
  XOR2_X1 U630 ( .A(G169GAT), .B(n564), .Z(G1348GAT) );
  NOR2_X1 U631 ( .A1(n569), .A2(n457), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n566) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  INV_X1 U636 ( .A(KEYINPUT124), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G183GAT), .B(n573), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(n576), .Z(n581) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n589) );
  INV_X1 U645 ( .A(n589), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n587), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U649 ( .A1(n587), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U651 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

