//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1251, new_n1252, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT66), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n205), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT64), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(new_n205), .B2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G13), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n222), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT65), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n213), .B(new_n219), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT67), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n228), .B(new_n230), .C1(new_n227), .C2(new_n226), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT68), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  OAI21_X1  g0047(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G150), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n217), .A2(G33), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n248), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n216), .ZN(new_n255));
  INV_X1    g0055(.A(G50), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n253), .A2(new_n255), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n258), .A2(new_n216), .A3(new_n254), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(KEYINPUT70), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n262), .B(new_n263), .C1(G1), .C2(new_n217), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n260), .B1(new_n264), .B2(new_n256), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  OAI211_X1 g0067(.A(G1), .B(G13), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n266), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n273), .A2(G223), .B1(new_n276), .B2(G77), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n271), .A2(new_n272), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G222), .A3(new_n269), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n268), .B1(new_n280), .B2(KEYINPUT69), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(KEYINPUT69), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(new_n268), .A3(G274), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n268), .A2(new_n283), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(G226), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n265), .B1(new_n290), .B2(G169), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(new_n290), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(G190), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n265), .B(KEYINPUT9), .ZN(new_n295));
  INV_X1    g0095(.A(G200), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n294), .B(new_n295), .C1(new_n296), .C2(new_n290), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n293), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G223), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n269), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n278), .B(new_n302), .C1(G226), .C2(new_n269), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G87), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n268), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G232), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n285), .B1(new_n287), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G179), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n308), .ZN(new_n311));
  INV_X1    g0111(.A(G68), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n271), .A2(new_n217), .A3(new_n272), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT7), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n217), .A4(new_n272), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G58), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n312), .ZN(new_n320));
  OAI21_X1  g0120(.A(G20), .B1(new_n320), .B2(new_n201), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n249), .A2(G159), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(KEYINPUT16), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n255), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n315), .A2(KEYINPUT75), .A3(new_n316), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n316), .A2(KEYINPUT75), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(G68), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT76), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n327), .A2(new_n328), .A3(new_n331), .A4(G68), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n324), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT16), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n326), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n251), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(new_n259), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n264), .B2(new_n336), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n311), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT18), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT18), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n311), .C1(new_n335), .C2(new_n338), .ZN(new_n342));
  INV_X1    g0142(.A(new_n338), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n308), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(G200), .B2(new_n308), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n323), .B1(new_n329), .B2(KEYINPUT76), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT16), .B1(new_n347), .B2(new_n332), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n343), .B(new_n346), .C1(new_n348), .C2(new_n326), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT17), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n333), .A2(new_n334), .ZN(new_n352));
  INV_X1    g0152(.A(new_n326), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n354), .A2(KEYINPUT17), .A3(new_n343), .A4(new_n346), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n340), .A2(new_n342), .A3(new_n351), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n306), .A2(G1698), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G226), .B2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n358), .B1(new_n360), .B2(new_n276), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n268), .A2(G238), .A3(new_n283), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n285), .A2(new_n364), .A3(KEYINPUT73), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT73), .B1(new_n285), .B2(new_n364), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT13), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n363), .B(new_n369), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G200), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n259), .A2(new_n312), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT12), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n249), .A2(G50), .B1(G20), .B2(new_n312), .ZN(new_n375));
  INV_X1    g0175(.A(G77), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n252), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n261), .B(G68), .C1(G1), .C2(new_n217), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT11), .B1(new_n377), .B2(new_n255), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n368), .A2(G190), .A3(new_n370), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n372), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(KEYINPUT74), .A2(G169), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n368), .B2(new_n370), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT14), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n388), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n368), .A2(G179), .A3(new_n370), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n382), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n385), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n288), .A2(G244), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n273), .A2(G238), .B1(new_n276), .B2(G107), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n278), .A2(G232), .A3(new_n269), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n286), .B(new_n395), .C1(new_n398), .C2(new_n362), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n292), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n261), .B(G77), .C1(G1), .C2(new_n217), .ZN(new_n401));
  XOR2_X1   g0201(.A(new_n401), .B(KEYINPUT72), .Z(new_n402));
  AOI22_X1  g0202(.A1(new_n336), .A2(new_n249), .B1(G20), .B2(G77), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT15), .B(G87), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n252), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n255), .B1(new_n376), .B2(new_n259), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n400), .B(new_n407), .C1(G169), .C2(new_n399), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n399), .A2(G190), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT71), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n399), .A2(KEYINPUT71), .A3(G190), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n399), .A2(new_n296), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n407), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n409), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n300), .A2(new_n357), .A3(new_n394), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n258), .A2(G107), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT85), .B(KEYINPUT25), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n257), .A2(G33), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n258), .A2(new_n423), .A3(new_n216), .A4(new_n254), .ZN(new_n424));
  INV_X1    g0224(.A(G107), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(G20), .B1(new_n271), .B2(new_n272), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT22), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(G87), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n217), .B(G87), .C1(new_n274), .C2(new_n275), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT22), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G116), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(G20), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT23), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n217), .B2(G107), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n425), .A2(KEYINPUT23), .A3(G20), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT24), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT24), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n434), .A2(new_n443), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n428), .B1(new_n445), .B2(new_n255), .ZN(new_n446));
  OAI211_X1 g0246(.A(G250), .B(new_n269), .C1(new_n274), .C2(new_n275), .ZN(new_n447));
  OAI211_X1 g0247(.A(G257), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G294), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT86), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT86), .A4(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n454), .A2(KEYINPUT87), .A3(new_n362), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  AND2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(G264), .A3(new_n268), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(new_n268), .A3(G274), .A4(new_n457), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n455), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n268), .B1(new_n452), .B2(new_n453), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(KEYINPUT87), .ZN(new_n468));
  OAI21_X1  g0268(.A(G169), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n454), .A2(new_n362), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G179), .A3(new_n465), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n446), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n444), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n443), .B1(new_n434), .B2(new_n440), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n255), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n427), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT87), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n464), .B1(new_n467), .B2(KEYINPUT87), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n344), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n470), .A2(new_n465), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n296), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n476), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n472), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G283), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n266), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n273), .B2(G250), .ZN(new_n487));
  OAI211_X1 g0287(.A(G244), .B(new_n269), .C1(new_n274), .C2(new_n275), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n269), .A2(KEYINPUT4), .A3(G244), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT79), .B1(new_n276), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n491), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT79), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n278), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n487), .A2(new_n490), .A3(new_n492), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n362), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n460), .A2(G257), .A3(new_n268), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n463), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT80), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n499), .B1(new_n496), .B2(new_n362), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(G200), .A3(new_n505), .ZN(new_n506));
  AOI211_X1 g0306(.A(new_n344), .B(new_n499), .C1(new_n496), .C2(new_n362), .ZN(new_n507));
  INV_X1    g0307(.A(new_n255), .ZN(new_n508));
  XOR2_X1   g0308(.A(KEYINPUT77), .B(KEYINPUT6), .Z(new_n509));
  XNOR2_X1  g0309(.A(G97), .B(G107), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G97), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT78), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT78), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G97), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g0316(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n425), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(G20), .B1(G77), .B2(new_n249), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n327), .A2(G107), .A3(new_n328), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n508), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n259), .A2(new_n512), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n424), .B2(new_n512), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n507), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n503), .A2(G179), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n310), .B2(new_n503), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n520), .A2(new_n521), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n255), .ZN(new_n529));
  INV_X1    g0329(.A(new_n524), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n506), .A2(new_n525), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G257), .B(new_n269), .C1(new_n274), .C2(new_n275), .ZN(new_n533));
  INV_X1    g0333(.A(G303), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n274), .A2(new_n275), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT83), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n278), .A2(KEYINPUT83), .A3(G257), .A4(new_n269), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT84), .B1(new_n273), .B2(G264), .ZN(new_n539));
  OAI211_X1 g0339(.A(G264), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT84), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n362), .ZN(new_n544));
  MUX2_X1   g0344(.A(new_n258), .B(new_n424), .S(G116), .Z(new_n545));
  INV_X1    g0345(.A(G116), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n254), .A2(new_n216), .B1(G20), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(G33), .B1(new_n513), .B2(new_n515), .ZN(new_n548));
  AOI21_X1  g0348(.A(G20), .B1(G33), .B2(G283), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(KEYINPUT20), .B(new_n547), .C1(new_n548), .C2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g0352(.A(KEYINPUT78), .B(G97), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n553), .B2(G33), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT20), .B1(new_n554), .B2(new_n547), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n545), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n460), .A2(G270), .A3(new_n268), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n463), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n292), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n544), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(G169), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n558), .B1(new_n543), .B2(new_n362), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT21), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n558), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n544), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT21), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT20), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n550), .B1(new_n516), .B2(new_n266), .ZN(new_n569));
  INV_X1    g0369(.A(new_n547), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n551), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n310), .B1(new_n572), .B2(new_n545), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n561), .B1(new_n564), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n556), .B1(new_n566), .B2(G200), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n344), .B2(new_n566), .ZN(new_n577));
  INV_X1    g0377(.A(new_n404), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(new_n258), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G87), .A2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n513), .A2(new_n515), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n217), .B1(new_n358), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(G68), .A2(new_n429), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n252), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n516), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT81), .B1(new_n586), .B2(new_n582), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT81), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n588), .B(KEYINPUT19), .C1(new_n516), .C2(new_n585), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n584), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n579), .B1(new_n590), .B2(new_n255), .ZN(new_n591));
  OAI211_X1 g0391(.A(G244), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n592));
  OAI211_X1 g0392(.A(G238), .B(new_n269), .C1(new_n274), .C2(new_n275), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(new_n435), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n362), .ZN(new_n595));
  INV_X1    g0395(.A(G274), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n362), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(G250), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n457), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n597), .A2(new_n457), .B1(new_n268), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G200), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n261), .A2(G87), .A3(new_n423), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n595), .A2(new_n600), .A3(G190), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n591), .A2(new_n602), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n579), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n261), .A2(new_n578), .A3(KEYINPUT82), .A4(new_n423), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT82), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n424), .B2(new_n404), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n581), .A2(new_n583), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n217), .B(G68), .C1(new_n274), .C2(new_n275), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n582), .B1(new_n553), .B2(new_n252), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n588), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n586), .A2(KEYINPUT81), .A3(new_n582), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n606), .B(new_n610), .C1(new_n617), .C2(new_n508), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n601), .A2(new_n310), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n595), .A2(new_n600), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n292), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n605), .A2(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n532), .A2(new_n575), .A3(new_n577), .A4(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n419), .A2(new_n484), .A3(new_n624), .ZN(G372));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n621), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n595), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n594), .A2(KEYINPUT88), .A3(new_n362), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(G169), .B1(new_n631), .B2(new_n600), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n480), .A2(new_n482), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n446), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n606), .B(new_n603), .C1(new_n617), .C2(new_n508), .ZN(new_n637));
  INV_X1    g0437(.A(new_n604), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n631), .A2(new_n600), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G200), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n627), .A2(new_n633), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n532), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n564), .A2(new_n574), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n560), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n472), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n634), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n503), .A2(new_n310), .ZN(new_n648));
  AOI211_X1 g0448(.A(new_n292), .B(new_n499), .C1(new_n496), .C2(new_n362), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT89), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n526), .B(new_n651), .C1(new_n310), .C2(new_n503), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n652), .A3(new_n531), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n642), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n605), .A2(new_n622), .ZN(new_n657));
  OAI22_X1  g0457(.A1(new_n648), .A2(new_n649), .B1(new_n522), .B2(new_n524), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n647), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n419), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n390), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n391), .B1(new_n387), .B2(new_n388), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n393), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n408), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n355), .A2(new_n351), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n384), .ZN(new_n668));
  INV_X1    g0468(.A(new_n342), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n343), .B1(new_n348), .B2(new_n326), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n341), .B1(new_n670), .B2(new_n311), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n298), .A2(new_n299), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n293), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n662), .A2(new_n675), .ZN(G369));
  NAND3_X1  g0476(.A1(new_n257), .A2(new_n217), .A3(G13), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT90), .Z(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n484), .B1(new_n446), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n472), .A2(new_n684), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n684), .A2(new_n556), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n645), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n575), .A2(new_n577), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n575), .A2(new_n684), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n484), .A2(new_n697), .B1(new_n472), .B2(new_n685), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(G399));
  NOR2_X1   g0499(.A1(new_n581), .A2(G116), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT91), .Z(new_n701));
  INV_X1    g0501(.A(new_n224), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n701), .A2(new_n257), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n215), .B2(new_n703), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  NAND2_X1  g0506(.A1(new_n661), .A2(new_n685), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n591), .A2(new_n603), .A3(new_n604), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n296), .B1(new_n631), .B2(new_n600), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n710), .A2(new_n711), .B1(new_n626), .B2(new_n632), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n653), .A2(new_n712), .A3(new_n655), .ZN(new_n713));
  INV_X1    g0513(.A(new_n658), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT26), .B1(new_n623), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n685), .B1(new_n647), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n709), .B1(new_n708), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G330), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n575), .A2(new_n623), .A3(new_n577), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n484), .A3(new_n532), .A4(new_n685), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT93), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n624), .A2(KEYINPUT93), .A3(new_n484), .A4(new_n685), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n461), .A2(new_n557), .A3(new_n463), .A4(G179), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n543), .B2(new_n362), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n470), .A3(new_n503), .A4(new_n620), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n481), .A2(new_n566), .A3(new_n292), .A4(new_n501), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n631), .A2(KEYINPUT92), .A3(new_n600), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT92), .B1(new_n631), .B2(new_n600), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n684), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT31), .B(new_n684), .C1(new_n730), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n719), .B1(new_n725), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n718), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n706), .B1(new_n744), .B2(G1), .ZN(G364));
  NOR2_X1   g0545(.A1(new_n222), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n257), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n703), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n224), .A2(G116), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n224), .A2(G355), .A3(new_n278), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n243), .A2(new_n456), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n224), .A2(new_n276), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n456), .B2(new_n215), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n750), .B(new_n751), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n216), .B1(G20), .B2(new_n310), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT94), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n749), .B1(new_n755), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT95), .Z(new_n763));
  INV_X1    g0563(.A(new_n759), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n217), .A2(new_n292), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n344), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n766), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(KEYINPUT33), .A2(G317), .ZN(new_n773));
  NAND2_X1  g0573(.A1(KEYINPUT33), .A2(G317), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n344), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n217), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n770), .B(new_n775), .C1(G294), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n217), .A2(G190), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(new_n292), .A3(new_n296), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(new_n765), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n784), .A2(new_n344), .A3(G200), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n278), .B(new_n788), .C1(G322), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n292), .A2(G200), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT96), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n792), .A2(new_n217), .A3(G190), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G283), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n792), .A2(new_n217), .A3(new_n344), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G303), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n779), .A2(new_n790), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n777), .A2(new_n512), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n782), .A2(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(KEYINPUT32), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n798), .B(new_n800), .C1(G68), .C2(new_n771), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n278), .B1(new_n786), .B2(new_n376), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G58), .B2(new_n789), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n799), .A2(KEYINPUT32), .B1(G50), .B2(new_n767), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G87), .A2(new_n795), .B1(new_n793), .B2(G107), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n801), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n758), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n763), .B1(new_n764), .B2(new_n807), .C1(new_n693), .C2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT97), .Z(new_n810));
  NOR2_X1   g0610(.A1(new_n693), .A2(G330), .ZN(new_n811));
  INV_X1    g0611(.A(new_n694), .ZN(new_n812));
  INV_X1    g0612(.A(new_n703), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n811), .B(new_n812), .C1(new_n813), .C2(new_n747), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NOR2_X1   g0616(.A1(new_n408), .A2(new_n684), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n414), .A2(new_n416), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n684), .A2(new_n407), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n817), .B1(new_n820), .B2(new_n408), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n707), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n821), .B(new_n685), .C1(new_n647), .C2(new_n660), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n749), .B1(new_n825), .B2(new_n743), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n743), .B2(new_n825), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n764), .A2(new_n757), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n749), .B1(G77), .B2(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G137), .A2(new_n767), .B1(new_n771), .B2(G150), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT98), .Z(new_n831));
  INV_X1    g0631(.A(G143), .ZN(new_n832));
  INV_X1    g0632(.A(new_n789), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n831), .B1(new_n832), .B2(new_n833), .C1(new_n834), .C2(new_n786), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT34), .Z(new_n836));
  INV_X1    g0636(.A(new_n793), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n312), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n278), .B1(new_n781), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G58), .B2(new_n778), .ZN(new_n842));
  INV_X1    g0642(.A(new_n795), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n839), .B(new_n842), .C1(new_n256), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n798), .B1(G303), .B2(new_n767), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n485), .B2(new_n772), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n833), .A2(new_n847), .B1(new_n786), .B2(new_n546), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n278), .B(new_n848), .C1(G311), .C2(new_n782), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n793), .A2(G87), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n795), .A2(G107), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n836), .A2(new_n844), .B1(new_n846), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n829), .B1(new_n853), .B2(new_n759), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n757), .B2(new_n821), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n827), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT99), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  NOR2_X1   g0658(.A1(new_n746), .A2(new_n257), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n334), .B1(new_n317), .B2(new_n323), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n325), .A2(new_n255), .A3(new_n861), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n862), .A2(new_n338), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n681), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n672), .B2(new_n667), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n681), .B1(new_n335), .B2(new_n338), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n339), .A2(new_n866), .A3(new_n867), .A4(new_n349), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n311), .A2(new_n681), .B1(new_n862), .B2(new_n338), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n349), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n860), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n864), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n356), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(KEYINPUT39), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n339), .A2(new_n866), .A3(new_n349), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n880), .A2(new_n868), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n866), .B1(new_n672), .B2(new_n667), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n860), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n877), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n878), .B1(new_n885), .B2(KEYINPUT39), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n392), .A2(new_n393), .A3(new_n685), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n876), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n876), .B2(new_n872), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT101), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT101), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n874), .A2(new_n892), .A3(new_n877), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n665), .B(new_n384), .C1(new_n382), .C2(new_n685), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n393), .B(new_n684), .C1(new_n392), .C2(new_n385), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n817), .B(KEYINPUT100), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n824), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n682), .B1(new_n669), .B2(new_n671), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n888), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n675), .B1(new_n718), .B2(new_n418), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n903), .B(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n740), .B1(new_n723), .B2(new_n724), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n897), .A2(new_n821), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT40), .B1(new_n894), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n883), .B2(new_n877), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n909), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n418), .A2(new_n906), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n719), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n859), .B1(new_n905), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n905), .B2(new_n915), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n918), .A2(G116), .A3(new_n218), .A4(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT36), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n214), .A2(new_n376), .A3(new_n320), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n312), .A2(G50), .ZN(new_n923));
  OAI211_X1 g0723(.A(G1), .B(new_n222), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n917), .A2(new_n921), .A3(new_n924), .ZN(G367));
  XOR2_X1   g0725(.A(new_n703), .B(KEYINPUT41), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n654), .A2(new_n684), .ZN(new_n927));
  INV_X1    g0727(.A(new_n531), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n532), .B1(new_n928), .B2(new_n685), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n698), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT45), .Z(new_n932));
  NOR2_X1   g0732(.A1(new_n698), .A2(new_n930), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT44), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(new_n696), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n484), .A2(new_n697), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n937), .B1(new_n688), .B2(new_n697), .C1(new_n812), .C2(KEYINPUT105), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT105), .B1(new_n812), .B2(KEYINPUT104), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n938), .B(new_n939), .Z(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(new_n744), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n926), .B1(new_n941), .B2(new_n744), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n748), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n930), .A2(new_n472), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n685), .B1(new_n944), .B2(new_n714), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT42), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n930), .A2(new_n484), .A3(new_n697), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n945), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT102), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(KEYINPUT102), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(KEYINPUT42), .C2(new_n947), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n684), .A2(new_n637), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n642), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n634), .B2(new_n953), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n952), .A2(KEYINPUT43), .A3(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT103), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n955), .B(KEYINPUT43), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(KEYINPUT103), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n930), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n696), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n943), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n961), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n235), .A2(new_n753), .ZN(new_n967));
  INV_X1    g0767(.A(new_n761), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n224), .B2(new_n404), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n749), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(G317), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n833), .A2(new_n534), .B1(new_n781), .B2(new_n971), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n278), .B(new_n972), .C1(G283), .C2(new_n785), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n772), .A2(new_n847), .B1(new_n425), .B2(new_n777), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G311), .B2(new_n767), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n973), .B(new_n975), .C1(new_n553), .C2(new_n837), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT106), .B1(new_n843), .B2(new_n546), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT46), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n795), .A2(G58), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G50), .A2(new_n785), .B1(new_n789), .B2(G150), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n793), .A2(G77), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n276), .B1(new_n782), .B2(G137), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n777), .A2(new_n312), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n772), .B2(new_n834), .C1(new_n832), .C2(new_n768), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n976), .A2(new_n978), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n970), .B1(new_n988), .B2(new_n759), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n808), .B2(new_n955), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n966), .A2(new_n990), .ZN(G387));
  AOI22_X1  g0791(.A1(G303), .A2(new_n785), .B1(new_n789), .B2(G317), .ZN(new_n992));
  INV_X1    g0792(.A(G322), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n787), .B2(new_n772), .C1(new_n993), .C2(new_n768), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT48), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n485), .B2(new_n777), .C1(new_n847), .C2(new_n843), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n994), .A2(new_n995), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n999), .A2(KEYINPUT49), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(KEYINPUT49), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n276), .B1(new_n781), .B2(new_n769), .C1(new_n837), .C2(new_n546), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n795), .A2(G77), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n276), .B1(new_n782), .B2(G150), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n837), .C2(new_n512), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT107), .Z(new_n1007));
  NOR2_X1   g0807(.A1(new_n777), .A2(new_n404), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G50), .A2(new_n789), .B1(new_n785), .B2(G68), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n251), .B2(new_n772), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(G159), .C2(new_n767), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT108), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n759), .B1(new_n1003), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g0814(.A1(new_n239), .A2(new_n456), .A3(new_n278), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n251), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT50), .B1(new_n251), .B2(G50), .ZN(new_n1017));
  AOI21_X1  g0817(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n701), .B1(new_n276), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n224), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n968), .C1(new_n425), .C2(new_n224), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1014), .A2(new_n749), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n689), .B2(new_n758), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n940), .B2(new_n748), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n744), .A2(new_n940), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n703), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n744), .A2(new_n940), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(G393));
  INV_X1    g0829(.A(KEYINPUT109), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n936), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n935), .A2(KEYINPUT109), .A3(new_n695), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n1026), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT111), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n703), .A3(new_n941), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1033), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n962), .A2(new_n758), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n968), .B1(new_n224), .B2(new_n553), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n246), .A2(new_n753), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n749), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n789), .A2(G159), .B1(new_n767), .B2(G150), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT51), .Z(new_n1043));
  NAND2_X1  g0843(.A1(new_n778), .A2(G77), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n276), .B1(new_n782), .B2(G143), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n850), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1043), .B(new_n1046), .C1(new_n312), .C2(new_n843), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n336), .A2(new_n785), .B1(new_n771), .B2(G50), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT110), .Z(new_n1049));
  OAI22_X1  g0849(.A1(new_n485), .A2(new_n843), .B1(new_n837), .B2(new_n425), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n276), .B1(new_n993), .B2(new_n781), .C1(new_n786), .C2(new_n847), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n772), .A2(new_n534), .B1(new_n546), .B2(new_n777), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n789), .A2(G311), .B1(new_n767), .B2(G317), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1047), .A2(new_n1049), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1041), .B1(new_n1056), .B2(new_n759), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1037), .A2(new_n748), .B1(new_n1038), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1036), .A2(new_n1058), .ZN(G390));
  NAND3_X1  g0859(.A1(new_n742), .A2(new_n821), .A3(new_n897), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n820), .A2(new_n408), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n685), .B(new_n1061), .C1(new_n647), .C2(new_n716), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n817), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n897), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n887), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n883), .B2(new_n877), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1067), .A3(KEYINPUT112), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT112), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n866), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n356), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n880), .A2(new_n868), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT38), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n887), .B1(new_n889), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n898), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1069), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1068), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n878), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT39), .B1(new_n883), .B2(new_n877), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1078), .A2(new_n1079), .B1(new_n900), .B2(new_n1066), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(KEYINPUT113), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT113), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1077), .A2(new_n1083), .A3(new_n1080), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1060), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1083), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1086));
  NOR4_X1   g0886(.A1(new_n906), .A2(new_n719), .A3(new_n898), .A4(new_n822), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n886), .A2(new_n756), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n749), .B1(new_n336), .B2(new_n828), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n795), .A2(G87), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n278), .B1(new_n782), .B2(G294), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n516), .A2(new_n785), .B1(new_n789), .B2(G116), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1044), .B1(new_n772), .B2(new_n425), .C1(new_n485), .C2(new_n768), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1095), .A2(new_n1096), .A3(new_n838), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1098), .A2(KEYINPUT115), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n795), .A2(G150), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT53), .Z(new_n1101));
  INV_X1    g0901(.A(G128), .ZN(new_n1102));
  INV_X1    g0902(.A(G137), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1102), .A2(new_n768), .B1(new_n772), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G159), .B2(new_n778), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n278), .B1(new_n786), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n782), .A2(G125), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n833), .B2(new_n840), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1107), .B(new_n1109), .C1(G50), .C2(new_n793), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1101), .A2(new_n1105), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1098), .A2(KEYINPUT115), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1099), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1091), .B1(new_n1113), .B2(new_n759), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1089), .A2(new_n748), .B1(new_n1090), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n419), .A2(new_n742), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1116), .B(new_n675), .C1(new_n718), .C2(new_n418), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n824), .A2(new_n899), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n897), .B1(new_n742), .B2(new_n821), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n1087), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1121), .A2(KEYINPUT114), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT114), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1123), .B(new_n1119), .C1(new_n1120), .C2(new_n1087), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n725), .A2(new_n741), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(G330), .A3(new_n821), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n898), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1064), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1060), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1118), .B1(new_n1122), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1121), .A2(KEYINPUT114), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1117), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1077), .A2(new_n1083), .A3(new_n1080), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1087), .B1(new_n1136), .B2(new_n1086), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1082), .A2(new_n1060), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1132), .A2(new_n703), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1115), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT116), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1115), .A2(new_n1140), .A3(KEYINPUT116), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n265), .A2(new_n681), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n300), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n300), .A2(new_n1147), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OR3_X1    g0952(.A1(new_n1149), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT118), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT101), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n892), .B1(new_n874), .B2(new_n877), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n908), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n910), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n719), .B1(new_n911), .B2(new_n908), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1157), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n907), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1125), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT40), .B1(new_n889), .B2(new_n1073), .ZN(new_n1166));
  OAI21_X1  g0966(.A(G330), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n909), .A2(KEYINPUT118), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1156), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n903), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT118), .B1(new_n909), .B2(new_n1167), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1155), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1165), .B1(new_n891), .B2(new_n893), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1157), .B(new_n1162), .C1(new_n1174), .C2(KEYINPUT40), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1155), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1156), .B1(new_n1177), .B2(KEYINPUT118), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n903), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1156), .A2(new_n756), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n749), .B1(G50), .B2(new_n828), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n985), .B1(new_n546), .B2(new_n768), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n793), .A2(G58), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G41), .B(new_n278), .C1(new_n785), .C2(new_n578), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n789), .A2(G107), .B1(G283), .B2(new_n782), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1004), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1183), .B(new_n1187), .C1(G97), .C2(new_n771), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT117), .Z(new_n1189));
  INV_X1    g0989(.A(KEYINPUT58), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(G33), .A2(G41), .ZN(new_n1193));
  AOI211_X1 g0993(.A(G50), .B(new_n1193), .C1(new_n276), .C2(new_n267), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n833), .A2(new_n1102), .B1(new_n786), .B2(new_n1103), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G132), .B2(new_n771), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G150), .A2(new_n778), .B1(new_n767), .B2(G125), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n843), .C2(new_n1106), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n782), .A2(G124), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1193), .B(new_n1200), .C1(new_n837), .C2(new_n834), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1198), .B2(KEYINPUT59), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1194), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1191), .A2(new_n1192), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1182), .B1(new_n1204), .B2(new_n759), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1180), .A2(new_n748), .B1(new_n1181), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1139), .B2(new_n1118), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT119), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT119), .B1(new_n1211), .B2(new_n1170), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1208), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1118), .A2(new_n1139), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n703), .B1(new_n1215), .B2(KEYINPUT57), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1206), .B1(new_n1214), .B2(new_n1216), .ZN(G375));
  NOR2_X1   g1017(.A1(new_n1122), .A2(new_n1130), .ZN(new_n1218));
  OR3_X1    g1018(.A1(new_n1218), .A2(KEYINPUT121), .A3(new_n747), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n749), .B1(G68), .B2(new_n828), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n767), .A2(G132), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n256), .B2(new_n777), .C1(new_n772), .C2(new_n1106), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n795), .A2(G159), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n276), .B1(new_n789), .B2(G137), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n785), .A2(G150), .B1(G128), .B2(new_n782), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1184), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n795), .A2(G97), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n278), .B1(new_n785), .B2(G107), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n789), .A2(G283), .B1(G303), .B2(new_n782), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n981), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1008), .B1(G294), .B2(new_n767), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n546), .B2(new_n772), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1222), .A2(new_n1226), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1220), .B1(new_n1233), .B2(new_n759), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n897), .B2(new_n757), .ZN(new_n1235));
  OAI21_X1  g1035(.A(KEYINPUT121), .B1(new_n1218), .B2(new_n747), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1219), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1133), .A2(new_n1117), .A3(new_n1134), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT120), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT120), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1218), .A2(new_n1240), .A3(new_n1117), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1135), .A2(new_n926), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1237), .B1(new_n1242), .B2(new_n1243), .ZN(G381));
  OR3_X1    g1044(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1141), .ZN(new_n1247));
  INV_X1    g1047(.A(G375), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(G407));
  NAND2_X1  g1049(.A1(new_n683), .A2(G213), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT122), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1248), .A2(new_n1247), .A3(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G407), .A2(G213), .A3(new_n1252), .ZN(G409));
  INV_X1    g1053(.A(KEYINPUT123), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1251), .A2(G2897), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1238), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n813), .B1(new_n1256), .B2(KEYINPUT60), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1242), .B2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1237), .A2(new_n1259), .A3(G384), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G384), .B1(new_n1237), .B2(new_n1259), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1254), .B(new_n1255), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n683), .A2(G213), .A3(G2897), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1254), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1262), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1260), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1255), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1264), .B1(new_n1267), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1250), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1213), .B(new_n703), .C1(KEYINPUT57), .C2(new_n1215), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G378), .A2(new_n1273), .A3(new_n1206), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1181), .A2(new_n1205), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1139), .A2(new_n1118), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1180), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1277), .B2(new_n926), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1180), .A2(KEYINPUT119), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1212), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n747), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1247), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1272), .B1(new_n1274), .B2(new_n1282), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1271), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(G390), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G393), .B(new_n815), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT124), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(G387), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1286), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n966), .B2(new_n990), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1285), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1290), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT124), .B1(new_n966), .B2(new_n990), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1292), .B(G390), .C1(new_n1286), .C2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT61), .B1(new_n1291), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1282), .B1(G375), .B2(new_n1145), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1296), .A2(new_n1250), .A3(new_n1265), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1251), .B1(new_n1274), .B2(new_n1282), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1265), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1284), .A2(new_n1295), .A3(new_n1299), .A4(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1271), .B2(new_n1300), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1269), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1251), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1306), .A2(new_n1296), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1297), .A2(new_n1305), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT125), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1297), .A2(KEYINPUT125), .A3(new_n1305), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1304), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1302), .B1(new_n1313), .B2(new_n1314), .ZN(G405));
  OAI21_X1  g1115(.A(KEYINPUT126), .B1(new_n1248), .B2(new_n1141), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(G375), .A2(new_n1317), .A3(new_n1247), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1316), .A2(new_n1318), .A3(new_n1274), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT127), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1265), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1319), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1274), .A2(new_n1318), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1324), .A2(new_n1320), .A3(new_n1265), .A4(new_n1316), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1314), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1323), .A2(new_n1325), .A3(new_n1291), .A4(new_n1294), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(G402));
endmodule


