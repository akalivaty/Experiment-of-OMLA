

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777;

  XNOR2_X1 U375 ( .A(n464), .B(n463), .ZN(n758) );
  INV_X1 U376 ( .A(G125), .ZN(n433) );
  XNOR2_X1 U377 ( .A(n766), .B(n512), .ZN(n371) );
  XOR2_X1 U378 ( .A(n534), .B(n533), .Z(n353) );
  XNOR2_X2 U379 ( .A(n422), .B(KEYINPUT35), .ZN(n587) );
  AND2_X2 U380 ( .A1(n421), .A2(n418), .ZN(n354) );
  INV_X2 U381 ( .A(n507), .ZN(n534) );
  XNOR2_X2 U382 ( .A(G128), .B(G143), .ZN(n507) );
  XNOR2_X2 U383 ( .A(n571), .B(n570), .ZN(n680) );
  INV_X1 U384 ( .A(n606), .ZN(n712) );
  XNOR2_X1 U385 ( .A(n530), .B(n502), .ZN(n504) );
  AND2_X1 U386 ( .A1(n359), .A2(n357), .ZN(n356) );
  NOR2_X1 U387 ( .A1(n606), .A2(n586), .ZN(n671) );
  XNOR2_X1 U388 ( .A(n479), .B(n478), .ZN(n775) );
  NOR2_X1 U389 ( .A1(n630), .A2(n618), .ZN(n677) );
  XNOR2_X1 U390 ( .A(n610), .B(KEYINPUT79), .ZN(n569) );
  XNOR2_X1 U391 ( .A(n633), .B(n603), .ZN(n681) );
  XNOR2_X1 U392 ( .A(n470), .B(n468), .ZN(n575) );
  OR2_X1 U393 ( .A1(n656), .A2(G902), .ZN(n388) );
  XNOR2_X1 U394 ( .A(n500), .B(n499), .ZN(n503) );
  XOR2_X1 U395 ( .A(G122), .B(G113), .Z(n559) );
  XNOR2_X1 U396 ( .A(G128), .B(G143), .ZN(n355) );
  INV_X2 U397 ( .A(G116), .ZN(n467) );
  AND2_X2 U398 ( .A1(n426), .A2(n427), .ZN(n363) );
  OR2_X1 U399 ( .A1(n666), .A2(KEYINPUT103), .ZN(n417) );
  NOR2_X1 U400 ( .A1(n416), .A2(n415), .ZN(n414) );
  NOR2_X1 U401 ( .A1(n680), .A2(n417), .ZN(n416) );
  XNOR2_X2 U402 ( .A(n467), .B(G107), .ZN(n548) );
  OR2_X2 U403 ( .A1(n775), .A2(n671), .ZN(n588) );
  XNOR2_X1 U404 ( .A(n535), .B(n487), .ZN(n558) );
  INV_X1 U405 ( .A(KEYINPUT10), .ZN(n487) );
  AND2_X1 U406 ( .A1(n447), .A2(n681), .ZN(n637) );
  AND2_X1 U407 ( .A1(n604), .A2(n448), .ZN(n447) );
  INV_X1 U408 ( .A(n612), .ZN(n448) );
  INV_X1 U409 ( .A(n605), .ZN(n386) );
  NAND2_X1 U410 ( .A1(n710), .A2(n709), .ZN(n707) );
  XNOR2_X1 U411 ( .A(n476), .B(n475), .ZN(n547) );
  INV_X1 U412 ( .A(KEYINPUT8), .ZN(n475) );
  NAND2_X1 U413 ( .A1(n493), .A2(G234), .ZN(n476) );
  AND2_X2 U414 ( .A1(n655), .A2(n654), .ZN(n743) );
  XNOR2_X1 U415 ( .A(n637), .B(KEYINPUT108), .ZN(n387) );
  INV_X1 U416 ( .A(KEYINPUT36), .ZN(n385) );
  XNOR2_X1 U417 ( .A(n628), .B(n446), .ZN(n378) );
  NOR2_X1 U418 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U419 ( .A1(G953), .A2(G237), .ZN(n556) );
  XNOR2_X1 U420 ( .A(G140), .B(KEYINPUT11), .ZN(n560) );
  XNOR2_X1 U421 ( .A(KEYINPUT77), .B(G107), .ZN(n439) );
  NAND2_X1 U422 ( .A1(n354), .A2(n393), .ZN(n392) );
  XNOR2_X1 U423 ( .A(n712), .B(KEYINPUT6), .ZN(n581) );
  INV_X1 U424 ( .A(KEYINPUT34), .ZN(n428) );
  INV_X1 U425 ( .A(KEYINPUT30), .ZN(n442) );
  INV_X1 U426 ( .A(n607), .ZN(n408) );
  XNOR2_X1 U427 ( .A(n495), .B(n496), .ZN(n710) );
  BUF_X1 U428 ( .A(n581), .Z(n604) );
  INV_X1 U429 ( .A(G953), .ZN(n752) );
  XNOR2_X1 U430 ( .A(n492), .B(KEYINPUT24), .ZN(n482) );
  XNOR2_X1 U431 ( .A(G119), .B(G110), .ZN(n492) );
  XNOR2_X1 U432 ( .A(n558), .B(n488), .ZN(n764) );
  XOR2_X1 U433 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n550) );
  INV_X1 U434 ( .A(G134), .ZN(n508) );
  XNOR2_X1 U435 ( .A(n371), .B(n513), .ZN(n739) );
  XNOR2_X1 U436 ( .A(n529), .B(n559), .ZN(n463) );
  XNOR2_X1 U437 ( .A(n465), .B(n530), .ZN(n464) );
  XNOR2_X1 U438 ( .A(n548), .B(n466), .ZN(n465) );
  XNOR2_X1 U439 ( .A(n404), .B(n364), .ZN(n645) );
  NOR2_X1 U440 ( .A1(n386), .A2(n385), .ZN(n382) );
  AND2_X1 U441 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n544), .B(KEYINPUT19), .ZN(n545) );
  XNOR2_X1 U443 ( .A(n451), .B(n449), .ZN(n574) );
  XNOR2_X1 U444 ( .A(n568), .B(n450), .ZN(n449) );
  OR2_X1 U445 ( .A1(n744), .A2(G902), .ZN(n451) );
  INV_X1 U446 ( .A(G475), .ZN(n450) );
  XNOR2_X1 U447 ( .A(n553), .B(n469), .ZN(n468) );
  OR2_X1 U448 ( .A1(n745), .A2(G902), .ZN(n470) );
  INV_X1 U449 ( .A(G478), .ZN(n553) );
  XNOR2_X1 U450 ( .A(n580), .B(n579), .ZN(n584) );
  XNOR2_X1 U451 ( .A(KEYINPUT70), .B(KEYINPUT22), .ZN(n579) );
  INV_X1 U452 ( .A(KEYINPUT1), .ZN(n456) );
  BUF_X1 U453 ( .A(n710), .Z(n431) );
  NOR2_X2 U454 ( .A1(n584), .A2(n604), .ZN(n409) );
  XNOR2_X1 U455 ( .A(n454), .B(n366), .ZN(n453) );
  NAND2_X1 U456 ( .A1(n743), .A2(G472), .ZN(n454) );
  INV_X1 U457 ( .A(KEYINPUT64), .ZN(n477) );
  BUF_X1 U458 ( .A(n743), .Z(n746) );
  AND2_X1 U459 ( .A1(n728), .A2(n365), .ZN(n473) );
  NAND2_X1 U460 ( .A1(n694), .A2(n480), .ZN(n474) );
  NOR2_X1 U461 ( .A1(n420), .A2(KEYINPUT103), .ZN(n415) );
  NAND2_X1 U462 ( .A1(G237), .A2(G234), .ZN(n524) );
  OR2_X1 U463 ( .A1(G902), .A2(G237), .ZN(n540) );
  XOR2_X1 U464 ( .A(G902), .B(KEYINPUT15), .Z(n539) );
  XNOR2_X1 U465 ( .A(G137), .B(G116), .ZN(n518) );
  XOR2_X1 U466 ( .A(G113), .B(KEYINPUT5), .Z(n520) );
  INV_X1 U467 ( .A(n689), .ZN(n400) );
  NAND2_X1 U468 ( .A1(n376), .A2(n375), .ZN(n374) );
  AND2_X1 U469 ( .A1(n635), .A2(n636), .ZN(n373) );
  OR2_X1 U470 ( .A1(n635), .A2(n636), .ZN(n377) );
  AND2_X1 U471 ( .A1(n774), .A2(n589), .ZN(n401) );
  XOR2_X1 U472 ( .A(G137), .B(G140), .Z(n502) );
  XNOR2_X1 U473 ( .A(n558), .B(n557), .ZN(n565) );
  XNOR2_X1 U474 ( .A(KEYINPUT99), .B(KEYINPUT12), .ZN(n561) );
  XOR2_X1 U475 ( .A(KEYINPUT66), .B(G131), .Z(n554) );
  XNOR2_X1 U476 ( .A(n439), .B(n438), .ZN(n499) );
  INV_X1 U477 ( .A(KEYINPUT96), .ZN(n438) );
  INV_X1 U478 ( .A(KEYINPUT16), .ZN(n466) );
  NOR2_X1 U479 ( .A1(n356), .A2(KEYINPUT72), .ZN(n649) );
  INV_X1 U480 ( .A(n574), .ZN(n576) );
  INV_X1 U481 ( .A(KEYINPUT101), .ZN(n469) );
  INV_X1 U482 ( .A(KEYINPUT33), .ZN(n523) );
  NOR2_X1 U483 ( .A1(n608), .A2(n440), .ZN(n632) );
  NOR2_X1 U484 ( .A1(n434), .A2(n408), .ZN(n407) );
  XNOR2_X1 U485 ( .A(n406), .B(n442), .ZN(n405) );
  BUF_X1 U486 ( .A(n614), .Z(n434) );
  BUF_X1 U487 ( .A(n707), .Z(n440) );
  INV_X1 U488 ( .A(KEYINPUT0), .ZN(n410) );
  XNOR2_X1 U489 ( .A(n432), .B(n494), .ZN(n659) );
  XNOR2_X1 U490 ( .A(n764), .B(n481), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n491), .B(n482), .ZN(n481) );
  XNOR2_X1 U492 ( .A(n437), .B(n552), .ZN(n745) );
  NAND2_X1 U493 ( .A1(n743), .A2(G475), .ZN(n461) );
  NOR2_X1 U494 ( .A1(n645), .A2(n633), .ZN(n403) );
  OR2_X1 U495 ( .A1(n380), .A2(n379), .ZN(n686) );
  NAND2_X1 U496 ( .A1(n383), .A2(n381), .ZN(n380) );
  NOR2_X1 U497 ( .A1(n382), .A2(n706), .ZN(n381) );
  INV_X1 U498 ( .A(KEYINPUT32), .ZN(n478) );
  NAND2_X1 U499 ( .A1(n409), .A2(n361), .ZN(n479) );
  XNOR2_X1 U500 ( .A(n452), .B(n368), .ZN(G57) );
  NAND2_X1 U501 ( .A1(n453), .A2(n459), .ZN(n452) );
  XNOR2_X1 U502 ( .A(n458), .B(n457), .ZN(G60) );
  INV_X1 U503 ( .A(KEYINPUT60), .ZN(n457) );
  NAND2_X1 U504 ( .A1(n460), .A2(n459), .ZN(n458) );
  XNOR2_X1 U505 ( .A(n461), .B(n358), .ZN(n460) );
  XNOR2_X1 U506 ( .A(n445), .B(n367), .ZN(n742) );
  NAND2_X1 U507 ( .A1(n746), .A2(G469), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n435), .B(n736), .ZN(n737) );
  XNOR2_X1 U509 ( .A(n472), .B(n471), .ZN(n730) );
  INV_X1 U510 ( .A(KEYINPUT119), .ZN(n471) );
  AND2_X1 U511 ( .A1(n377), .A2(n399), .ZN(n357) );
  XOR2_X1 U512 ( .A(n744), .B(n369), .Z(n358) );
  AND2_X1 U513 ( .A1(n372), .A2(n374), .ZN(n359) );
  XOR2_X1 U514 ( .A(KEYINPUT97), .B(G472), .Z(n360) );
  XOR2_X1 U515 ( .A(n583), .B(KEYINPUT105), .Z(n361) );
  XOR2_X1 U516 ( .A(n520), .B(n519), .Z(n362) );
  XOR2_X1 U517 ( .A(KEYINPUT86), .B(KEYINPUT39), .Z(n364) );
  OR2_X1 U518 ( .A1(n729), .A2(n695), .ZN(n365) );
  INV_X1 U519 ( .A(KEYINPUT103), .ZN(n419) );
  XOR2_X1 U520 ( .A(n656), .B(KEYINPUT62), .Z(n366) );
  XOR2_X1 U521 ( .A(n741), .B(n740), .Z(n367) );
  NOR2_X1 U522 ( .A1(n493), .A2(G952), .ZN(n750) );
  INV_X1 U523 ( .A(n750), .ZN(n459) );
  XOR2_X1 U524 ( .A(n657), .B(KEYINPUT92), .Z(n368) );
  XNOR2_X1 U525 ( .A(KEYINPUT59), .B(KEYINPUT91), .ZN(n369) );
  INV_X1 U526 ( .A(KEYINPUT88), .ZN(n395) );
  XNOR2_X1 U527 ( .A(n443), .B(n758), .ZN(n735) );
  INV_X2 U528 ( .A(KEYINPUT4), .ZN(n430) );
  NAND2_X1 U529 ( .A1(n743), .A2(G210), .ZN(n435) );
  AND2_X1 U530 ( .A1(n411), .A2(KEYINPUT34), .ZN(n424) );
  NOR2_X2 U531 ( .A1(n582), .A2(n639), .ZN(n663) );
  NAND2_X1 U532 ( .A1(n588), .A2(KEYINPUT44), .ZN(n397) );
  XNOR2_X1 U533 ( .A(n634), .B(KEYINPUT46), .ZN(n635) );
  NAND2_X1 U534 ( .A1(n407), .A2(n405), .ZN(n608) );
  XNOR2_X1 U535 ( .A(n565), .B(n564), .ZN(n566) );
  NAND2_X1 U536 ( .A1(n370), .A2(n414), .ZN(n418) );
  NAND2_X1 U537 ( .A1(n412), .A2(n413), .ZN(n370) );
  NOR2_X2 U538 ( .A1(n575), .A2(n574), .ZN(n683) );
  XNOR2_X1 U539 ( .A(n566), .B(n567), .ZN(n744) );
  NOR2_X1 U540 ( .A1(n701), .A2(n419), .ZN(n412) );
  INV_X1 U541 ( .A(n701), .ZN(n420) );
  XNOR2_X1 U542 ( .A(n371), .B(n522), .ZN(n656) );
  NAND2_X1 U543 ( .A1(n373), .A2(n378), .ZN(n372) );
  INV_X1 U544 ( .A(n636), .ZN(n375) );
  INV_X1 U545 ( .A(n378), .ZN(n376) );
  NOR2_X1 U546 ( .A1(n387), .A2(n385), .ZN(n379) );
  NAND2_X1 U547 ( .A1(n387), .A2(n384), .ZN(n383) );
  XNOR2_X2 U548 ( .A(n388), .B(n360), .ZN(n606) );
  NAND2_X1 U549 ( .A1(n389), .A2(n581), .ZN(n455) );
  AND2_X2 U550 ( .A1(n517), .A2(n639), .ZN(n389) );
  NAND2_X1 U551 ( .A1(n389), .A2(n606), .ZN(n717) );
  NAND2_X1 U552 ( .A1(n390), .A2(n395), .ZN(n394) );
  NAND2_X1 U553 ( .A1(n354), .A2(n391), .ZN(n390) );
  INV_X1 U554 ( .A(n663), .ZN(n391) );
  NAND2_X1 U555 ( .A1(n394), .A2(n392), .ZN(n398) );
  NOR2_X1 U556 ( .A1(n663), .A2(n395), .ZN(n393) );
  XNOR2_X1 U557 ( .A(n396), .B(KEYINPUT87), .ZN(n592) );
  NAND2_X1 U558 ( .A1(n398), .A2(n397), .ZN(n396) );
  NOR2_X1 U559 ( .A1(n400), .A2(n688), .ZN(n399) );
  NOR2_X1 U560 ( .A1(n584), .A2(n431), .ZN(n585) );
  NAND2_X1 U561 ( .A1(n590), .A2(n401), .ZN(n591) );
  NAND2_X1 U562 ( .A1(n695), .A2(n428), .ZN(n427) );
  OR2_X2 U563 ( .A1(n411), .A2(KEYINPUT34), .ZN(n426) );
  NAND2_X1 U564 ( .A1(n363), .A2(n425), .ZN(n429) );
  XNOR2_X2 U565 ( .A(n402), .B(n511), .ZN(n766) );
  XNOR2_X1 U566 ( .A(n402), .B(n551), .ZN(n437) );
  NAND2_X2 U567 ( .A1(n509), .A2(n510), .ZN(n402) );
  XNOR2_X1 U568 ( .A(n403), .B(KEYINPUT40), .ZN(n776) );
  NAND2_X1 U569 ( .A1(n632), .A2(n696), .ZN(n404) );
  NAND2_X1 U570 ( .A1(n606), .A2(n697), .ZN(n406) );
  NAND2_X1 U571 ( .A1(n617), .A2(n546), .ZN(n462) );
  XNOR2_X2 U572 ( .A(n605), .B(n545), .ZN(n617) );
  NAND2_X1 U573 ( .A1(n609), .A2(n697), .ZN(n605) );
  XNOR2_X1 U574 ( .A(n543), .B(n542), .ZN(n609) );
  NAND2_X1 U575 ( .A1(n409), .A2(n431), .ZN(n582) );
  AND2_X2 U576 ( .A1(n444), .A2(n411), .ZN(n571) );
  XNOR2_X2 U577 ( .A(n462), .B(n410), .ZN(n411) );
  NAND2_X1 U578 ( .A1(n411), .A2(n572), .ZN(n573) );
  NAND2_X1 U579 ( .A1(n578), .A2(n411), .ZN(n580) );
  OR2_X1 U580 ( .A1(n680), .A2(n666), .ZN(n413) );
  NAND2_X1 U581 ( .A1(n587), .A2(KEYINPUT44), .ZN(n421) );
  NAND2_X1 U582 ( .A1(n429), .A2(n569), .ZN(n422) );
  NAND2_X1 U583 ( .A1(n424), .A2(n423), .ZN(n425) );
  INV_X1 U584 ( .A(n695), .ZN(n423) );
  XNOR2_X2 U585 ( .A(n430), .B(G101), .ZN(n533) );
  NOR2_X2 U586 ( .A1(n573), .A2(n434), .ZN(n666) );
  XNOR2_X2 U587 ( .A(n433), .B(G146), .ZN(n535) );
  NOR2_X2 U588 ( .A1(n739), .A2(G902), .ZN(n516) );
  NAND2_X1 U589 ( .A1(n436), .A2(n503), .ZN(n506) );
  INV_X1 U590 ( .A(n504), .ZN(n436) );
  AND2_X2 U591 ( .A1(n648), .A2(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U592 ( .A1(n441), .A2(n506), .ZN(n513) );
  NAND2_X1 U593 ( .A1(n505), .A2(n504), .ZN(n441) );
  NOR2_X1 U594 ( .A1(n776), .A2(n777), .ZN(n634) );
  XNOR2_X1 U595 ( .A(n537), .B(n538), .ZN(n443) );
  INV_X1 U596 ( .A(n717), .ZN(n444) );
  INV_X1 U597 ( .A(KEYINPUT67), .ZN(n446) );
  XNOR2_X2 U598 ( .A(n455), .B(n523), .ZN(n695) );
  XNOR2_X2 U599 ( .A(n614), .B(n456), .ZN(n639) );
  XNOR2_X2 U600 ( .A(n501), .B(KEYINPUT93), .ZN(n530) );
  NAND2_X1 U601 ( .A1(n474), .A2(n473), .ZN(n472) );
  XNOR2_X2 U602 ( .A(n477), .B(G953), .ZN(n493) );
  INV_X1 U603 ( .A(n647), .ZN(n480) );
  NOR2_X2 U604 ( .A1(n737), .A2(n750), .ZN(n738) );
  NOR2_X2 U605 ( .A1(n660), .A2(n750), .ZN(n662) );
  XNOR2_X2 U606 ( .A(G110), .B(G104), .ZN(n501) );
  INV_X1 U607 ( .A(KEYINPUT47), .ZN(n621) );
  XNOR2_X1 U608 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n636) );
  INV_X1 U609 ( .A(n502), .ZN(n488) );
  INV_X1 U610 ( .A(n554), .ZN(n511) );
  XNOR2_X1 U611 ( .A(n521), .B(n362), .ZN(n522) );
  XNOR2_X1 U612 ( .A(n541), .B(KEYINPUT80), .ZN(n542) );
  INV_X1 U613 ( .A(KEYINPUT106), .ZN(n603) );
  INV_X1 U614 ( .A(KEYINPUT63), .ZN(n657) );
  INV_X1 U615 ( .A(KEYINPUT123), .ZN(n661) );
  XOR2_X1 U616 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n485) );
  INV_X1 U617 ( .A(n539), .ZN(n646) );
  NAND2_X1 U618 ( .A1(G234), .A2(n646), .ZN(n483) );
  XNOR2_X1 U619 ( .A(KEYINPUT20), .B(n483), .ZN(n497) );
  NAND2_X1 U620 ( .A1(n497), .A2(G217), .ZN(n484) );
  XNOR2_X1 U621 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U622 ( .A(KEYINPUT25), .B(n486), .ZN(n496) );
  XOR2_X1 U623 ( .A(KEYINPUT76), .B(KEYINPUT23), .Z(n490) );
  XNOR2_X1 U624 ( .A(G128), .B(KEYINPUT83), .ZN(n489) );
  XNOR2_X1 U625 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U626 ( .A1(G221), .A2(n547), .ZN(n494) );
  NOR2_X1 U627 ( .A1(n659), .A2(G902), .ZN(n495) );
  NAND2_X1 U628 ( .A1(n497), .A2(G221), .ZN(n498) );
  XNOR2_X1 U629 ( .A(n498), .B(KEYINPUT21), .ZN(n594) );
  INV_X1 U630 ( .A(n594), .ZN(n709) );
  INV_X1 U631 ( .A(n707), .ZN(n517) );
  NAND2_X1 U632 ( .A1(G227), .A2(n493), .ZN(n500) );
  INV_X1 U633 ( .A(n503), .ZN(n505) );
  NAND2_X1 U634 ( .A1(G134), .A2(n355), .ZN(n510) );
  NAND2_X1 U635 ( .A1(n508), .A2(n534), .ZN(n509) );
  XOR2_X1 U636 ( .A(n533), .B(G146), .Z(n512) );
  XNOR2_X1 U637 ( .A(G469), .B(KEYINPUT69), .ZN(n514) );
  XOR2_X1 U638 ( .A(n514), .B(KEYINPUT68), .Z(n515) );
  XNOR2_X2 U639 ( .A(n516), .B(n515), .ZN(n614) );
  XOR2_X1 U640 ( .A(G119), .B(KEYINPUT3), .Z(n529) );
  XOR2_X1 U641 ( .A(n518), .B(n529), .Z(n521) );
  NAND2_X1 U642 ( .A1(n556), .A2(G210), .ZN(n519) );
  NOR2_X1 U643 ( .A1(G898), .A2(n752), .ZN(n760) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(KEYINPUT94), .Z(n525) );
  XOR2_X1 U645 ( .A(n525), .B(n524), .Z(n527) );
  NAND2_X1 U646 ( .A1(n527), .A2(G902), .ZN(n526) );
  XNOR2_X1 U647 ( .A(n526), .B(KEYINPUT95), .ZN(n596) );
  NAND2_X1 U648 ( .A1(n760), .A2(n596), .ZN(n528) );
  AND2_X1 U649 ( .A1(n527), .A2(G952), .ZN(n726) );
  NAND2_X1 U650 ( .A1(n726), .A2(n752), .ZN(n595) );
  NAND2_X1 U651 ( .A1(n528), .A2(n595), .ZN(n546) );
  NAND2_X1 U652 ( .A1(G214), .A2(n540), .ZN(n697) );
  XOR2_X1 U653 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n532) );
  NAND2_X1 U654 ( .A1(G224), .A2(n493), .ZN(n531) );
  XNOR2_X1 U655 ( .A(n532), .B(n531), .ZN(n538) );
  XNOR2_X1 U656 ( .A(n535), .B(KEYINPUT78), .ZN(n536) );
  XNOR2_X1 U657 ( .A(n353), .B(n536), .ZN(n537) );
  NOR2_X1 U658 ( .A1(n735), .A2(n539), .ZN(n543) );
  NAND2_X1 U659 ( .A1(G210), .A2(n540), .ZN(n541) );
  XNOR2_X1 U660 ( .A(KEYINPUT65), .B(KEYINPUT73), .ZN(n544) );
  NAND2_X1 U661 ( .A1(n547), .A2(G217), .ZN(n552) );
  XNOR2_X1 U662 ( .A(n548), .B(G122), .ZN(n549) );
  XNOR2_X1 U663 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U664 ( .A(G104), .B(G143), .ZN(n555) );
  XNOR2_X1 U665 ( .A(n555), .B(n554), .ZN(n567) );
  NAND2_X1 U666 ( .A1(n556), .A2(G214), .ZN(n557) );
  XNOR2_X1 U667 ( .A(n559), .B(KEYINPUT98), .ZN(n563) );
  XNOR2_X1 U668 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U669 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U670 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n568) );
  OR2_X1 U671 ( .A1(n575), .A2(n576), .ZN(n610) );
  INV_X1 U672 ( .A(KEYINPUT31), .ZN(n570) );
  NOR2_X1 U673 ( .A1(n606), .A2(n440), .ZN(n572) );
  NAND2_X1 U674 ( .A1(n575), .A2(n574), .ZN(n633) );
  XOR2_X1 U675 ( .A(KEYINPUT102), .B(n683), .Z(n644) );
  AND2_X1 U676 ( .A1(n633), .A2(n644), .ZN(n701) );
  NAND2_X1 U677 ( .A1(n576), .A2(n575), .ZN(n699) );
  NOR2_X1 U678 ( .A1(n594), .A2(n699), .ZN(n577) );
  XNOR2_X1 U679 ( .A(KEYINPUT104), .B(n577), .ZN(n578) );
  INV_X1 U680 ( .A(n639), .ZN(n706) );
  NOR2_X1 U681 ( .A1(n431), .A2(n706), .ZN(n583) );
  NAND2_X1 U682 ( .A1(n585), .A2(n706), .ZN(n586) );
  INV_X1 U683 ( .A(n587), .ZN(n774) );
  XNOR2_X1 U684 ( .A(n588), .B(KEYINPUT89), .ZN(n590) );
  INV_X1 U685 ( .A(KEYINPUT44), .ZN(n589) );
  NAND2_X1 U686 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X2 U687 ( .A(n593), .B(KEYINPUT45), .ZN(n751) );
  NOR2_X1 U688 ( .A1(n710), .A2(n594), .ZN(n602) );
  INV_X1 U689 ( .A(n595), .ZN(n600) );
  INV_X1 U690 ( .A(n493), .ZN(n597) );
  NAND2_X1 U691 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U692 ( .A1(G900), .A2(n598), .ZN(n599) );
  NOR2_X1 U693 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U694 ( .A(KEYINPUT81), .B(n601), .ZN(n607) );
  NAND2_X1 U695 ( .A1(n602), .A2(n607), .ZN(n612) );
  INV_X1 U696 ( .A(n609), .ZN(n643) );
  NOR2_X1 U697 ( .A1(n643), .A2(n610), .ZN(n611) );
  NAND2_X1 U698 ( .A1(n632), .A2(n611), .ZN(n675) );
  NAND2_X1 U699 ( .A1(n686), .A2(n675), .ZN(n627) );
  NOR2_X1 U700 ( .A1(n701), .A2(KEYINPUT71), .ZN(n619) );
  NOR2_X1 U701 ( .A1(n712), .A2(n612), .ZN(n613) );
  XNOR2_X1 U702 ( .A(n613), .B(KEYINPUT28), .ZN(n616) );
  INV_X1 U703 ( .A(n434), .ZN(n615) );
  NAND2_X1 U704 ( .A1(n616), .A2(n615), .ZN(n630) );
  INV_X1 U705 ( .A(n617), .ZN(n618) );
  NAND2_X1 U706 ( .A1(n619), .A2(n677), .ZN(n620) );
  NAND2_X1 U707 ( .A1(n620), .A2(KEYINPUT47), .ZN(n625) );
  XOR2_X1 U708 ( .A(KEYINPUT71), .B(n701), .Z(n623) );
  NAND2_X1 U709 ( .A1(n677), .A2(n621), .ZN(n622) );
  OR2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U712 ( .A(KEYINPUT38), .B(n643), .ZN(n696) );
  NAND2_X1 U713 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U714 ( .A1(n699), .A2(n700), .ZN(n629) );
  XNOR2_X1 U715 ( .A(n629), .B(KEYINPUT41), .ZN(n729) );
  NOR2_X1 U716 ( .A1(n630), .A2(n729), .ZN(n631) );
  XNOR2_X1 U717 ( .A(n631), .B(KEYINPUT42), .ZN(n777) );
  XNOR2_X1 U718 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n637), .A2(n697), .ZN(n638) );
  NOR2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U721 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n689) );
  NOR2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n688) );
  AND2_X2 U724 ( .A1(n751), .A2(n356), .ZN(n648) );
  NOR2_X2 U725 ( .A1(n647), .A2(n646), .ZN(n655) );
  NAND2_X1 U726 ( .A1(n648), .A2(KEYINPUT72), .ZN(n653) );
  INV_X1 U727 ( .A(KEYINPUT2), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n649), .A2(n751), .ZN(n650) );
  AND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U731 ( .A1(G217), .A2(n743), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(n659), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(G66) );
  XOR2_X1 U734 ( .A(n663), .B(G101), .Z(G3) );
  XOR2_X1 U735 ( .A(G104), .B(KEYINPUT109), .Z(n665) );
  NAND2_X1 U736 ( .A1(n666), .A2(n681), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(G6) );
  XNOR2_X1 U738 ( .A(G107), .B(KEYINPUT110), .ZN(n670) );
  XOR2_X1 U739 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n668) );
  NAND2_X1 U740 ( .A1(n666), .A2(n683), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n670), .B(n669), .ZN(G9) );
  XOR2_X1 U743 ( .A(G110), .B(n671), .Z(G12) );
  XOR2_X1 U744 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n673) );
  NAND2_X1 U745 ( .A1(n677), .A2(n683), .ZN(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(n674) );
  XOR2_X1 U747 ( .A(G128), .B(n674), .Z(G30) );
  XNOR2_X1 U748 ( .A(G143), .B(KEYINPUT112), .ZN(n676) );
  XNOR2_X1 U749 ( .A(n676), .B(n675), .ZN(G45) );
  XOR2_X1 U750 ( .A(G146), .B(KEYINPUT113), .Z(n679) );
  NAND2_X1 U751 ( .A1(n677), .A2(n681), .ZN(n678) );
  XNOR2_X1 U752 ( .A(n679), .B(n678), .ZN(G48) );
  NAND2_X1 U753 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n682), .B(G113), .ZN(G15) );
  NAND2_X1 U755 ( .A1(n680), .A2(n683), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n684), .B(G116), .ZN(G18) );
  XOR2_X1 U757 ( .A(KEYINPUT114), .B(KEYINPUT37), .Z(n685) );
  XNOR2_X1 U758 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U759 ( .A(G125), .B(n687), .ZN(G27) );
  XOR2_X1 U760 ( .A(G134), .B(n688), .Z(G36) );
  XNOR2_X1 U761 ( .A(G140), .B(n689), .ZN(G42) );
  XNOR2_X1 U762 ( .A(KEYINPUT2), .B(KEYINPUT82), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n751), .A2(n691), .ZN(n690) );
  XNOR2_X1 U764 ( .A(n690), .B(KEYINPUT84), .ZN(n693) );
  NOR2_X1 U765 ( .A1(n691), .A2(n356), .ZN(n692) );
  NOR2_X1 U766 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U767 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U771 ( .A(KEYINPUT117), .B(n704), .Z(n705) );
  NOR2_X1 U772 ( .A1(n695), .A2(n705), .ZN(n723) );
  XNOR2_X1 U773 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n720) );
  NAND2_X1 U774 ( .A1(n440), .A2(n706), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n708), .B(KEYINPUT50), .ZN(n716) );
  NOR2_X1 U776 ( .A1(n431), .A2(n709), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n711), .B(KEYINPUT49), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U779 ( .A(KEYINPUT115), .B(n714), .ZN(n715) );
  NAND2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n718) );
  NAND2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U782 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U783 ( .A1(n729), .A2(n721), .ZN(n722) );
  NOR2_X1 U784 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U785 ( .A(KEYINPUT52), .B(n724), .Z(n725) );
  NAND2_X1 U786 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U787 ( .A(KEYINPUT118), .B(n727), .ZN(n728) );
  NOR2_X1 U788 ( .A1(G953), .A2(n730), .ZN(n731) );
  XNOR2_X1 U789 ( .A(KEYINPUT53), .B(n731), .ZN(G75) );
  XOR2_X1 U790 ( .A(KEYINPUT55), .B(KEYINPUT90), .Z(n733) );
  XNOR2_X1 U791 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n732) );
  XNOR2_X1 U792 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U793 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U794 ( .A(n738), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U795 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n741) );
  XNOR2_X1 U796 ( .A(n739), .B(KEYINPUT121), .ZN(n740) );
  NOR2_X1 U797 ( .A1(n750), .A2(n742), .ZN(G54) );
  XNOR2_X1 U798 ( .A(n745), .B(KEYINPUT122), .ZN(n748) );
  NAND2_X1 U799 ( .A1(G478), .A2(n746), .ZN(n747) );
  XNOR2_X1 U800 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U801 ( .A1(n750), .A2(n749), .ZN(G63) );
  NAND2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n756) );
  NAND2_X1 U803 ( .A1(G953), .A2(G224), .ZN(n753) );
  XNOR2_X1 U804 ( .A(KEYINPUT61), .B(n753), .ZN(n754) );
  NAND2_X1 U805 ( .A1(n754), .A2(G898), .ZN(n755) );
  NAND2_X1 U806 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U807 ( .A(n757), .B(KEYINPUT125), .ZN(n763) );
  XOR2_X1 U808 ( .A(n758), .B(G101), .Z(n759) );
  NOR2_X1 U809 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U810 ( .A(n761), .B(KEYINPUT124), .Z(n762) );
  XNOR2_X1 U811 ( .A(n763), .B(n762), .ZN(G69) );
  XOR2_X1 U812 ( .A(n764), .B(KEYINPUT4), .Z(n765) );
  XOR2_X1 U813 ( .A(n766), .B(n765), .Z(n770) );
  XOR2_X1 U814 ( .A(KEYINPUT126), .B(n770), .Z(n767) );
  XNOR2_X1 U815 ( .A(G227), .B(n767), .ZN(n768) );
  NAND2_X1 U816 ( .A1(n768), .A2(G900), .ZN(n769) );
  NAND2_X1 U817 ( .A1(n769), .A2(G953), .ZN(n773) );
  XNOR2_X1 U818 ( .A(n356), .B(n770), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n771), .A2(n493), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n773), .A2(n772), .ZN(G72) );
  XNOR2_X1 U821 ( .A(G122), .B(n774), .ZN(G24) );
  XOR2_X1 U822 ( .A(G119), .B(n775), .Z(G21) );
  XOR2_X1 U823 ( .A(G131), .B(n776), .Z(G33) );
  XOR2_X1 U824 ( .A(G137), .B(n777), .Z(G39) );
endmodule

