//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  XOR2_X1   g000(.A(G71gat), .B(G99gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT24), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n215), .A2(G169gat), .A3(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n215), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT65), .A3(new_n217), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n213), .A2(new_n219), .A3(new_n220), .A4(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT25), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT27), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT27), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n231), .A2(new_n232), .B1(G183gat), .B2(G190gat), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n230), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  INV_X1    g037(.A(new_n221), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n217), .B1(new_n239), .B2(KEYINPUT26), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n233), .B(new_n236), .C1(new_n238), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n243), .A2(new_n244), .B1(new_n207), .B2(new_n209), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n222), .A2(new_n246), .A3(new_n220), .A4(new_n217), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n225), .A2(new_n241), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(G113gat), .B2(G120gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(G113gat), .A2(G120gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(G127gat), .A2(G134gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(G127gat), .A2(G134gat), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n256), .A2(new_n257), .B1(KEYINPUT68), .B2(KEYINPUT1), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  INV_X1    g060(.A(G134gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G127gat), .A2(G134gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G113gat), .ZN(new_n266));
  INV_X1    g065(.A(G120gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(new_n251), .A3(new_n253), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n259), .A2(new_n270), .A3(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n250), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n248), .B1(new_n224), .B2(KEYINPUT25), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n277), .A2(new_n274), .A3(new_n273), .A4(new_n241), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n205), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n280), .A2(KEYINPUT33), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n204), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n278), .ZN(new_n283));
  INV_X1    g082(.A(new_n205), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n280), .B1(new_n204), .B2(KEYINPUT33), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT70), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n288));
  INV_X1    g087(.A(new_n286), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n279), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n282), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT34), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n276), .A2(new_n278), .A3(new_n292), .A4(new_n205), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n278), .A3(new_n205), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT34), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n285), .A2(KEYINPUT70), .A3(new_n286), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n288), .B1(new_n279), .B2(new_n289), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n297), .A2(new_n296), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n282), .A2(new_n302), .B1(new_n303), .B2(new_n294), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n306), .A2(KEYINPUT74), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(KEYINPUT74), .ZN(new_n308));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n307), .A2(new_n311), .A3(new_n308), .A4(new_n309), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G226gat), .ZN(new_n317));
  INV_X1    g116(.A(G233gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n277), .A2(new_n241), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n277), .A2(new_n241), .B1(new_n323), .B2(new_n320), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n316), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n323), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n250), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(new_n315), .A3(new_n321), .ZN(new_n328));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT75), .ZN(new_n330));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  NAND3_X1  g131(.A1(new_n325), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n325), .A2(new_n328), .A3(KEYINPUT30), .A4(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n328), .ZN(new_n337));
  INV_X1    g136(.A(new_n332), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT76), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n340));
  AOI211_X1 g139(.A(new_n340), .B(new_n332), .C1(new_n325), .C2(new_n328), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n335), .B(new_n336), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G228gat), .A2(G233gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  INV_X1    g145(.A(G155gat), .ZN(new_n347));
  INV_X1    g146(.A(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G141gat), .B(G148gat), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n346), .B(new_n349), .C1(new_n350), .C2(KEYINPUT2), .ZN(new_n351));
  INV_X1    g150(.A(G141gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G148gat), .ZN(new_n353));
  INV_X1    g152(.A(G148gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G141gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n349), .A2(new_n346), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n346), .A2(KEYINPUT2), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n351), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n313), .B2(new_n314), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(KEYINPUT3), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n351), .A2(new_n363), .A3(new_n359), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n323), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n316), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n362), .A2(new_n366), .A3(G22gat), .ZN(new_n367));
  AOI21_X1  g166(.A(G22gat), .B1(new_n362), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n345), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(new_n366), .ZN(new_n370));
  INV_X1    g169(.A(G22gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n362), .A2(G22gat), .A3(new_n366), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n344), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(KEYINPUT31), .ZN(new_n376));
  INV_X1    g175(.A(G50gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n369), .A2(new_n374), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n378), .B(new_n379), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n369), .B2(new_n374), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n360), .A2(new_n259), .A3(new_n270), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n271), .A2(new_n351), .A3(new_n359), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n385), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n351), .A2(new_n359), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n273), .A2(KEYINPUT4), .A3(new_n392), .A4(new_n274), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n259), .A2(new_n270), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n364), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  OAI22_X1  g196(.A1(new_n395), .A2(new_n360), .B1(new_n397), .B2(new_n390), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n391), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n273), .A2(new_n392), .A3(new_n274), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n397), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n392), .A2(new_n271), .A3(KEYINPUT4), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n390), .A2(KEYINPUT5), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n402), .A2(new_n396), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G57gat), .B(G85gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n405), .A3(new_n411), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n406), .A2(KEYINPUT83), .A3(new_n412), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n415), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n413), .A2(new_n417), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n305), .A2(new_n343), .A3(new_n384), .A4(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT35), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n406), .B2(new_n412), .ZN(new_n427));
  AOI211_X1 g226(.A(KEYINPUT78), .B(new_n411), .C1(new_n400), .C2(new_n405), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n418), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n421), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n418), .B(KEYINPUT79), .C1(new_n427), .C2(new_n428), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n342), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n302), .A2(new_n303), .A3(new_n294), .A4(new_n282), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n291), .A2(new_n298), .ZN(new_n435));
  AND4_X1   g234(.A1(KEYINPUT35), .A2(new_n384), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n424), .A2(new_n425), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT40), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n259), .A2(new_n270), .A3(KEYINPUT69), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT69), .B1(new_n259), .B2(new_n270), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT4), .B1(new_n441), .B2(new_n392), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n396), .A2(new_n403), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n390), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT82), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n446), .B(new_n390), .C1(new_n442), .C2(new_n443), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n388), .A2(new_n390), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n411), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT39), .B1(new_n445), .B2(new_n447), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n438), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n445), .A2(new_n447), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n449), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n456), .A2(KEYINPUT40), .A3(new_n411), .A4(new_n451), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n415), .A2(new_n419), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n454), .A2(new_n342), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n384), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n325), .A2(new_n328), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n315), .B1(new_n327), .B2(new_n321), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(KEYINPUT84), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n325), .A2(new_n328), .A3(new_n463), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(new_n338), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT85), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n467), .A2(new_n338), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n462), .A2(new_n465), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n468), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n467), .A2(new_n338), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n463), .B1(new_n325), .B2(new_n328), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT38), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n420), .A2(new_n478), .A3(new_n422), .A4(new_n333), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n384), .A2(KEYINPUT81), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT81), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n381), .B2(new_n383), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI22_X1  g283(.A1(new_n460), .A2(new_n480), .B1(new_n433), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n435), .A2(KEYINPUT36), .A3(new_n434), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n435), .B2(new_n434), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n488), .B2(KEYINPUT73), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT73), .ZN(new_n490));
  AOI211_X1 g289(.A(new_n490), .B(new_n487), .C1(new_n435), .C2(new_n434), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n437), .B1(new_n485), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT86), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT86), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n437), .B(new_n495), .C1(new_n485), .C2(new_n492), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT16), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(G1gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G1gat), .B2(new_n497), .ZN(new_n500));
  INV_X1    g299(.A(G8gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G29gat), .ZN(new_n504));
  INV_X1    g303(.A(G36gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT14), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT14), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n506), .B(new_n508), .C1(new_n504), .C2(new_n505), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n377), .A2(G43gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT87), .B(G50gat), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G43gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G43gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G50gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(new_n510), .A3(KEYINPUT15), .ZN(new_n517));
  MUX2_X1   g316(.A(new_n509), .B(new_n514), .S(new_n517), .Z(new_n518));
  AND2_X1   g317(.A1(new_n503), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(KEYINPUT17), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(new_n502), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n518), .B(new_n502), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n522), .B(KEYINPUT13), .Z(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT11), .ZN(new_n532));
  INV_X1    g331(.A(G169gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G197gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT12), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT18), .A3(new_n522), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n530), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n536), .B1(new_n530), .B2(new_n537), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n494), .A2(new_n496), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G64gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(G57gat), .ZN(new_n545));
  INV_X1    g344(.A(G57gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(G64gat), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(KEYINPUT88), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(KEYINPUT88), .B2(new_n547), .ZN(new_n549));
  NAND2_X1  g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  OR2_X1    g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT9), .B1(new_n547), .B2(new_n545), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n550), .A3(new_n551), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G127gat), .B(G155gat), .Z(new_n562));
  XOR2_X1   g361(.A(new_n562), .B(KEYINPUT20), .Z(new_n563));
  XNOR2_X1  g362(.A(new_n561), .B(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n503), .B1(KEYINPUT21), .B2(new_n558), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(new_n226), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n564), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G211gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n567), .B(new_n569), .Z(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT90), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  NOR2_X1   g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(KEYINPUT8), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G99gat), .B(G106gat), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n574), .A2(new_n582), .A3(new_n575), .A4(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n520), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  AND2_X1   g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n586), .A2(new_n518), .B1(KEYINPUT41), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n587), .A2(KEYINPUT41), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT91), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n591), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n570), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n557), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n558), .A2(new_n581), .A3(new_n583), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n586), .A2(KEYINPUT10), .A3(new_n558), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n602), .B1(new_n604), .B2(new_n606), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT92), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G176gat), .ZN(new_n614));
  INV_X1    g413(.A(G204gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n612), .B1(new_n611), .B2(new_n616), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n611), .A2(new_n616), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n601), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n543), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n431), .A2(new_n432), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n342), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT16), .B(G8gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(KEYINPUT42), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(G8gat), .B2(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(KEYINPUT42), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(G1325gat));
  OAI21_X1  g436(.A(KEYINPUT93), .B1(new_n489), .B2(new_n491), .ZN(new_n638));
  INV_X1    g437(.A(new_n487), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n299), .B2(new_n304), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n490), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n488), .A2(KEYINPUT73), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .A4(new_n486), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(G15gat), .B1(new_n625), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n305), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n648), .A2(G15gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n625), .B2(new_n649), .ZN(G1326gat));
  OR3_X1    g449(.A1(new_n625), .A2(KEYINPUT94), .A3(new_n484), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT94), .B1(new_n625), .B2(new_n484), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT43), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G22gat), .ZN(G1327gat));
  NOR3_X1   g454(.A1(new_n570), .A2(new_n600), .A3(new_n623), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n543), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n657), .A2(G29gat), .A3(new_n627), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT45), .ZN(new_n659));
  INV_X1    g458(.A(new_n600), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n494), .A2(new_n496), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT44), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n627), .A2(new_n343), .ZN(new_n663));
  INV_X1    g462(.A(new_n484), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n459), .B(new_n384), .C1(new_n479), .C2(new_n475), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n638), .A2(new_n644), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n437), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT44), .ZN(new_n669));
  AND4_X1   g468(.A1(KEYINPUT96), .A2(new_n668), .A3(new_n669), .A4(new_n660), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n600), .B1(new_n667), .B2(new_n437), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT96), .B1(new_n671), .B2(new_n669), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n662), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT95), .B1(new_n539), .B2(new_n540), .ZN(new_n674));
  INV_X1    g473(.A(new_n540), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT95), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n538), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(new_n570), .A3(new_n623), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n504), .B1(new_n680), .B2(new_n628), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n659), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT97), .ZN(G1328gat));
  NAND2_X1  g482(.A1(new_n673), .A2(new_n679), .ZN(new_n684));
  OAI21_X1  g483(.A(G36gat), .B1(new_n684), .B2(new_n343), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n657), .A2(G36gat), .A3(new_n343), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(KEYINPUT98), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT98), .B(KEYINPUT46), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n685), .B(new_n688), .C1(new_n686), .C2(new_n689), .ZN(G1329gat));
  NOR2_X1   g489(.A1(new_n684), .A2(new_n646), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT101), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n684), .B2(new_n646), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(G43gat), .A3(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n543), .A2(new_n515), .A3(new_n305), .A4(new_n656), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT99), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(KEYINPUT47), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n691), .B2(new_n515), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n699), .B2(new_n701), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n698), .B1(new_n702), .B2(new_n703), .ZN(G1330gat));
  INV_X1    g503(.A(new_n384), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n511), .B1(new_n680), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  INV_X1    g506(.A(new_n511), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n657), .A2(new_n484), .A3(new_n708), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n680), .A2(new_n664), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n711), .A2(KEYINPUT102), .A3(new_n708), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT102), .B1(new_n711), .B2(new_n708), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n712), .A2(new_n713), .A3(new_n709), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n710), .B1(new_n714), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g514(.A(new_n678), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(new_n601), .A3(new_n622), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n668), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n627), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(new_n546), .ZN(G1332gat));
  INV_X1    g519(.A(new_n718), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n343), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT103), .ZN(new_n724));
  NOR2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n718), .B2(new_n646), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n648), .A2(G71gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n718), .B2(new_n728), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g529(.A1(new_n721), .A2(new_n664), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g531(.A1(new_n716), .A2(new_n570), .A3(new_n622), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n673), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734), .B2(new_n627), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n716), .A2(new_n570), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n671), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n671), .A2(KEYINPUT51), .A3(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n623), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n627), .A2(G85gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n735), .B1(new_n742), .B2(new_n743), .ZN(G1336gat));
  OAI21_X1  g543(.A(G92gat), .B1(new_n734), .B2(new_n343), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n343), .A2(G92gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n742), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT52), .ZN(G1337gat));
  OR3_X1    g547(.A1(new_n742), .A2(G99gat), .A3(new_n648), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n673), .A2(new_n645), .A3(new_n733), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT104), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G99gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(KEYINPUT104), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(G1338gat));
  OAI21_X1  g553(.A(G106gat), .B1(new_n734), .B2(new_n384), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n384), .A2(G106gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n623), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n760));
  INV_X1    g559(.A(new_n758), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n673), .A2(new_n664), .A3(new_n733), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G106gat), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(KEYINPUT105), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n765), .A3(G106gat), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n760), .B(new_n756), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(KEYINPUT105), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n766), .A3(new_n758), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT106), .B1(new_n769), .B2(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n759), .B1(new_n767), .B2(new_n770), .ZN(G1339gat));
  NOR3_X1   g570(.A1(new_n716), .A2(new_n601), .A3(new_n623), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n528), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n526), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT107), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n521), .A2(new_n522), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n535), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n538), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n607), .A2(new_n608), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n602), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n607), .A2(new_n608), .A3(new_n603), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(KEYINPUT54), .A3(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n616), .B1(new_n609), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n618), .A2(new_n619), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n791), .A2(new_n597), .A3(new_n599), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n781), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n622), .A2(new_n779), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT109), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n622), .B2(new_n779), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n791), .A2(new_n792), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n796), .B(new_n798), .C1(new_n678), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n794), .B1(new_n800), .B2(new_n600), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n773), .B1(new_n801), .B2(new_n570), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n484), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n627), .A2(new_n342), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n305), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n805), .A2(new_n266), .A3(new_n541), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n802), .A2(new_n628), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n648), .A2(new_n705), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n807), .A2(new_n342), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n716), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n806), .A2(new_n811), .ZN(G1340gat));
  NOR3_X1   g611(.A1(new_n805), .A2(new_n267), .A3(new_n622), .ZN(new_n813));
  AOI21_X1  g612(.A(G120gat), .B1(new_n810), .B2(new_n623), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(G1341gat));
  INV_X1    g614(.A(new_n570), .ZN(new_n816));
  OAI21_X1  g615(.A(G127gat), .B1(new_n805), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n810), .A2(new_n261), .A3(new_n570), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1342gat));
  NAND3_X1  g618(.A1(new_n810), .A2(new_n262), .A3(new_n660), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n820), .A2(KEYINPUT56), .ZN(new_n822));
  OAI21_X1  g621(.A(G134gat), .B1(new_n805), .B2(new_n600), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(KEYINPUT110), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(KEYINPUT110), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n821), .B(new_n822), .C1(new_n824), .C2(new_n825), .ZN(G1343gat));
  NAND2_X1  g625(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n802), .A2(new_n828), .A3(new_n628), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n645), .A2(new_n342), .A3(new_n384), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n542), .A2(new_n352), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834));
  INV_X1    g633(.A(new_n794), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n788), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n785), .A2(new_n787), .A3(KEYINPUT111), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n789), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT55), .B1(new_n788), .B2(new_n836), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(KEYINPUT112), .A3(new_n838), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT113), .B1(new_n844), .B2(new_n791), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n790), .B1(new_n841), .B2(new_n843), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n541), .B1(new_n847), .B2(KEYINPUT113), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n795), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n835), .B1(new_n849), .B2(new_n660), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n772), .B1(new_n850), .B2(new_n816), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n484), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n834), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n795), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n842), .A2(KEYINPUT112), .A3(new_n838), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT112), .B1(new_n842), .B2(new_n838), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT113), .B(new_n791), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n542), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n860), .B2(new_n845), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n600), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n570), .B1(new_n862), .B2(new_n835), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT114), .B(new_n853), .C1(new_n863), .C2(new_n772), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n802), .A2(new_n705), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n852), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n855), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n646), .A2(new_n804), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n716), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n833), .B1(new_n870), .B2(G141gat), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n853), .B1(new_n863), .B2(new_n772), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n873), .A2(new_n834), .B1(new_n852), .B2(new_n865), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n868), .B1(new_n874), .B2(new_n864), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n352), .B1(new_n875), .B2(new_n542), .ZN(new_n876));
  XNOR2_X1  g675(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n831), .B2(new_n832), .ZN(new_n878));
  OAI22_X1  g677(.A1(new_n871), .A2(new_n872), .B1(new_n876), .B2(new_n878), .ZN(G1344gat));
  INV_X1    g678(.A(new_n831), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n354), .A3(new_n623), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G148gat), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n875), .B2(new_n623), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n624), .A2(new_n541), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n793), .A2(KEYINPUT118), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n781), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(KEYINPUT118), .B2(new_n793), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n862), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n885), .B1(new_n889), .B2(new_n570), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n484), .A2(KEYINPUT57), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n890), .A2(new_n891), .B1(KEYINPUT57), .B2(new_n865), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n868), .B(KEYINPUT117), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n623), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n882), .B1(new_n894), .B2(G148gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n881), .B1(new_n884), .B2(new_n895), .ZN(G1345gat));
  NAND2_X1  g695(.A1(new_n570), .A2(G155gat), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT119), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n867), .A2(new_n869), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n347), .B1(new_n831), .B2(new_n816), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n899), .A2(KEYINPUT120), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1346gat));
  NAND3_X1  g704(.A1(new_n880), .A2(new_n348), .A3(new_n660), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n875), .A2(new_n660), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n348), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n628), .A2(new_n343), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n305), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT121), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n803), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n533), .A3(new_n541), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n802), .A2(new_n627), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n809), .A2(new_n343), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n716), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n913), .B1(new_n533), .B2(new_n918), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n912), .B2(new_n622), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n622), .A2(G176gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n916), .B2(new_n921), .ZN(G1349gat));
  NAND4_X1  g721(.A1(new_n914), .A2(new_n235), .A3(new_n570), .A4(new_n915), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n802), .A2(new_n484), .A3(new_n570), .A4(new_n911), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G183gat), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n926), .A2(KEYINPUT122), .A3(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n923), .A2(new_n925), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(KEYINPUT60), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n932), .B1(new_n926), .B2(new_n927), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n930), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n928), .A2(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n917), .A2(new_n230), .A3(new_n660), .ZN(new_n936));
  OAI21_X1  g735(.A(G190gat), .B1(new_n912), .B2(new_n600), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1351gat));
  AND4_X1   g739(.A1(new_n342), .A2(new_n914), .A3(new_n705), .A4(new_n646), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n716), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n646), .A2(new_n909), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT124), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n892), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n542), .A2(G197gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n941), .A2(new_n615), .A3(new_n623), .ZN(new_n949));
  AND2_X1   g748(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n950));
  NOR2_X1   g749(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(G204gat), .B1(new_n945), .B2(new_n622), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n952), .B(new_n953), .C1(new_n950), .C2(new_n949), .ZN(G1353gat));
  INV_X1    g753(.A(G211gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n941), .A2(new_n955), .A3(new_n570), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n892), .A2(new_n570), .A3(new_n944), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  AOI21_X1  g759(.A(G218gat), .B1(new_n941), .B2(new_n660), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n660), .A2(G218gat), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT127), .Z(new_n963));
  AOI21_X1  g762(.A(new_n963), .B1(new_n946), .B2(KEYINPUT126), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n945), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n961), .B1(new_n964), .B2(new_n966), .ZN(G1355gat));
endmodule


