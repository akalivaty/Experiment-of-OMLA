//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n593, new_n596, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G137), .A3(new_n459), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G136), .ZN(new_n473));
  INV_X1    g048(.A(new_n470), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n459), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n459), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n473), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n469), .B2(new_n470), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n462), .A2(KEYINPUT70), .A3(new_n484), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(KEYINPUT4), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n459), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n469), .C2(new_n470), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n489), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  XNOR2_X1  g072(.A(KEYINPUT5), .B(G543), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT6), .B(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n504), .A2(new_n507), .ZN(G303));
  INV_X1    g083(.A(G303), .ZN(G166));
  XNOR2_X1  g084(.A(KEYINPUT71), .B(G89), .ZN(new_n510));
  INV_X1    g085(.A(G51), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n500), .A2(new_n510), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT7), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n498), .A2(G63), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(G168));
  NAND2_X1  g092(.A1(G77), .A2(G543), .ZN(new_n518));
  XOR2_X1   g093(.A(KEYINPUT5), .B(G543), .Z(new_n519));
  INV_X1    g094(.A(G64), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n506), .B1(new_n521), .B2(KEYINPUT72), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n522), .B1(KEYINPUT72), .B2(new_n521), .ZN(new_n523));
  INV_X1    g098(.A(new_n500), .ZN(new_n524));
  INV_X1    g099(.A(new_n502), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT73), .B(G52), .Z(new_n526));
  AOI22_X1  g101(.A1(G90), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n523), .A2(new_n527), .ZN(G301));
  INV_X1    g103(.A(G301), .ZN(G171));
  INV_X1    g104(.A(G81), .ZN(new_n530));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n500), .A2(new_n530), .B1(new_n502), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n498), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n506), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g112(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n538));
  NAND2_X1  g113(.A1(G1), .A2(G3), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND4_X1  g115(.A1(G319), .A2(G483), .A3(G661), .A4(new_n540), .ZN(G188));
  INV_X1    g116(.A(G53), .ZN(new_n542));
  OR3_X1    g117(.A1(new_n502), .A2(KEYINPUT9), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(KEYINPUT9), .B1(new_n502), .B2(new_n542), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(G78), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G65), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n519), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G651), .B1(new_n524), .B2(G91), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(G299));
  INV_X1    g125(.A(G168), .ZN(G286));
  OAI21_X1  g126(.A(G651), .B1(new_n498), .B2(G74), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n499), .A2(G49), .A3(G543), .ZN(new_n553));
  INV_X1    g128(.A(G87), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n552), .B(new_n553), .C1(new_n554), .C2(new_n500), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(KEYINPUT75), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(KEYINPUT75), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n557), .A2(new_n558), .ZN(G288));
  NAND2_X1  g134(.A1(G73), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G61), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n519), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(new_n525), .B2(G48), .ZN(new_n563));
  INV_X1    g138(.A(G86), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT76), .B1(new_n500), .B2(new_n564), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n500), .A2(KEYINPUT76), .A3(new_n564), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G305));
  INV_X1    g143(.A(G85), .ZN(new_n569));
  INV_X1    g144(.A(G47), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n500), .A2(new_n569), .B1(new_n502), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n506), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n571), .B2(new_n573), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G290));
  INV_X1    g152(.A(G868), .ZN(new_n578));
  OR3_X1    g153(.A1(G171), .A2(KEYINPUT78), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT78), .B1(G171), .B2(new_n578), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n498), .A2(new_n499), .A3(G92), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT10), .ZN(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n519), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n525), .B2(G54), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n579), .B(new_n580), .C1(G868), .C2(new_n588), .ZN(G284));
  OAI211_X1 g164(.A(new_n579), .B(new_n580), .C1(G868), .C2(new_n588), .ZN(G321));
  OR3_X1    g165(.A1(G168), .A2(KEYINPUT79), .A3(new_n578), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT79), .B1(G168), .B2(new_n578), .ZN(new_n592));
  INV_X1    g167(.A(G299), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(G868), .C2(new_n593), .ZN(G297));
  OAI211_X1 g169(.A(new_n591), .B(new_n592), .C1(G868), .C2(new_n593), .ZN(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n588), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n588), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n535), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g176(.A1(new_n472), .A2(G135), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT80), .Z(new_n603));
  NAND2_X1  g178(.A1(new_n476), .A2(G123), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT81), .ZN(new_n605));
  OR2_X1    g180(.A1(G99), .A2(G2105), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n606), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT82), .B(G2096), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n459), .A2(G2104), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n462), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2100), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n611), .A2(new_n612), .A3(new_n617), .ZN(G156));
  XOR2_X1   g193(.A(KEYINPUT15), .B(G2435), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2438), .ZN(new_n620));
  XOR2_X1   g195(.A(G2427), .B(G2430), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT84), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT83), .B(KEYINPUT14), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n620), .A2(new_n622), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n626), .B(new_n630), .Z(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(G14), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n632), .ZN(G401));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT85), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT17), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2084), .B(G2090), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n638), .B2(new_n640), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n639), .B2(new_n640), .ZN(new_n644));
  INV_X1    g219(.A(new_n640), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n645), .A2(new_n641), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT18), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n642), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1971), .B(G1976), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n653), .A2(new_n658), .A3(new_n656), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n653), .A2(new_n658), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n661));
  AOI211_X1 g236(.A(new_n657), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n660), .B2(new_n661), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G6), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n567), .B2(new_n671), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT32), .B(G1981), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n671), .A2(G22), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT89), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G303), .B2(G16), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G1971), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n671), .A2(G23), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n556), .B2(new_n671), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT33), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n675), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n685));
  AOI22_X1  g260(.A1(new_n472), .A2(G131), .B1(new_n476), .B2(G119), .ZN(new_n686));
  INV_X1    g261(.A(G95), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n687), .A2(new_n459), .A3(KEYINPUT87), .ZN(new_n688));
  AOI21_X1  g263(.A(KEYINPUT87), .B1(new_n687), .B2(new_n459), .ZN(new_n689));
  OAI221_X1 g264(.A(G2104), .B1(G107), .B2(new_n459), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(G25), .B(new_n693), .S(G29), .Z(new_n694));
  XOR2_X1   g269(.A(KEYINPUT35), .B(G1991), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n671), .A2(G24), .ZN(new_n698));
  INV_X1    g273(.A(G290), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n671), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1986), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n685), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n685), .A2(new_n702), .A3(KEYINPUT90), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(KEYINPUT36), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n707), .A2(new_n711), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n472), .A2(G141), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n476), .A2(G129), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n613), .A2(G105), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT98), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT26), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n723), .B2(G32), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT99), .Z(new_n728));
  INV_X1    g303(.A(G160), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G34), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n723), .B1(new_n730), .B2(G34), .ZN(new_n732));
  OAI22_X1  g307(.A1(new_n729), .A2(new_n723), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n728), .B1(G2084), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n723), .A2(G33), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT25), .Z(new_n738));
  INV_X1    g313(.A(new_n472), .ZN(new_n739));
  INV_X1    g314(.A(G139), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT95), .Z(new_n742));
  NAND2_X1  g317(.A1(G115), .A2(G2104), .ZN(new_n743));
  INV_X1    g318(.A(G127), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n471), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n459), .B1(new_n745), .B2(KEYINPUT96), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(KEYINPUT96), .B2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n736), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT97), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2072), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(G2072), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n735), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT100), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT31), .B(G11), .Z(new_n756));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n723), .B1(new_n757), .B2(G28), .ZN(new_n758));
  AOI21_X1  g333(.A(KEYINPUT101), .B1(new_n757), .B2(G28), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(KEYINPUT101), .A3(G28), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n756), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n608), .B2(new_n723), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n671), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n671), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1966), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n671), .A2(G5), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G171), .B2(new_n671), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT102), .Z(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT103), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n671), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT105), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1956), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT94), .B(G2067), .Z(new_n781));
  XOR2_X1   g356(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n723), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n476), .A2(G128), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT92), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n472), .A2(G140), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(G104), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n787), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n785), .B1(new_n793), .B2(G29), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n780), .B1(new_n781), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n770), .A2(G1961), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n796), .B(new_n797), .C1(new_n781), .C2(new_n795), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n773), .A2(new_n774), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n725), .A2(new_n726), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n734), .A2(G2084), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n588), .A2(new_n671), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G4), .B2(new_n671), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n671), .A2(G19), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n535), .B2(new_n671), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G1341), .Z(new_n808));
  NAND4_X1  g383(.A1(new_n800), .A2(new_n801), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n723), .A2(G35), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G162), .B2(new_n723), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT29), .B(G2090), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G164), .A2(new_n723), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G27), .B2(new_n723), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT104), .B(G2078), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n803), .B2(new_n804), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n809), .A2(new_n813), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  AND4_X1   g395(.A1(new_n775), .A2(new_n798), .A3(new_n799), .A4(new_n820), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n713), .A2(new_n755), .A3(new_n821), .ZN(G311));
  NAND3_X1  g397(.A1(new_n713), .A2(new_n755), .A3(new_n821), .ZN(G150));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n500), .A2(new_n824), .B1(new_n502), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n498), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(new_n506), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT106), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n535), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  INV_X1    g407(.A(new_n829), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n833), .A2(KEYINPUT106), .A3(new_n535), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n587), .A2(new_n596), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n829), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n721), .B(G164), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n793), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n748), .A2(KEYINPUT107), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n748), .A2(KEYINPUT107), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n476), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n459), .A2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G142), .B2(new_n472), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n615), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(new_n691), .Z(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n851), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n848), .A2(new_n858), .A3(new_n850), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n481), .B(new_n729), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n608), .ZN(new_n864));
  AOI21_X1  g439(.A(G37), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT108), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n861), .A2(new_n866), .ZN(new_n868));
  INV_X1    g443(.A(new_n864), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n860), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n865), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g447(.A1(new_n829), .A2(new_n578), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n699), .A2(G305), .ZN(new_n874));
  NAND2_X1  g449(.A1(G290), .A2(new_n567), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G303), .B(new_n555), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n877), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT110), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n835), .B(new_n598), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n587), .B(G299), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n889), .A2(KEYINPUT109), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(KEYINPUT109), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n888), .B1(new_n885), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n884), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n873), .B1(new_n894), .B2(new_n578), .ZN(G295));
  OAI21_X1  g470(.A(new_n873), .B1(new_n894), .B2(new_n578), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT111), .ZN(new_n897));
  XNOR2_X1  g472(.A(G301), .B(G286), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n835), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n832), .A2(new_n834), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n898), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n897), .B1(new_n903), .B2(new_n887), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n900), .B(new_n902), .C1(new_n890), .C2(new_n891), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n906), .B(new_n882), .C1(KEYINPUT111), .C2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n887), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n900), .A2(new_n889), .A3(new_n902), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n881), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n881), .B1(new_n908), .B2(new_n909), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT44), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n882), .B1(new_n905), .B2(KEYINPUT111), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n905), .B2(new_n904), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n921), .B2(new_n912), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT112), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT112), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n924), .B(KEYINPUT43), .C1(new_n921), .C2(new_n912), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n912), .A2(KEYINPUT43), .A3(new_n916), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n919), .B1(new_n927), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g503(.A(KEYINPUT127), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT114), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n793), .A2(G2067), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n793), .A2(G2067), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n933), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(KEYINPUT114), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n721), .A2(G1996), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n487), .A2(KEYINPUT4), .A3(new_n488), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n465), .A2(new_n466), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(G2105), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(G40), .A3(new_n463), .A4(new_n461), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  OR3_X1    g523(.A1(new_n944), .A2(G1996), .A3(new_n947), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT113), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n938), .A2(new_n948), .B1(new_n950), .B2(new_n722), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n691), .B(new_n696), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n948), .ZN(new_n954));
  XOR2_X1   g529(.A(G290), .B(G1986), .Z(new_n955));
  OAI211_X1 g530(.A(new_n951), .B(new_n953), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1981), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n563), .A2(new_n566), .A3(new_n957), .A4(new_n565), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n498), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n959));
  INV_X1    g534(.A(G48), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n959), .A2(new_n506), .B1(new_n960), .B2(new_n502), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n500), .A2(new_n564), .ZN(new_n962));
  OAI21_X1  g537(.A(G1981), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n958), .A2(KEYINPUT49), .A3(new_n963), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT118), .B(G8), .ZN(new_n968));
  INV_X1    g543(.A(new_n941), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n969), .B2(new_n489), .ZN(new_n970));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n464), .A2(new_n467), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n968), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n966), .A2(new_n967), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(G288), .A2(G1976), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n974), .A2(new_n975), .B1(new_n957), .B2(new_n567), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n973), .B(KEYINPUT119), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G8), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n947), .B1(new_n942), .B2(new_n943), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n943), .A2(G1384), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n940), .B2(new_n941), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT115), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n496), .A2(new_n984), .A3(new_n981), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n980), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1971), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n942), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n496), .A2(new_n939), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n947), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G2090), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n979), .B1(new_n988), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G303), .A2(G8), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n970), .A2(new_n972), .ZN(new_n1002));
  INV_X1    g577(.A(new_n968), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n556), .A2(G1976), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT52), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n557), .A2(new_n1007), .A3(new_n558), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n973), .A3(new_n1009), .A4(new_n1004), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n974), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n978), .B1(new_n1001), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n1015));
  INV_X1    g590(.A(G2078), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n980), .A2(new_n1016), .A3(new_n983), .A4(new_n985), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n496), .A2(new_n939), .A3(new_n992), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT50), .B1(new_n496), .B2(new_n939), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n972), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n772), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1018), .A2(G2078), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n980), .A2(new_n983), .A3(new_n985), .A4(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1019), .A2(G301), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1015), .B1(new_n1026), .B2(KEYINPUT124), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n947), .B1(new_n496), .B2(new_n981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(new_n944), .A3(new_n1024), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n1019), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G171), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1026), .A2(KEYINPUT124), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1027), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1025), .B1(G1961), .B2(new_n994), .ZN(new_n1036));
  OAI21_X1  g611(.A(G171), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1019), .A2(G301), .A3(new_n1023), .A4(new_n1029), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(KEYINPUT54), .A3(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT121), .B(G2084), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n972), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1042));
  INV_X1    g617(.A(G1966), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n982), .A2(new_n972), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT45), .B1(new_n496), .B2(new_n939), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n968), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(G168), .B2(new_n968), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1047), .B2(G286), .ZN(new_n1051));
  NOR2_X1   g626(.A1(G168), .A2(new_n968), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1028), .A2(new_n944), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n990), .A2(new_n993), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1056), .A2(new_n1043), .B1(new_n1057), .B2(new_n1041), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1055), .B1(new_n1058), .B2(new_n979), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1050), .B1(new_n1051), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1039), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1011), .B1(new_n997), .B2(new_n1000), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n942), .A2(new_n992), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n496), .A2(new_n989), .A3(new_n939), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(new_n995), .A3(new_n972), .A4(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n968), .B1(new_n988), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1063), .B1(new_n1067), .B2(new_n1000), .ZN(new_n1068));
  INV_X1    g643(.A(new_n985), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n984), .B1(new_n496), .B2(new_n981), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1971), .B1(new_n1071), .B2(new_n980), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1066), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1003), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1000), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(KEYINPUT120), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1062), .A2(new_n1068), .A3(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1034), .A2(new_n1061), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1064), .A2(new_n972), .A3(new_n1065), .ZN(new_n1079));
  INV_X1    g654(.A(G1956), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n980), .A2(new_n983), .A3(new_n985), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n1085));
  XNOR2_X1  g660(.A(G299), .B(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n994), .A2(G1348), .B1(G2067), .B2(new_n1002), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n588), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1081), .A2(new_n1083), .A3(new_n1086), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(G1341), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1002), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n986), .B2(G1996), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1097), .A2(KEYINPUT59), .A3(new_n535), .ZN(new_n1098));
  OAI221_X1 g673(.A(KEYINPUT60), .B1(G2067), .B2(new_n1002), .C1(new_n994), .C2(G1348), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(new_n588), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT59), .B1(new_n1097), .B2(new_n535), .ZN(new_n1101));
  OR3_X1    g676(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1092), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1086), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1088), .A2(KEYINPUT61), .A3(new_n1092), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1089), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(new_n588), .A3(new_n1099), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1093), .B1(new_n1102), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1014), .B1(new_n1078), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1060), .A2(new_n1114), .A3(KEYINPUT62), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1003), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1049), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(G1966), .B1(new_n1028), .B2(new_n944), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n972), .A2(new_n1040), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n990), .B2(new_n993), .ZN(new_n1122));
  OAI211_X1 g697(.A(G286), .B(new_n1003), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT51), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1054), .B1(new_n1116), .B2(G8), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1119), .B(KEYINPUT62), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT125), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1115), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(G301), .B1(new_n1030), .B2(new_n1019), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1062), .A2(new_n1068), .A3(new_n1076), .A4(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1060), .A2(KEYINPUT62), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1117), .A2(G286), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1062), .A2(new_n1068), .A3(new_n1076), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT63), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1117), .A2(new_n1135), .A3(G286), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1062), .B(new_n1137), .C1(new_n1000), .C2(new_n997), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1128), .A2(new_n1132), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n956), .B1(new_n1113), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n693), .A2(new_n696), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n933), .B1(new_n951), .B2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1142), .A2(new_n954), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n954), .A2(G1986), .A3(G290), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1144), .B(KEYINPUT48), .Z(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(new_n951), .A3(new_n953), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n949), .A2(KEYINPUT113), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n949), .A2(KEYINPUT113), .ZN(new_n1148));
  OR3_X1    g723(.A1(new_n1147), .A2(new_n1148), .A3(KEYINPUT46), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT47), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n934), .A2(new_n936), .A3(new_n722), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1153), .A2(new_n948), .B1(new_n950), .B2(KEYINPUT46), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1152), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1143), .B(new_n1146), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n929), .B1(new_n1140), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n956), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1026), .A2(KEYINPUT124), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1026), .A2(KEYINPUT124), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1160), .B(new_n1015), .C1(new_n1129), .C2(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1062), .A2(new_n1068), .A3(new_n1076), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1162), .A2(new_n1163), .A3(new_n1060), .A4(new_n1039), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1106), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1165), .A2(new_n1166), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1013), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1130), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1060), .A2(KEYINPUT62), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1169), .A2(new_n1170), .A3(new_n1115), .A4(new_n1127), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1159), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1146), .B1(new_n1142), .B2(new_n954), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT47), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1175), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1174), .A2(KEYINPUT127), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1158), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g756(.A(G319), .ZN(new_n1183));
  NOR3_X1   g757(.A1(G401), .A2(new_n1183), .A3(G227), .ZN(new_n1184));
  NAND4_X1  g758(.A1(new_n871), .A2(new_n918), .A3(new_n669), .A4(new_n1184), .ZN(G225));
  INV_X1    g759(.A(G225), .ZN(G308));
endmodule


