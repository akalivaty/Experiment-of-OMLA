

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U547 ( .A(n675), .B(n674), .ZN(n710) );
  INV_X1 U548 ( .A(n933), .ZN(n772) );
  AND2_X1 U549 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X2 U550 ( .A1(n710), .A2(n709), .ZN(n756) );
  INV_X1 U551 ( .A(KEYINPUT92), .ZN(n674) );
  XOR2_X1 U552 ( .A(KEYINPUT17), .B(n529), .Z(n854) );
  NOR2_X1 U553 ( .A1(G651), .A2(G543), .ZN(n632) );
  INV_X1 U554 ( .A(G651), .ZN(n518) );
  NOR2_X1 U555 ( .A1(G543), .A2(n518), .ZN(n512) );
  XNOR2_X1 U556 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n511) );
  XNOR2_X1 U557 ( .A(n512), .B(n511), .ZN(n631) );
  NAND2_X1 U558 ( .A1(G63), .A2(n631), .ZN(n515) );
  XOR2_X1 U559 ( .A(KEYINPUT0), .B(G543), .Z(n626) );
  NOR2_X1 U560 ( .A1(G651), .A2(n626), .ZN(n513) );
  XNOR2_X1 U561 ( .A(KEYINPUT64), .B(n513), .ZN(n629) );
  NAND2_X1 U562 ( .A1(G51), .A2(n629), .ZN(n514) );
  NAND2_X1 U563 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U564 ( .A(KEYINPUT6), .B(n516), .ZN(n523) );
  NAND2_X1 U565 ( .A1(n632), .A2(G89), .ZN(n517) );
  XNOR2_X1 U566 ( .A(n517), .B(KEYINPUT4), .ZN(n520) );
  NOR2_X1 U567 ( .A1(n626), .A2(n518), .ZN(n635) );
  NAND2_X1 U568 ( .A1(G76), .A2(n635), .ZN(n519) );
  NAND2_X1 U569 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U570 ( .A(n521), .B(KEYINPUT5), .Z(n522) );
  NOR2_X1 U571 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U572 ( .A(KEYINPUT78), .B(n524), .Z(n525) );
  XNOR2_X1 U573 ( .A(KEYINPUT7), .B(n525), .ZN(G168) );
  XOR2_X1 U574 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n857) );
  NAND2_X1 U576 ( .A1(n857), .A2(G113), .ZN(n528) );
  INV_X1 U577 ( .A(G2105), .ZN(n530) );
  AND2_X1 U578 ( .A1(n530), .A2(G2104), .ZN(n853) );
  NAND2_X1 U579 ( .A1(G101), .A2(n853), .ZN(n526) );
  XOR2_X1 U580 ( .A(KEYINPUT23), .B(n526), .Z(n527) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n534) );
  NOR2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  NAND2_X1 U583 ( .A1(G137), .A2(n854), .ZN(n532) );
  NOR2_X1 U584 ( .A1(G2104), .A2(n530), .ZN(n858) );
  NAND2_X1 U585 ( .A1(G125), .A2(n858), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U587 ( .A1(n534), .A2(n533), .ZN(G160) );
  NAND2_X1 U588 ( .A1(G85), .A2(n632), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G72), .A2(n635), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G60), .A2(n631), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G47), .A2(n629), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  OR2_X1 U594 ( .A1(n540), .A2(n539), .ZN(G290) );
  NAND2_X1 U595 ( .A1(G64), .A2(n631), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G52), .A2(n629), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n548) );
  NAND2_X1 U598 ( .A1(G90), .A2(n632), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G77), .A2(n635), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n545), .Z(n546) );
  XNOR2_X1 U602 ( .A(KEYINPUT66), .B(n546), .ZN(n547) );
  NOR2_X1 U603 ( .A1(n548), .A2(n547), .ZN(G171) );
  INV_X1 U604 ( .A(G132), .ZN(G219) );
  INV_X1 U605 ( .A(G57), .ZN(G237) );
  INV_X1 U606 ( .A(G120), .ZN(G236) );
  INV_X1 U607 ( .A(G108), .ZN(G238) );
  NAND2_X1 U608 ( .A1(G94), .A2(G452), .ZN(n549) );
  XNOR2_X1 U609 ( .A(n549), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U610 ( .A1(G7), .A2(G661), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n550), .B(KEYINPUT10), .ZN(n551) );
  XNOR2_X1 U612 ( .A(KEYINPUT70), .B(n551), .ZN(G223) );
  XOR2_X1 U613 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n553) );
  XNOR2_X1 U614 ( .A(KEYINPUT71), .B(G223), .ZN(n806) );
  NAND2_X1 U615 ( .A1(n806), .A2(G567), .ZN(n552) );
  XNOR2_X1 U616 ( .A(n553), .B(n552), .ZN(G234) );
  INV_X1 U617 ( .A(G860), .ZN(n588) );
  NAND2_X1 U618 ( .A1(G81), .A2(n632), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT12), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT74), .ZN(n557) );
  NAND2_X1 U621 ( .A1(G68), .A2(n635), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT13), .B(n558), .Z(n562) );
  NAND2_X1 U624 ( .A1(G56), .A2(n631), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT14), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT73), .ZN(n561) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G43), .A2(n629), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n924) );
  NOR2_X1 U630 ( .A1(n588), .A2(n924), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT75), .ZN(G153) );
  XOR2_X1 U632 ( .A(G171), .B(KEYINPUT76), .Z(G301) );
  NAND2_X1 U633 ( .A1(G868), .A2(G301), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G54), .A2(n629), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G92), .A2(n632), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G79), .A2(n635), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G66), .A2(n631), .ZN(n568) );
  XNOR2_X1 U639 ( .A(KEYINPUT77), .B(n568), .ZN(n569) );
  NOR2_X1 U640 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U642 ( .A(KEYINPUT15), .B(n573), .Z(n735) );
  INV_X1 U643 ( .A(G868), .ZN(n652) );
  NAND2_X1 U644 ( .A1(n735), .A2(n652), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(G284) );
  NAND2_X1 U646 ( .A1(G65), .A2(n631), .ZN(n577) );
  NAND2_X1 U647 ( .A1(G78), .A2(n635), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n632), .A2(G91), .ZN(n578) );
  XOR2_X1 U650 ( .A(KEYINPUT68), .B(n578), .Z(n579) );
  NOR2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G53), .A2(n629), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(G299) );
  XNOR2_X1 U654 ( .A(KEYINPUT79), .B(G868), .ZN(n583) );
  NOR2_X1 U655 ( .A1(G286), .A2(n583), .ZN(n586) );
  NOR2_X1 U656 ( .A1(G868), .A2(G299), .ZN(n584) );
  XNOR2_X1 U657 ( .A(n584), .B(KEYINPUT80), .ZN(n585) );
  NOR2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U659 ( .A(KEYINPUT81), .B(n587), .Z(G297) );
  NAND2_X1 U660 ( .A1(n588), .A2(G559), .ZN(n589) );
  INV_X1 U661 ( .A(n735), .ZN(n922) );
  NAND2_X1 U662 ( .A1(n589), .A2(n922), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U664 ( .A1(G868), .A2(n924), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n922), .A2(G868), .ZN(n591) );
  NOR2_X1 U666 ( .A1(G559), .A2(n591), .ZN(n592) );
  NOR2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U668 ( .A(KEYINPUT82), .B(n594), .ZN(G282) );
  NAND2_X1 U669 ( .A1(G123), .A2(n858), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n595), .B(KEYINPUT18), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n857), .A2(G111), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G99), .A2(n853), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G135), .A2(n854), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n973) );
  XNOR2_X1 U677 ( .A(n973), .B(G2096), .ZN(n603) );
  INV_X1 U678 ( .A(G2100), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(G156) );
  NAND2_X1 U680 ( .A1(G67), .A2(n631), .ZN(n605) );
  NAND2_X1 U681 ( .A1(G55), .A2(n629), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U683 ( .A(KEYINPUT84), .B(n606), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G93), .A2(n632), .ZN(n608) );
  NAND2_X1 U685 ( .A1(G80), .A2(n635), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n609) );
  OR2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n651) );
  NAND2_X1 U688 ( .A1(n922), .A2(G559), .ZN(n641) );
  XOR2_X1 U689 ( .A(KEYINPUT83), .B(n924), .Z(n611) );
  XNOR2_X1 U690 ( .A(n641), .B(n611), .ZN(n612) );
  NOR2_X1 U691 ( .A1(G860), .A2(n612), .ZN(n613) );
  XOR2_X1 U692 ( .A(n651), .B(n613), .Z(G145) );
  NAND2_X1 U693 ( .A1(G75), .A2(n635), .ZN(n614) );
  XOR2_X1 U694 ( .A(KEYINPUT88), .B(n614), .Z(n619) );
  NAND2_X1 U695 ( .A1(G62), .A2(n631), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G50), .A2(n629), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U698 ( .A(KEYINPUT87), .B(n617), .Z(n618) );
  NOR2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n632), .A2(G88), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(G303) );
  INV_X1 U702 ( .A(G303), .ZN(G166) );
  NAND2_X1 U703 ( .A1(G651), .A2(G74), .ZN(n623) );
  NAND2_X1 U704 ( .A1(G49), .A2(n629), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U706 ( .A1(n631), .A2(n624), .ZN(n625) );
  XOR2_X1 U707 ( .A(KEYINPUT85), .B(n625), .Z(n628) );
  NAND2_X1 U708 ( .A1(n626), .A2(G87), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(G288) );
  NAND2_X1 U710 ( .A1(n629), .A2(G48), .ZN(n630) );
  XNOR2_X1 U711 ( .A(n630), .B(KEYINPUT86), .ZN(n640) );
  NAND2_X1 U712 ( .A1(G61), .A2(n631), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G86), .A2(n632), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n635), .A2(G73), .ZN(n636) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(G305) );
  XOR2_X1 U719 ( .A(KEYINPUT90), .B(n641), .Z(n649) );
  XNOR2_X1 U720 ( .A(G166), .B(G288), .ZN(n646) );
  XOR2_X1 U721 ( .A(KEYINPUT89), .B(KEYINPUT19), .Z(n642) );
  XNOR2_X1 U722 ( .A(G290), .B(n642), .ZN(n643) );
  XOR2_X1 U723 ( .A(n651), .B(n643), .Z(n644) );
  XNOR2_X1 U724 ( .A(n644), .B(n924), .ZN(n645) );
  XNOR2_X1 U725 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U726 ( .A(n647), .B(G299), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(G305), .ZN(n876) );
  XNOR2_X1 U728 ( .A(n649), .B(n876), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n650), .A2(G868), .ZN(n654) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n654), .A2(n653), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2078), .A2(G2084), .ZN(n655) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n658), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U738 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NOR2_X1 U739 ( .A1(G238), .A2(G236), .ZN(n659) );
  NAND2_X1 U740 ( .A1(G69), .A2(n659), .ZN(n660) );
  NOR2_X1 U741 ( .A1(n660), .A2(G237), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n661), .B(KEYINPUT91), .ZN(n811) );
  NAND2_X1 U743 ( .A1(G567), .A2(n811), .ZN(n666) );
  NOR2_X1 U744 ( .A1(G219), .A2(G220), .ZN(n662) );
  XOR2_X1 U745 ( .A(KEYINPUT22), .B(n662), .Z(n663) );
  NOR2_X1 U746 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U747 ( .A1(G96), .A2(n664), .ZN(n812) );
  NAND2_X1 U748 ( .A1(G2106), .A2(n812), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n666), .A2(n665), .ZN(n813) );
  NAND2_X1 U750 ( .A1(G483), .A2(G661), .ZN(n667) );
  NOR2_X1 U751 ( .A1(n813), .A2(n667), .ZN(n810) );
  NAND2_X1 U752 ( .A1(n810), .A2(G36), .ZN(G176) );
  NAND2_X1 U753 ( .A1(G102), .A2(n853), .ZN(n669) );
  NAND2_X1 U754 ( .A1(G138), .A2(n854), .ZN(n668) );
  NAND2_X1 U755 ( .A1(n669), .A2(n668), .ZN(n673) );
  NAND2_X1 U756 ( .A1(G114), .A2(n857), .ZN(n671) );
  NAND2_X1 U757 ( .A1(G126), .A2(n858), .ZN(n670) );
  NAND2_X1 U758 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U759 ( .A1(n673), .A2(n672), .ZN(G164) );
  XNOR2_X1 U760 ( .A(G1986), .B(G290), .ZN(n936) );
  NAND2_X1 U761 ( .A1(G40), .A2(G160), .ZN(n675) );
  INV_X1 U762 ( .A(n710), .ZN(n676) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n676), .A2(n709), .ZN(n801) );
  NAND2_X1 U765 ( .A1(n936), .A2(n801), .ZN(n791) );
  XOR2_X1 U766 ( .A(G2067), .B(KEYINPUT37), .Z(n677) );
  XNOR2_X1 U767 ( .A(KEYINPUT93), .B(n677), .ZN(n799) );
  XNOR2_X1 U768 ( .A(KEYINPUT94), .B(KEYINPUT34), .ZN(n681) );
  NAND2_X1 U769 ( .A1(G104), .A2(n853), .ZN(n679) );
  NAND2_X1 U770 ( .A1(G140), .A2(n854), .ZN(n678) );
  NAND2_X1 U771 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U772 ( .A(n681), .B(n680), .ZN(n688) );
  NAND2_X1 U773 ( .A1(n858), .A2(G128), .ZN(n682) );
  XNOR2_X1 U774 ( .A(KEYINPUT95), .B(n682), .ZN(n685) );
  NAND2_X1 U775 ( .A1(n857), .A2(G116), .ZN(n683) );
  XOR2_X1 U776 ( .A(KEYINPUT96), .B(n683), .Z(n684) );
  NOR2_X1 U777 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U778 ( .A(n686), .B(KEYINPUT35), .ZN(n687) );
  NOR2_X1 U779 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U780 ( .A(KEYINPUT36), .B(n689), .ZN(n872) );
  NOR2_X1 U781 ( .A1(n799), .A2(n872), .ZN(n971) );
  NAND2_X1 U782 ( .A1(n801), .A2(n971), .ZN(n797) );
  NAND2_X1 U783 ( .A1(G107), .A2(n857), .ZN(n691) );
  NAND2_X1 U784 ( .A1(G119), .A2(n858), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U786 ( .A1(G131), .A2(n854), .ZN(n692) );
  XNOR2_X1 U787 ( .A(KEYINPUT97), .B(n692), .ZN(n693) );
  NOR2_X1 U788 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n853), .A2(G95), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n867) );
  NAND2_X1 U791 ( .A1(G1991), .A2(n867), .ZN(n705) );
  NAND2_X1 U792 ( .A1(G117), .A2(n857), .ZN(n698) );
  NAND2_X1 U793 ( .A1(G141), .A2(n854), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n853), .A2(G105), .ZN(n699) );
  XOR2_X1 U796 ( .A(KEYINPUT38), .B(n699), .Z(n700) );
  NOR2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n858), .A2(G129), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n703), .A2(n702), .ZN(n849) );
  NAND2_X1 U800 ( .A1(G1996), .A2(n849), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U802 ( .A(KEYINPUT98), .B(n706), .Z(n974) );
  XNOR2_X1 U803 ( .A(KEYINPUT99), .B(n801), .ZN(n707) );
  NOR2_X1 U804 ( .A1(n974), .A2(n707), .ZN(n794) );
  INV_X1 U805 ( .A(n794), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n797), .A2(n708), .ZN(n789) );
  NAND2_X1 U807 ( .A1(G8), .A2(n756), .ZN(n782) );
  NOR2_X1 U808 ( .A1(G1981), .A2(G305), .ZN(n711) );
  XOR2_X1 U809 ( .A(n711), .B(KEYINPUT24), .Z(n712) );
  NOR2_X1 U810 ( .A1(n782), .A2(n712), .ZN(n787) );
  NOR2_X1 U811 ( .A1(G1976), .A2(G288), .ZN(n715) );
  NAND2_X1 U812 ( .A1(n715), .A2(KEYINPUT33), .ZN(n713) );
  NOR2_X1 U813 ( .A1(n782), .A2(n713), .ZN(n777) );
  NOR2_X1 U814 ( .A1(G1971), .A2(G303), .ZN(n714) );
  NOR2_X1 U815 ( .A1(n715), .A2(n714), .ZN(n941) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n782), .ZN(n767) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n756), .ZN(n764) );
  NOR2_X1 U818 ( .A1(n767), .A2(n764), .ZN(n716) );
  XNOR2_X1 U819 ( .A(n716), .B(KEYINPUT104), .ZN(n717) );
  NAND2_X1 U820 ( .A1(n717), .A2(G8), .ZN(n718) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n718), .ZN(n719) );
  NOR2_X1 U822 ( .A1(G168), .A2(n719), .ZN(n724) );
  XOR2_X1 U823 ( .A(KEYINPUT25), .B(G2078), .Z(n951) );
  NOR2_X1 U824 ( .A1(n951), .A2(n756), .ZN(n720) );
  XOR2_X1 U825 ( .A(KEYINPUT100), .B(n720), .Z(n722) );
  INV_X1 U826 ( .A(G1961), .ZN(n898) );
  NAND2_X1 U827 ( .A1(n756), .A2(n898), .ZN(n721) );
  NAND2_X1 U828 ( .A1(n722), .A2(n721), .ZN(n751) );
  NOR2_X1 U829 ( .A1(G171), .A2(n751), .ZN(n723) );
  NOR2_X1 U830 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U831 ( .A(KEYINPUT31), .B(n725), .Z(n755) );
  NAND2_X1 U832 ( .A1(G1348), .A2(n756), .ZN(n727) );
  INV_X1 U833 ( .A(n756), .ZN(n738) );
  NAND2_X1 U834 ( .A1(n738), .A2(G2067), .ZN(n726) );
  NAND2_X1 U835 ( .A1(n727), .A2(n726), .ZN(n734) );
  NOR2_X1 U836 ( .A1(n735), .A2(n734), .ZN(n733) );
  XNOR2_X1 U837 ( .A(KEYINPUT102), .B(G1996), .ZN(n948) );
  NAND2_X1 U838 ( .A1(n948), .A2(n738), .ZN(n728) );
  XNOR2_X1 U839 ( .A(n728), .B(KEYINPUT26), .ZN(n730) );
  NAND2_X1 U840 ( .A1(n756), .A2(G1341), .ZN(n729) );
  NAND2_X1 U841 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U842 ( .A1(n731), .A2(n924), .ZN(n732) );
  NOR2_X1 U843 ( .A1(n733), .A2(n732), .ZN(n737) );
  AND2_X1 U844 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U845 ( .A1(n737), .A2(n736), .ZN(n745) );
  NAND2_X1 U846 ( .A1(n738), .A2(G2072), .ZN(n739) );
  XOR2_X1 U847 ( .A(KEYINPUT27), .B(n739), .Z(n742) );
  NAND2_X1 U848 ( .A1(G1956), .A2(n756), .ZN(n740) );
  XOR2_X1 U849 ( .A(KEYINPUT101), .B(n740), .Z(n741) );
  NAND2_X1 U850 ( .A1(n742), .A2(n741), .ZN(n746) );
  NOR2_X1 U851 ( .A1(G299), .A2(n746), .ZN(n743) );
  XOR2_X1 U852 ( .A(KEYINPUT103), .B(n743), .Z(n744) );
  NOR2_X1 U853 ( .A1(n745), .A2(n744), .ZN(n749) );
  NAND2_X1 U854 ( .A1(G299), .A2(n746), .ZN(n747) );
  XOR2_X1 U855 ( .A(KEYINPUT28), .B(n747), .Z(n748) );
  NOR2_X1 U856 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U857 ( .A(n750), .B(KEYINPUT29), .ZN(n753) );
  NAND2_X1 U858 ( .A1(G171), .A2(n751), .ZN(n752) );
  NAND2_X1 U859 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U860 ( .A1(n755), .A2(n754), .ZN(n765) );
  NAND2_X1 U861 ( .A1(n765), .A2(G286), .ZN(n761) );
  NOR2_X1 U862 ( .A1(G1971), .A2(n782), .ZN(n758) );
  NOR2_X1 U863 ( .A1(G2090), .A2(n756), .ZN(n757) );
  NOR2_X1 U864 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U865 ( .A1(n759), .A2(G303), .ZN(n760) );
  NAND2_X1 U866 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U867 ( .A1(G8), .A2(n762), .ZN(n763) );
  XNOR2_X1 U868 ( .A(n763), .B(KEYINPUT32), .ZN(n771) );
  NAND2_X1 U869 ( .A1(G8), .A2(n764), .ZN(n769) );
  INV_X1 U870 ( .A(n765), .ZN(n766) );
  NOR2_X1 U871 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U872 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U873 ( .A1(n771), .A2(n770), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n941), .A2(n781), .ZN(n774) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n933) );
  NOR2_X1 U876 ( .A1(n782), .A2(n772), .ZN(n773) );
  NOR2_X1 U877 ( .A1(KEYINPUT33), .A2(n775), .ZN(n776) );
  NOR2_X1 U878 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U879 ( .A(G1981), .B(G305), .Z(n928) );
  NAND2_X1 U880 ( .A1(n778), .A2(n928), .ZN(n785) );
  NOR2_X1 U881 ( .A1(G2090), .A2(G303), .ZN(n779) );
  NAND2_X1 U882 ( .A1(G8), .A2(n779), .ZN(n780) );
  NAND2_X1 U883 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U884 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U885 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U886 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U887 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n804) );
  NOR2_X1 U889 ( .A1(G1996), .A2(n849), .ZN(n980) );
  NOR2_X1 U890 ( .A1(G1986), .A2(G290), .ZN(n792) );
  NOR2_X1 U891 ( .A1(G1991), .A2(n867), .ZN(n977) );
  NOR2_X1 U892 ( .A1(n792), .A2(n977), .ZN(n793) );
  NOR2_X1 U893 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U894 ( .A1(n980), .A2(n795), .ZN(n796) );
  XNOR2_X1 U895 ( .A(n796), .B(KEYINPUT39), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U897 ( .A1(n799), .A2(n872), .ZN(n969) );
  NAND2_X1 U898 ( .A1(n800), .A2(n969), .ZN(n802) );
  NAND2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U901 ( .A(KEYINPUT40), .B(n805), .ZN(G329) );
  NAND2_X1 U902 ( .A1(G2106), .A2(n806), .ZN(G217) );
  AND2_X1 U903 ( .A1(G15), .A2(G2), .ZN(n807) );
  NAND2_X1 U904 ( .A1(G661), .A2(n807), .ZN(G259) );
  NAND2_X1 U905 ( .A1(G3), .A2(G1), .ZN(n808) );
  XOR2_X1 U906 ( .A(KEYINPUT107), .B(n808), .Z(n809) );
  NAND2_X1 U907 ( .A1(n810), .A2(n809), .ZN(G188) );
  XOR2_X1 U908 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  NOR2_X1 U909 ( .A1(n812), .A2(n811), .ZN(G325) );
  XNOR2_X1 U910 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U912 ( .A(G96), .ZN(G221) );
  XOR2_X1 U913 ( .A(KEYINPUT110), .B(n813), .Z(G319) );
  XOR2_X1 U914 ( .A(KEYINPUT111), .B(G2678), .Z(n815) );
  XNOR2_X1 U915 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n814) );
  XNOR2_X1 U916 ( .A(n815), .B(n814), .ZN(n819) );
  XOR2_X1 U917 ( .A(KEYINPUT112), .B(G2090), .Z(n817) );
  XNOR2_X1 U918 ( .A(G2067), .B(G2072), .ZN(n816) );
  XNOR2_X1 U919 ( .A(n817), .B(n816), .ZN(n818) );
  XOR2_X1 U920 ( .A(n819), .B(n818), .Z(n821) );
  XNOR2_X1 U921 ( .A(G2096), .B(G2100), .ZN(n820) );
  XNOR2_X1 U922 ( .A(n821), .B(n820), .ZN(n823) );
  XOR2_X1 U923 ( .A(G2078), .B(G2084), .Z(n822) );
  XNOR2_X1 U924 ( .A(n823), .B(n822), .ZN(G227) );
  XOR2_X1 U925 ( .A(G1991), .B(G1986), .Z(n825) );
  XNOR2_X1 U926 ( .A(G1961), .B(G1956), .ZN(n824) );
  XNOR2_X1 U927 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U928 ( .A(G1976), .B(G1981), .Z(n827) );
  XNOR2_X1 U929 ( .A(G1966), .B(G1971), .ZN(n826) );
  XNOR2_X1 U930 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U931 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U932 ( .A(G2474), .B(KEYINPUT41), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n833) );
  XOR2_X1 U934 ( .A(G1996), .B(KEYINPUT113), .Z(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(G229) );
  NAND2_X1 U936 ( .A1(n853), .A2(G100), .ZN(n840) );
  NAND2_X1 U937 ( .A1(G112), .A2(n857), .ZN(n835) );
  NAND2_X1 U938 ( .A1(G136), .A2(n854), .ZN(n834) );
  NAND2_X1 U939 ( .A1(n835), .A2(n834), .ZN(n838) );
  NAND2_X1 U940 ( .A1(n858), .A2(G124), .ZN(n836) );
  XOR2_X1 U941 ( .A(KEYINPUT44), .B(n836), .Z(n837) );
  NOR2_X1 U942 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U943 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U944 ( .A(KEYINPUT114), .B(n841), .Z(G162) );
  NAND2_X1 U945 ( .A1(G118), .A2(n857), .ZN(n843) );
  NAND2_X1 U946 ( .A1(G130), .A2(n858), .ZN(n842) );
  NAND2_X1 U947 ( .A1(n843), .A2(n842), .ZN(n848) );
  NAND2_X1 U948 ( .A1(G106), .A2(n853), .ZN(n845) );
  NAND2_X1 U949 ( .A1(G142), .A2(n854), .ZN(n844) );
  NAND2_X1 U950 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U951 ( .A(KEYINPUT45), .B(n846), .Z(n847) );
  NOR2_X1 U952 ( .A1(n848), .A2(n847), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n973), .B(n849), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n850), .B(G162), .ZN(n851) );
  XOR2_X1 U955 ( .A(n852), .B(n851), .Z(n865) );
  NAND2_X1 U956 ( .A1(G103), .A2(n853), .ZN(n856) );
  NAND2_X1 U957 ( .A1(G139), .A2(n854), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G115), .A2(n857), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G127), .A2(n858), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(KEYINPUT47), .B(n861), .Z(n862) );
  NOR2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n984) );
  XNOR2_X1 U964 ( .A(G160), .B(n984), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n874) );
  XOR2_X1 U966 ( .A(KEYINPUT116), .B(KEYINPUT115), .Z(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(n868), .B(KEYINPUT48), .Z(n870) );
  XNOR2_X1 U969 ( .A(G164), .B(KEYINPUT46), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n875) );
  NOR2_X1 U973 ( .A1(G37), .A2(n875), .ZN(G395) );
  XNOR2_X1 U974 ( .A(G286), .B(n876), .ZN(n878) );
  XNOR2_X1 U975 ( .A(G171), .B(n922), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n879) );
  NOR2_X1 U977 ( .A1(G37), .A2(n879), .ZN(G397) );
  XNOR2_X1 U978 ( .A(G2435), .B(G2443), .ZN(n889) );
  XOR2_X1 U979 ( .A(G2454), .B(G2430), .Z(n881) );
  XNOR2_X1 U980 ( .A(G2446), .B(KEYINPUT105), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n885) );
  XOR2_X1 U982 ( .A(G2451), .B(G2427), .Z(n883) );
  XNOR2_X1 U983 ( .A(G1341), .B(G1348), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U985 ( .A(n885), .B(n884), .Z(n887) );
  XNOR2_X1 U986 ( .A(KEYINPUT106), .B(G2438), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n890) );
  NAND2_X1 U989 ( .A1(n890), .A2(G14), .ZN(n897) );
  NAND2_X1 U990 ( .A1(n897), .A2(G319), .ZN(n894) );
  NOR2_X1 U991 ( .A1(G227), .A2(G229), .ZN(n891) );
  XOR2_X1 U992 ( .A(KEYINPUT117), .B(n891), .Z(n892) );
  XNOR2_X1 U993 ( .A(n892), .B(KEYINPUT49), .ZN(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n896) );
  NOR2_X1 U995 ( .A1(G395), .A2(G397), .ZN(n895) );
  NAND2_X1 U996 ( .A1(n896), .A2(n895), .ZN(G225) );
  INV_X1 U997 ( .A(G225), .ZN(G308) );
  INV_X1 U998 ( .A(n897), .ZN(G401) );
  XNOR2_X1 U999 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1002) );
  XNOR2_X1 U1000 ( .A(n898), .B(G5), .ZN(n918) );
  XOR2_X1 U1001 ( .A(G1966), .B(G21), .Z(n909) );
  XNOR2_X1 U1002 ( .A(G1348), .B(KEYINPUT59), .ZN(n899) );
  XNOR2_X1 U1003 ( .A(n899), .B(G4), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(G1956), .B(G20), .ZN(n901) );
  XNOR2_X1 U1005 ( .A(G6), .B(G1981), .ZN(n900) );
  NOR2_X1 U1006 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U1007 ( .A1(n903), .A2(n902), .ZN(n906) );
  XNOR2_X1 U1008 ( .A(KEYINPUT124), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1009 ( .A(G19), .B(n904), .ZN(n905) );
  NOR2_X1 U1010 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1011 ( .A(KEYINPUT60), .B(n907), .ZN(n908) );
  NAND2_X1 U1012 ( .A1(n909), .A2(n908), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(G1971), .B(G22), .ZN(n911) );
  XNOR2_X1 U1014 ( .A(G23), .B(G1976), .ZN(n910) );
  NOR2_X1 U1015 ( .A1(n911), .A2(n910), .ZN(n913) );
  XOR2_X1 U1016 ( .A(G1986), .B(G24), .Z(n912) );
  NAND2_X1 U1017 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1018 ( .A(KEYINPUT58), .B(n914), .ZN(n915) );
  NOR2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(n919), .B(KEYINPUT61), .ZN(n920) );
  XOR2_X1 U1022 ( .A(KEYINPUT125), .B(n920), .Z(n921) );
  NOR2_X1 U1023 ( .A1(G16), .A2(n921), .ZN(n1000) );
  XOR2_X1 U1024 ( .A(KEYINPUT56), .B(G16), .Z(n946) );
  XNOR2_X1 U1025 ( .A(n922), .B(G1348), .ZN(n923) );
  XNOR2_X1 U1026 ( .A(n923), .B(KEYINPUT123), .ZN(n944) );
  XOR2_X1 U1027 ( .A(G1341), .B(n924), .Z(n926) );
  NAND2_X1 U1028 ( .A1(G1971), .A2(G303), .ZN(n925) );
  NAND2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(G1966), .B(KEYINPUT122), .ZN(n927) );
  XNOR2_X1 U1031 ( .A(n927), .B(G168), .ZN(n929) );
  NAND2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(n930), .B(KEYINPUT57), .ZN(n938) );
  XOR2_X1 U1034 ( .A(G171), .B(G1961), .Z(n932) );
  XNOR2_X1 U1035 ( .A(G299), .B(G1956), .ZN(n931) );
  NOR2_X1 U1036 ( .A1(n932), .A2(n931), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n997) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n947) );
  NAND2_X1 U1045 ( .A1(n947), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G32), .B(n948), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n959) );
  XNOR2_X1 U1048 ( .A(n951), .B(G27), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(G2072), .B(KEYINPUT120), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(n952), .B(G33), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G26), .B(G2067), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(KEYINPUT121), .B(n955), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(n960), .B(KEYINPUT53), .ZN(n963) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(G35), .B(G2090), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(G29), .A2(n966), .ZN(n968) );
  XOR2_X1 U1063 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n967) );
  XNOR2_X1 U1064 ( .A(n968), .B(n967), .ZN(n995) );
  INV_X1 U1065 ( .A(n969), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n991) );
  XOR2_X1 U1067 ( .A(G2084), .B(G160), .Z(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n983) );
  XOR2_X1 U1071 ( .A(G2090), .B(KEYINPUT118), .Z(n978) );
  XNOR2_X1 U1072 ( .A(G162), .B(n978), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1074 ( .A(KEYINPUT51), .B(n981), .Z(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n989) );
  XOR2_X1 U1076 ( .A(G2072), .B(n984), .Z(n986) );
  XOR2_X1 U1077 ( .A(G164), .B(G2078), .Z(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1079 ( .A(KEYINPUT50), .B(n987), .Z(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT52), .B(n992), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(G29), .A2(n993), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n998), .A2(G11), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1002), .B(n1001), .ZN(G311) );
  XNOR2_X1 U1089 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

