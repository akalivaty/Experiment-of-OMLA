//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  AND2_X1   g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT0), .B(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n197), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n190), .A3(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT65), .B1(new_n188), .B2(G137), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n190), .A2(G134), .ZN(new_n212));
  OAI211_X1 g026(.A(G131), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n196), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n199), .B(new_n201), .C1(KEYINPUT1), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n200), .A2(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n198), .A2(G143), .ZN(new_n221));
  OAI211_X1 g035(.A(G128), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n218), .B(new_n222), .C1(new_n213), .C2(new_n214), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n208), .B(KEYINPUT30), .C1(new_n216), .C2(new_n223), .ZN(new_n224));
  OR2_X1    g038(.A1(KEYINPUT2), .A2(G113), .ZN(new_n225));
  AND3_X1   g039(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(G116), .B(G119), .Z(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G116), .B(G119), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(new_n225), .C1(new_n227), .C2(new_n226), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n206), .B1(new_n196), .B2(new_n194), .ZN(new_n234));
  INV_X1    g048(.A(new_n223), .ZN(new_n235));
  INV_X1    g049(.A(new_n193), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n236), .A2(new_n195), .B1(new_n213), .B2(new_n214), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n224), .B(new_n233), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n208), .B1(new_n216), .B2(new_n223), .ZN(new_n242));
  INV_X1    g056(.A(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n233), .A4(new_n224), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(G237), .A2(G953), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G210), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n242), .A2(new_n233), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n247), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT31), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n262));
  INV_X1    g076(.A(new_n233), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT72), .B1(new_n238), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n242), .A2(new_n265), .A3(new_n233), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n238), .A2(new_n263), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT71), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n255), .B(new_n262), .C1(new_n269), .C2(new_n260), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n247), .A2(new_n271), .A3(new_n257), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n259), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(G472), .A2(G902), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT32), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n273), .A2(KEYINPUT32), .A3(new_n274), .ZN(new_n278));
  INV_X1    g092(.A(new_n255), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n262), .C1(new_n269), .C2(new_n260), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n256), .B1(new_n241), .B2(new_n246), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n255), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT29), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n268), .A2(KEYINPUT28), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n242), .B(new_n263), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(KEYINPUT28), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n279), .A2(KEYINPUT29), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G472), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n277), .A2(new_n278), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G140), .ZN(new_n292));
  INV_X1    g106(.A(G125), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(KEYINPUT75), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(G125), .A3(G140), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(KEYINPUT16), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT16), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(new_n293), .B2(G140), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n198), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G125), .B(G140), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n198), .ZN(new_n303));
  XNOR2_X1  g117(.A(G119), .B(G128), .ZN(new_n304));
  INV_X1    g118(.A(G110), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(KEYINPUT24), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(KEYINPUT24), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT73), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT24), .B(G110), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n304), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(G128), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n315), .B(new_n316), .C1(G119), .C2(new_n217), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT76), .B(G110), .Z(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n301), .B(new_n303), .C1(new_n312), .C2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n308), .A2(new_n311), .A3(new_n304), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT74), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n308), .A2(new_n311), .A3(new_n323), .A4(new_n304), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n317), .A2(G110), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n297), .A2(new_n198), .A3(new_n299), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n328), .B2(new_n300), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n320), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT77), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT22), .B(G137), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n322), .A2(new_n324), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n301), .A2(new_n327), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n326), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n320), .A3(new_n335), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n284), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n337), .A2(KEYINPUT25), .A3(new_n284), .A4(new_n341), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G234), .ZN(new_n347));
  OAI21_X1  g161(.A(G217), .B1(new_n347), .B2(G902), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n340), .A2(new_n320), .A3(new_n335), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n335), .B1(new_n340), .B2(new_n320), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n349), .A2(G902), .ZN(new_n356));
  XOR2_X1   g170(.A(new_n356), .B(KEYINPUT78), .Z(new_n357));
  NOR2_X1   g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n350), .A2(new_n351), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n348), .B1(new_n344), .B2(new_n345), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT79), .B1(new_n361), .B2(new_n358), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT9), .B(G234), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n364), .A2(new_n365), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n284), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G221), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n370), .B(KEYINPUT81), .Z(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT90), .ZN(new_n374));
  INV_X1    g188(.A(G237), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n331), .A3(G214), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n200), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n248), .A2(G143), .A3(G214), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G131), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT17), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n379), .A2(KEYINPUT90), .A3(KEYINPUT17), .A4(G131), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n195), .A3(new_n378), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n380), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT91), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n328), .A2(new_n300), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n380), .A2(KEYINPUT91), .A3(new_n381), .A4(new_n385), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n384), .A2(new_n388), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G113), .B(G122), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n294), .A2(G146), .A3(new_n296), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n303), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT88), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT88), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n303), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT18), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n379), .A2(new_n401), .B1(new_n402), .B2(new_n195), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n195), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n377), .A2(KEYINPUT89), .A3(new_n404), .A4(new_n378), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n400), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n391), .A2(new_n394), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT19), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n302), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n294), .A2(KEYINPUT19), .A3(new_n296), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n198), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n380), .A2(new_n385), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n301), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n394), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n408), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G475), .A2(G902), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n373), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n419), .ZN(new_n421));
  AOI211_X1 g235(.A(KEYINPUT20), .B(new_n421), .C1(new_n408), .C2(new_n417), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n391), .A2(new_n407), .ZN(new_n423));
  INV_X1    g237(.A(new_n394), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(G902), .B1(new_n425), .B2(new_n408), .ZN(new_n426));
  INV_X1    g240(.A(G475), .ZN(new_n427));
  OAI22_X1  g241(.A1(new_n420), .A2(new_n422), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G478), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(KEYINPUT15), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n200), .A2(G128), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n217), .A2(G143), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n431), .A2(new_n432), .A3(new_n188), .ZN(new_n433));
  INV_X1    g247(.A(G122), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G116), .ZN(new_n435));
  INV_X1    g249(.A(G116), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G122), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G107), .ZN(new_n439));
  INV_X1    g253(.A(G107), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n433), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT13), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n431), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n432), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n431), .A2(new_n443), .ZN(new_n446));
  OAI21_X1  g260(.A(G134), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n436), .A2(KEYINPUT14), .A3(G122), .ZN(new_n449));
  OAI211_X1 g263(.A(G107), .B(new_n449), .C1(new_n438), .C2(KEYINPUT14), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n188), .B1(new_n431), .B2(new_n432), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n450), .B(new_n441), .C1(new_n433), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n331), .A2(G217), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n366), .A2(new_n367), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(new_n452), .A3(new_n455), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(KEYINPUT92), .ZN(new_n460));
  INV_X1    g274(.A(new_n458), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n455), .B1(new_n448), .B2(new_n452), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT92), .B(new_n284), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n430), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n331), .A2(G952), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n347), .B2(new_n375), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n284), .B(new_n331), .C1(G234), .C2(G237), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OAI22_X1  g286(.A1(new_n459), .A2(KEYINPUT92), .B1(KEYINPUT15), .B2(new_n429), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n428), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT83), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT3), .B1(new_n393), .B2(G107), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n440), .A3(G104), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n393), .A2(G107), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G101), .ZN(new_n482));
  INV_X1    g296(.A(G101), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n477), .A2(new_n479), .A3(new_n483), .A4(new_n480), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(KEYINPUT4), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n486), .A3(G101), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n207), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n440), .A2(KEYINPUT82), .A3(G104), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n393), .B2(G107), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n440), .A2(G104), .ZN(new_n492));
  OAI211_X1 g306(.A(G101), .B(new_n489), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n493), .A2(new_n484), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n494), .A2(KEYINPUT10), .A3(new_n218), .A4(new_n222), .ZN(new_n495));
  INV_X1    g309(.A(new_n197), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n493), .A2(new_n222), .A3(new_n484), .A4(new_n218), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT10), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n488), .A2(new_n495), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(new_n484), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n222), .A2(new_n218), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n497), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n504), .A2(KEYINPUT12), .A3(new_n197), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT12), .B1(new_n504), .B2(new_n197), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G110), .B(G140), .ZN(new_n508));
  INV_X1    g322(.A(G227), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(G953), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n508), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n511), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n500), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n488), .A2(new_n495), .A3(new_n499), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n197), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(G902), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G469), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n476), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n507), .A2(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n521));
  OAI211_X1 g335(.A(KEYINPUT83), .B(G469), .C1(new_n521), .C2(G902), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n500), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n511), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n504), .A2(new_n197), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n504), .A2(KEYINPUT12), .A3(new_n197), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n514), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n519), .A3(new_n284), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n520), .A2(new_n522), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(G214), .B1(G237), .B2(G902), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT84), .Z(new_n535));
  OAI21_X1  g349(.A(G210), .B1(G237), .B2(G902), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT86), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n537), .B(KEYINPUT87), .Z(new_n538));
  XNOR2_X1  g352(.A(G110), .B(G122), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n539), .B(KEYINPUT8), .Z(new_n540));
  INV_X1    g354(.A(KEYINPUT5), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n314), .A3(G116), .ZN(new_n542));
  OAI211_X1 g356(.A(G113), .B(new_n542), .C1(new_n229), .C2(new_n541), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n232), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n501), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n494), .A2(new_n232), .A3(new_n543), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n331), .A2(G224), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n207), .A2(G125), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n222), .A2(new_n293), .A3(new_n218), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n551), .A3(new_n549), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT85), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT85), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n550), .A2(new_n556), .A3(new_n551), .A4(new_n549), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n485), .A2(new_n233), .A3(new_n487), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n546), .A3(new_n539), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n284), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n546), .ZN(new_n563));
  INV_X1    g377(.A(new_n539), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT6), .A3(new_n560), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT6), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n550), .A2(new_n551), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n548), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n566), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n538), .B1(new_n562), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n555), .A2(new_n557), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n574), .A2(new_n552), .A3(new_n547), .ZN(new_n575));
  AOI21_X1  g389(.A(G902), .B1(new_n575), .B2(new_n560), .ZN(new_n576));
  INV_X1    g390(.A(new_n537), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n577), .A3(new_n571), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n535), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  AND4_X1   g393(.A1(new_n372), .A2(new_n475), .A3(new_n533), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n291), .A2(new_n363), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  INV_X1    g396(.A(KEYINPUT94), .ZN(new_n583));
  OAI21_X1  g397(.A(G469), .B1(new_n521), .B2(G902), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n511), .A2(new_n523), .B1(new_n514), .B2(new_n529), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(G902), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n584), .A2(new_n476), .B1(new_n586), .B2(new_n519), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n371), .B1(new_n587), .B2(new_n522), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n363), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n273), .A2(new_n284), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n591));
  INV_X1    g405(.A(G472), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n273), .B(new_n284), .C1(new_n591), .C2(new_n592), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n583), .B1(new_n589), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n360), .A2(new_n362), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n533), .A2(new_n372), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n600), .A2(KEYINPUT94), .A3(new_n595), .A4(new_n594), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n578), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n577), .B1(new_n576), .B2(new_n571), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n534), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n459), .A2(new_n429), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n429), .B2(new_n284), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n457), .A2(new_n458), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(KEYINPUT33), .Z(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n609), .B2(G478), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n428), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n605), .A2(new_n471), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  AOI22_X1  g429(.A1(new_n382), .A2(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n389), .A2(new_n390), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n616), .A2(new_n617), .B1(new_n400), .B2(new_n406), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n416), .B1(new_n618), .B2(new_n394), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT20), .B1(new_n619), .B2(new_n421), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n418), .A2(new_n373), .A3(new_n419), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n408), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n394), .B1(new_n391), .B2(new_n407), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n284), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(G475), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n465), .A2(new_n473), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n622), .A2(new_n626), .A3(new_n472), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT95), .ZN(new_n629));
  INV_X1    g443(.A(new_n534), .ZN(new_n630));
  INV_X1    g444(.A(new_n604), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(new_n631), .B2(new_n578), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n620), .A2(new_n621), .B1(new_n625), .B2(G475), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT95), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n633), .A2(new_n634), .A3(new_n472), .A4(new_n627), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n629), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n602), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT96), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT35), .B(G107), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  XNOR2_X1  g454(.A(new_n330), .B(KEYINPUT97), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n336), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n357), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n361), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n580), .A2(new_n595), .A3(new_n594), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n469), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n467), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n633), .A2(new_n627), .A3(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n605), .A2(new_n653), .A3(new_n645), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n291), .A2(new_n588), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n291), .A2(KEYINPUT98), .A3(new_n654), .A4(new_n588), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  XNOR2_X1  g474(.A(new_n652), .B(KEYINPUT39), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n588), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT40), .Z(new_n663));
  AND3_X1   g477(.A1(new_n273), .A2(KEYINPUT32), .A3(new_n274), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT32), .B1(new_n273), .B2(new_n274), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n281), .A2(new_n255), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n286), .A2(new_n255), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n284), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n428), .A2(new_n627), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n646), .A2(new_n630), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT99), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n573), .A2(new_n578), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n663), .A2(new_n671), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  AOI21_X1  g492(.A(new_n599), .B1(new_n666), .B2(new_n290), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n428), .A2(new_n610), .A3(new_n652), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n679), .A2(new_n632), .A3(new_n646), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  OAI21_X1  g497(.A(G469), .B1(new_n585), .B2(G902), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n532), .A3(new_n372), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n684), .A2(new_n532), .A3(KEYINPUT100), .A4(new_n372), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n291), .A2(new_n363), .A3(new_n612), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT101), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT41), .B(G113), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n291), .A2(new_n636), .A3(new_n363), .A4(new_n689), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  AND3_X1   g509(.A1(new_n632), .A2(new_n687), .A3(new_n688), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n645), .A2(new_n428), .A3(new_n474), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n291), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  AND3_X1   g513(.A1(new_n687), .A2(new_n472), .A3(new_n688), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n287), .A2(new_n255), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n259), .A2(new_n272), .A3(new_n701), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n590), .A2(G472), .B1(new_n274), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n605), .A2(new_n672), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n361), .A2(new_n358), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n700), .A2(new_n703), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NAND2_X1  g521(.A1(new_n703), .A2(new_n646), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n681), .A3(new_n696), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  NAND2_X1  g525(.A1(new_n584), .A2(new_n532), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n372), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n573), .A2(new_n578), .A3(new_n534), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n680), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AND4_X1   g529(.A1(KEYINPUT42), .A2(new_n291), .A3(new_n705), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n291), .A2(new_n363), .A3(new_n715), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT42), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n719), .B1(new_n718), .B2(new_n720), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n717), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G131), .ZN(G33));
  NOR3_X1   g538(.A1(new_n653), .A2(new_n713), .A3(new_n714), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n291), .A2(new_n363), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n188), .ZN(G36));
  OR2_X1    g541(.A1(new_n521), .A2(KEYINPUT45), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n521), .A2(KEYINPUT45), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(G469), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(G469), .A2(G902), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n532), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(new_n372), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n661), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT103), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n739), .A3(new_n661), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n633), .A2(new_n610), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT43), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n596), .A3(new_n646), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n714), .B1(new_n743), .B2(new_n744), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n738), .A2(new_n740), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT104), .B(G137), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G39));
  XNOR2_X1  g563(.A(new_n736), .B(KEYINPUT47), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n291), .A2(new_n363), .A3(new_n680), .A4(new_n714), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT105), .Z(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT106), .B(G140), .Z(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G42));
  XOR2_X1   g569(.A(new_n652), .B(KEYINPUT112), .Z(new_n756));
  NOR3_X1   g570(.A1(new_n646), .A2(new_n713), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n671), .A2(new_n704), .A3(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n659), .A2(new_n682), .A3(new_n710), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT52), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n696), .A2(new_n681), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n657), .A2(new_n658), .B1(new_n709), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n682), .A4(new_n758), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n718), .A2(new_n720), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT102), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n716), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n715), .A2(new_n703), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n291), .A2(new_n588), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n465), .A2(new_n473), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n652), .ZN(new_n775));
  OR3_X1    g589(.A1(new_n775), .A2(KEYINPUT110), .A3(new_n428), .ZN(new_n776));
  INV_X1    g590(.A(new_n714), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT110), .B1(new_n775), .B2(new_n428), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n772), .B1(new_n773), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n646), .ZN(new_n781));
  INV_X1    g595(.A(new_n726), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n771), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n428), .B2(new_n774), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n622), .A2(new_n626), .A3(KEYINPUT108), .A4(new_n627), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n579), .A3(new_n472), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n535), .B(new_n471), .C1(new_n573), .C2(new_n578), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(KEYINPUT109), .A3(new_n786), .A4(new_n787), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT107), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n611), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n428), .A2(KEYINPUT107), .A3(new_n610), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n790), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n597), .A2(new_n797), .A3(new_n601), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n581), .A2(new_n698), .A3(new_n647), .A4(new_n706), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n694), .A2(new_n690), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n767), .B1(new_n784), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n726), .B1(new_n780), .B2(new_n646), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n767), .A2(new_n801), .A3(new_n723), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n766), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n762), .A2(new_n763), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n798), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n799), .A2(new_n800), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n723), .A2(new_n809), .A3(new_n810), .A4(new_n803), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT111), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n801), .A2(new_n767), .A3(new_n723), .A4(new_n803), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n765), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n808), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT54), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n805), .A2(new_n818), .A3(new_n806), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT113), .B1(new_n814), .B2(KEYINPUT53), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n765), .A2(new_n821), .A3(new_n811), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n823), .A2(KEYINPUT54), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n468), .A2(new_n742), .A3(new_n689), .A4(new_n777), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n291), .A2(new_n705), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n705), .A2(new_n742), .A3(new_n468), .A4(new_n703), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n696), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n689), .A2(new_n777), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n671), .A2(new_n832), .A3(new_n598), .A4(new_n467), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n831), .B(new_n466), .C1(new_n834), .C2(new_n611), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n684), .A2(new_n532), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n372), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n777), .B(new_n830), .C1(new_n750), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n428), .A2(new_n610), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n833), .A2(new_n840), .B1(new_n825), .B2(new_n709), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n676), .A2(new_n534), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n830), .A2(new_n689), .A3(new_n843), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n844), .B(KEYINPUT50), .Z(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT51), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n836), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n845), .B(KEYINPUT114), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n848), .A2(new_n842), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n817), .A2(new_n824), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(G952), .B2(G953), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n371), .A2(new_n535), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n741), .A2(new_n705), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n837), .B(KEYINPUT49), .ZN(new_n856));
  OR3_X1    g670(.A1(new_n676), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n853), .B1(new_n671), .B2(new_n857), .ZN(G75));
  NAND2_X1  g672(.A1(new_n566), .A2(new_n568), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(new_n570), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT55), .Z(new_n861));
  NAND2_X1  g675(.A1(new_n823), .A2(G902), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n577), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(new_n863), .B2(KEYINPUT56), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n331), .A2(G952), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n823), .A2(KEYINPUT116), .A3(G902), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n538), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(G51));
  XNOR2_X1  g687(.A(new_n823), .B(KEYINPUT54), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n731), .B(KEYINPUT57), .Z(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n531), .ZN(new_n877));
  INV_X1    g691(.A(new_n730), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n869), .A2(new_n878), .A3(new_n870), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n865), .B1(new_n877), .B2(new_n879), .ZN(G54));
  AND2_X1   g694(.A1(KEYINPUT58), .A2(G475), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n869), .A2(new_n870), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT117), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n882), .A2(new_n883), .A3(new_n619), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n882), .B2(new_n619), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n869), .A2(new_n418), .A3(new_n870), .A4(new_n881), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n866), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(G60));
  INV_X1    g702(.A(new_n609), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n817), .A2(new_n824), .ZN(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n429), .A2(new_n284), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n889), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n874), .A2(new_n889), .A3(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n865), .ZN(G63));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT120), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT121), .Z(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT60), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n823), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n865), .B1(new_n903), .B2(new_n355), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n643), .B(KEYINPUT119), .Z(new_n905));
  NAND3_X1  g719(.A1(new_n823), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n897), .A2(KEYINPUT120), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n900), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n907), .B(new_n899), .C1(KEYINPUT120), .C2(new_n897), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(G66));
  INV_X1    g726(.A(new_n470), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n331), .B1(new_n913), .B2(G224), .ZN(new_n914));
  INV_X1    g728(.A(new_n801), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n331), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n859), .B1(G898), .B2(new_n331), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT122), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n916), .B(new_n918), .ZN(G69));
  NAND2_X1  g733(.A1(new_n794), .A2(new_n795), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n786), .A2(new_n787), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT124), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n662), .A2(new_n714), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(new_n291), .A3(new_n363), .A4(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n753), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n677), .A2(new_n682), .A3(new_n762), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(KEYINPUT62), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n926), .A2(new_n747), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n930), .A2(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(KEYINPUT125), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n331), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT123), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n244), .A2(new_n224), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(new_n412), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n509), .B2(new_n650), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT123), .B1(new_n933), .B2(new_n331), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n650), .A2(G953), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n738), .A2(new_n704), .A3(new_n826), .A4(new_n740), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n747), .A2(new_n753), .A3(new_n943), .A4(new_n782), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n723), .A2(new_n682), .A3(new_n762), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n942), .B1(new_n946), .B2(G953), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n937), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n948), .B2(new_n947), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n938), .B(new_n940), .C1(new_n941), .C2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n941), .A2(new_n950), .ZN(new_n952));
  INV_X1    g766(.A(new_n937), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n934), .B2(KEYINPUT123), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n939), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(G72));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n946), .B2(new_n801), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n866), .B1(new_n960), .B2(new_n282), .ZN(new_n961));
  INV_X1    g775(.A(new_n667), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n931), .A2(new_n801), .A3(new_n932), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n958), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n282), .A3(new_n958), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT127), .Z(new_n966));
  AOI211_X1 g780(.A(new_n961), .B(new_n964), .C1(new_n816), .C2(new_n966), .ZN(G57));
endmodule


