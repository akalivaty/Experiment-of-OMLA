//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g003(.A(G8gat), .B1(new_n204), .B2(KEYINPUT96), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G1gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n207), .B2(new_n202), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n205), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT14), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  INV_X1    g017(.A(G43gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(G50gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n220), .B2(KEYINPUT94), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n218), .ZN(new_n223));
  INV_X1    g022(.A(G50gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G43gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n217), .B(new_n221), .C1(new_n220), .C2(new_n225), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n230));
  OR2_X1    g029(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n229), .B2(new_n230), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n209), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n229), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n209), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n209), .B(new_n235), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n237), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n236), .A4(new_n237), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G169gat), .B(G197gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n245), .B(new_n251), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n254));
  NAND2_X1  g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255));
  INV_X1    g054(.A(G169gat), .ZN(new_n256));
  INV_X1    g055(.A(G176gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT26), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT27), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(G183gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(KEYINPUT27), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n259), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(KEYINPUT27), .ZN(new_n265));
  AOI21_X1  g064(.A(G190gat), .B1(new_n265), .B2(KEYINPUT68), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT28), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n268));
  NOR4_X1   g067(.A1(new_n261), .A2(new_n263), .A3(new_n268), .A4(G190gat), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n255), .B(new_n258), .C1(new_n267), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n256), .A2(new_n257), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT26), .ZN(new_n272));
  NAND2_X1  g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n254), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT24), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT66), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n255), .A2(new_n283), .A3(new_n277), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n279), .A2(new_n281), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n273), .B1(new_n271), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n286), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n293), .B(new_n273), .C1(new_n271), .C2(new_n286), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n295));
  AND4_X1   g094(.A1(KEYINPUT25), .A2(new_n294), .A3(new_n295), .A4(new_n289), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n255), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n280), .B1(new_n261), .B2(new_n259), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n260), .A2(G183gat), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT68), .B1(new_n265), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n268), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n261), .A2(new_n263), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT28), .A3(new_n280), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n300), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n307), .A2(KEYINPUT69), .A3(new_n274), .A4(new_n258), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n276), .A2(new_n299), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G134gat), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT71), .B1(new_n310), .B2(G127gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT70), .B(G127gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(new_n310), .ZN(new_n313));
  INV_X1    g112(.A(G127gat), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n314), .A2(KEYINPUT70), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(KEYINPUT70), .ZN(new_n316));
  OAI211_X1 g115(.A(KEYINPUT71), .B(G134gat), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318));
  INV_X1    g117(.A(G113gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(G120gat), .ZN(new_n320));
  INV_X1    g119(.A(G120gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(G113gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n313), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n325));
  XOR2_X1   g124(.A(G113gat), .B(G120gat), .Z(new_n326));
  NAND2_X1  g125(.A1(new_n310), .A2(G127gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n314), .A2(G134gat), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n326), .A2(new_n318), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n325), .B1(new_n324), .B2(new_n329), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n309), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n332), .A2(new_n276), .A3(new_n299), .A4(new_n308), .ZN(new_n335));
  NAND2_X1  g134(.A1(G227gat), .A2(G233gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT64), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT32), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT33), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G15gat), .B(G43gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(G71gat), .B(G99gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n334), .A2(new_n335), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT34), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n337), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n334), .A2(new_n335), .B1(G227gat), .B2(G233gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n345), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n339), .B(KEYINPUT32), .C1(new_n341), .C2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n346), .A2(new_n351), .A3(KEYINPUT73), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n353), .A2(new_n346), .B1(new_n351), .B2(KEYINPUT73), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT36), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n358));
  NAND2_X1  g157(.A1(new_n347), .A2(new_n336), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT34), .B1(new_n334), .B2(new_n335), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n359), .A2(KEYINPUT34), .B1(new_n360), .B2(new_n337), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n346), .A2(new_n361), .A3(new_n353), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n346), .B2(new_n353), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366));
  INV_X1    g165(.A(G64gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n368), .B(G92gat), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n374));
  NAND2_X1  g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n374), .B1(new_n373), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G197gat), .ZN(new_n379));
  INV_X1    g178(.A(G204gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G197gat), .A2(G204gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n381), .A2(new_n382), .B1(new_n383), .B2(new_n375), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT77), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n384), .C1(new_n376), .C2(new_n377), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n384), .B(KEYINPUT75), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n378), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(KEYINPUT29), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n309), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n307), .A2(new_n274), .A3(new_n258), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n299), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n393), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n392), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n299), .B1(new_n275), .B2(new_n270), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n394), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n276), .A2(new_n299), .A3(new_n308), .A4(new_n393), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n401), .A2(new_n402), .A3(new_n392), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n370), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n392), .A3(new_n402), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n309), .A2(new_n394), .B1(new_n397), .B2(new_n393), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n405), .B(new_n369), .C1(new_n406), .C2(new_n392), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(KEYINPUT30), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n406), .B2(new_n392), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n370), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n414));
  XNOR2_X1  g213(.A(G155gat), .B(G162gat), .ZN(new_n415));
  XOR2_X1   g214(.A(KEYINPUT78), .B(KEYINPUT2), .Z(new_n416));
  INV_X1    g215(.A(G148gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G141gat), .ZN(new_n418));
  INV_X1    g217(.A(G141gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G148gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT2), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT79), .B(G162gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(G155gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n421), .A2(new_n415), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n426), .A2(new_n427), .A3(KEYINPUT80), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT80), .ZN(new_n429));
  INV_X1    g228(.A(G162gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(G155gat), .ZN(new_n431));
  INV_X1    g230(.A(G155gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G162gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G141gat), .B(G148gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(KEYINPUT79), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G162gat), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n439), .A3(G155gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT2), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n429), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n423), .B1(new_n428), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n324), .A2(new_n329), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT80), .B1(new_n426), .B2(new_n427), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n436), .A2(new_n441), .A3(new_n429), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n422), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(new_n324), .A3(new_n329), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n451), .B(KEYINPUT81), .Z(new_n452));
  AOI21_X1  g251(.A(new_n414), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n448), .B1(new_n330), .B2(new_n331), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n454), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT82), .B1(new_n454), .B2(KEYINPUT4), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n449), .A2(KEYINPUT4), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n448), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n444), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n452), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n453), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n447), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n460), .B1(new_n466), .B2(new_n423), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT3), .B(new_n422), .C1(new_n446), .C2(new_n447), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT4), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n469), .A2(new_n444), .B1(new_n470), .B2(new_n454), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n448), .A2(KEYINPUT4), .A3(new_n324), .A4(new_n329), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n471), .A2(KEYINPUT83), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n454), .A2(new_n470), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(new_n462), .A3(new_n473), .A4(new_n472), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT83), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n465), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT0), .B(G57gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G85gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(G1gat), .B(G29gat), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n482), .B(new_n483), .Z(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT6), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT84), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n454), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT82), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n457), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n454), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n464), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n495), .A2(new_n453), .B1(new_n474), .B2(new_n478), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n487), .B1(new_n496), .B2(new_n484), .ZN(new_n497));
  AND4_X1   g296(.A1(new_n487), .A2(new_n465), .A3(new_n484), .A4(new_n479), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n486), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n496), .A2(new_n500), .A3(new_n484), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n413), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G78gat), .B(G106gat), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(G22gat), .Z(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT29), .B1(new_n448), .B2(new_n460), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT86), .B1(new_n507), .B2(new_n392), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n386), .A2(new_n388), .B1(new_n390), .B2(new_n378), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT86), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n509), .B(new_n510), .C1(new_n468), .C2(KEYINPUT29), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT3), .B1(new_n392), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n508), .B(new_n511), .C1(new_n513), .C2(new_n448), .ZN(new_n514));
  AND2_X1   g313(.A1(G228gat), .A2(G233gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(new_n224), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n386), .A2(new_n388), .B1(new_n378), .B2(new_n385), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n460), .B1(new_n520), .B2(KEYINPUT29), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n443), .ZN(new_n522));
  NAND2_X1  g321(.A1(G228gat), .A2(G233gat), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n522), .B(new_n523), .C1(new_n392), .C2(new_n507), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n519), .B1(new_n516), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n506), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n516), .A2(new_n524), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n518), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(new_n505), .A3(new_n525), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n365), .B1(new_n503), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT87), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT88), .B1(new_n496), .B2(new_n484), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT88), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n480), .A2(new_n536), .A3(new_n485), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n465), .A2(new_n479), .A3(new_n484), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT84), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n496), .A2(new_n487), .A3(new_n484), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n542), .A3(new_n500), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT90), .B(KEYINPUT37), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n409), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT37), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n545), .B(new_n369), .C1(new_n409), .C2(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n547), .A2(KEYINPUT38), .B1(new_n409), .B2(new_n370), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n406), .A2(new_n392), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n401), .A2(new_n402), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n549), .B(KEYINPUT37), .C1(new_n392), .C2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT38), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n551), .A2(new_n545), .A3(new_n552), .A4(new_n369), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n543), .A2(new_n502), .A3(new_n548), .A4(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n528), .A2(new_n531), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT40), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT39), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n450), .A2(new_n452), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n475), .A2(new_n462), .A3(new_n473), .ZN(new_n559));
  AOI211_X1 g358(.A(new_n557), .B(new_n558), .C1(new_n559), .C2(new_n452), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n557), .A3(new_n452), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n484), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n556), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n408), .A3(new_n411), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n564), .B1(new_n535), .B2(new_n537), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n560), .A2(new_n562), .A3(new_n556), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n555), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT87), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n571), .B(new_n365), .C1(new_n503), .C2(new_n532), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n534), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n346), .A2(new_n353), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n351), .A2(KEYINPUT73), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n354), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT92), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n532), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n532), .B2(new_n577), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n362), .B2(new_n363), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n574), .A2(new_n351), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n346), .A2(new_n361), .A3(new_n353), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(KEYINPUT91), .A3(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n584), .A2(new_n587), .A3(new_n532), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n543), .A2(new_n502), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n412), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n503), .A2(new_n582), .B1(new_n590), .B2(new_n581), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n253), .B1(new_n573), .B2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G57gat), .B(G64gat), .Z(new_n593));
  INV_X1    g392(.A(G71gat), .ZN(new_n594));
  INV_X1    g393(.A(G78gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n593), .B1(KEYINPUT9), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G71gat), .B(G78gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n209), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G183gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT97), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(new_n371), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n608), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n607), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n611), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n603), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n609), .A2(new_n611), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n619), .A3(new_n602), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT8), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT100), .B(G92gat), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n624), .B1(new_n625), .B2(G85gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n631));
  OR2_X1    g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n623), .ZN(new_n633));
  OR3_X1    g432(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n629), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT100), .B(G92gat), .Z(new_n636));
  INV_X1    g435(.A(G85gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n635), .A2(new_n638), .A3(new_n633), .A4(new_n624), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n623), .B(new_n632), .C1(new_n626), .C2(new_n629), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n640), .A3(new_n631), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n634), .A2(KEYINPUT102), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT102), .B1(new_n634), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n644), .A2(new_n229), .B1(KEYINPUT41), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n232), .A2(new_n233), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT103), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649));
  OAI221_X1 g448(.A(new_n649), .B1(new_n232), .B2(new_n233), .C1(new_n642), .C2(new_n643), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n280), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n645), .A2(KEYINPUT41), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT98), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G218gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n653), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n646), .A2(new_n648), .A3(new_n650), .A4(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n654), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n657), .B1(new_n654), .B2(new_n659), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n622), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n599), .A2(KEYINPUT10), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n642), .A2(new_n643), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n597), .B(new_n598), .Z(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n634), .A3(new_n641), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT10), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n599), .A2(new_n640), .A3(new_n639), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n665), .B1(new_n667), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n665), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n634), .A2(new_n641), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n634), .A2(KEYINPUT102), .A3(new_n641), .ZN(new_n680));
  INV_X1    g479(.A(new_n666), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n676), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT104), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n675), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n676), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(new_n257), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(new_n380), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n686), .A2(new_n688), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n684), .A2(new_n695), .ZN(new_n696));
  AOI211_X1 g495(.A(KEYINPUT105), .B(new_n676), .C1(new_n682), .C2(new_n683), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n692), .B1(new_n698), .B2(new_n688), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n664), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n592), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n501), .B1(new_n542), .B2(new_n486), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g504(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n706));
  OR2_X1    g505(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n702), .A2(new_n413), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n702), .ZN(new_n711));
  OAI21_X1  g510(.A(G8gat), .B1(new_n711), .B2(new_n412), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n709), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(G1325gat));
  NAND2_X1  g513(.A1(new_n584), .A2(new_n587), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(G15gat), .B1(new_n702), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n702), .A2(G15gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n585), .A2(new_n586), .ZN(new_n719));
  AOI22_X1  g518(.A1(KEYINPUT36), .A2(new_n577), .B1(new_n719), .B2(new_n358), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n717), .B1(new_n718), .B2(new_n720), .ZN(G1326gat));
  NAND2_X1  g520(.A1(new_n702), .A2(new_n555), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  INV_X1    g523(.A(new_n700), .ZN(new_n725));
  AND4_X1   g524(.A1(new_n592), .A2(new_n621), .A3(new_n662), .A4(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(new_n210), .A3(new_n703), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT45), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n621), .B(KEYINPUT106), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n729), .A2(new_n252), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n663), .A2(KEYINPUT44), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n500), .B1(new_n496), .B2(new_n484), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n540), .B2(new_n541), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n412), .B1(new_n734), .B2(new_n501), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n720), .B1(new_n555), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n570), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n590), .A2(new_n581), .ZN(new_n738));
  INV_X1    g537(.A(new_n580), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n532), .A2(new_n577), .A3(new_n578), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n739), .A2(new_n503), .A3(KEYINPUT35), .A4(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n737), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n591), .A2(KEYINPUT107), .A3(new_n737), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n732), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n573), .A2(new_n591), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n662), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n725), .B(new_n730), .C1(new_n746), .C2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n703), .ZN(new_n751));
  OAI21_X1  g550(.A(G29gat), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n728), .A2(new_n752), .ZN(G1328gat));
  NAND3_X1  g552(.A1(new_n726), .A2(new_n211), .A3(new_n413), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT46), .Z(new_n755));
  OAI21_X1  g554(.A(G36gat), .B1(new_n750), .B2(new_n412), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1329gat));
  NAND3_X1  g556(.A1(new_n726), .A2(new_n219), .A3(new_n716), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n726), .A2(KEYINPUT108), .A3(new_n219), .A4(new_n716), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G43gat), .B1(new_n750), .B2(new_n365), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(KEYINPUT47), .A3(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(G1330gat));
  OAI21_X1  g567(.A(G50gat), .B1(new_n750), .B2(new_n532), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n726), .A2(new_n224), .A3(new_n555), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT48), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n771), .B(new_n773), .ZN(G1331gat));
  NAND2_X1  g573(.A1(new_n744), .A2(new_n745), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n664), .A2(new_n252), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n775), .A2(new_n700), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n703), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n413), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT110), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n777), .A2(new_n783), .A3(new_n413), .A4(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1333gat));
  NAND3_X1  g586(.A1(new_n777), .A2(G71gat), .A3(new_n720), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n775), .A2(new_n700), .A3(new_n776), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n594), .B1(new_n789), .B2(new_n715), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g591(.A1(new_n789), .A2(new_n532), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(new_n595), .ZN(G1335gat));
  NOR3_X1   g593(.A1(new_n622), .A2(new_n252), .A3(new_n663), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n742), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(new_n742), .A3(KEYINPUT51), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n703), .A2(new_n700), .A3(new_n637), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT112), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT107), .B1(new_n591), .B2(new_n737), .ZN(new_n804));
  AND4_X1   g603(.A1(KEYINPUT107), .A2(new_n737), .A3(new_n738), .A4(new_n741), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n731), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT6), .B1(new_n540), .B2(new_n541), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n501), .B1(new_n807), .B2(new_n538), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n584), .A2(new_n587), .A3(new_n532), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n808), .A2(new_n809), .A3(new_n413), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n741), .B1(new_n810), .B2(KEYINPUT35), .ZN(new_n811));
  INV_X1    g610(.A(new_n572), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n555), .B1(new_n703), .B2(new_n413), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n571), .B1(new_n813), .B2(new_n365), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n811), .B1(new_n815), .B2(new_n570), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT44), .B1(new_n816), .B2(new_n663), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n806), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n622), .A2(new_n252), .A3(new_n725), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT111), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(KEYINPUT111), .B(new_n819), .C1(new_n746), .C2(new_n749), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n751), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n803), .B1(new_n823), .B2(new_n637), .ZN(G1336gat));
  AOI21_X1  g623(.A(new_n725), .B1(new_n798), .B2(new_n799), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(G92gat), .A3(new_n412), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n819), .B1(new_n746), .B2(new_n749), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n625), .B1(new_n829), .B2(new_n412), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n822), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n413), .B1(new_n820), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n827), .B1(new_n833), .B2(new_n625), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(G1337gat));
  XOR2_X1   g635(.A(KEYINPUT113), .B(G99gat), .Z(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n825), .A2(new_n716), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n365), .B1(new_n821), .B2(new_n822), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n838), .ZN(G1338gat));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n829), .B2(new_n532), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n818), .A2(KEYINPUT115), .A3(new_n555), .A4(new_n819), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(G106gat), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n847));
  INV_X1    g646(.A(G106gat), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n825), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n847), .B1(new_n849), .B2(new_n532), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n825), .A2(KEYINPUT114), .A3(new_n848), .A4(new_n555), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n845), .A2(new_n846), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n849), .A2(new_n532), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n555), .B1(new_n820), .B2(new_n832), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(G106gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n855), .B2(new_n846), .ZN(G1339gat));
  XNOR2_X1  g655(.A(new_n684), .B(new_n695), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n692), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n667), .A2(new_n672), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n860), .B2(new_n676), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n684), .A2(KEYINPUT104), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n674), .B(new_n676), .C1(new_n682), .C2(new_n683), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT116), .B1(new_n686), .B2(new_n861), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n859), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n859), .B(KEYINPUT55), .C1(new_n866), .C2(new_n867), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n871), .A2(KEYINPUT117), .A3(new_n693), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n871), .B2(new_n693), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n252), .B(new_n870), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n240), .A2(new_n243), .A3(new_n244), .A4(new_n251), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n237), .B1(new_n234), .B2(new_n236), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n241), .A2(new_n242), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n250), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n700), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n662), .B1(new_n874), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT118), .B1(new_n875), .B2(new_n878), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n660), .A2(new_n661), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n875), .A2(KEYINPUT118), .A3(new_n878), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n858), .B1(new_n696), .B2(new_n697), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n691), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n864), .A2(new_n865), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n686), .A2(KEYINPUT116), .A3(new_n861), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n882), .B(new_n883), .C1(new_n888), .C2(KEYINPUT55), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n871), .A2(new_n693), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n871), .A2(KEYINPUT117), .A3(new_n693), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n729), .B1(new_n880), .B2(new_n894), .ZN(new_n895));
  NOR4_X1   g694(.A1(new_n621), .A2(new_n252), .A3(new_n662), .A4(new_n700), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n751), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n579), .A2(new_n580), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n898), .A2(new_n412), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n319), .A3(new_n252), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n895), .A2(new_n897), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n902), .A2(new_n703), .A3(new_n588), .A4(new_n412), .ZN(new_n903));
  OAI21_X1  g702(.A(G113gat), .B1(new_n903), .B2(new_n253), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1340gat));
  NAND3_X1  g704(.A1(new_n900), .A2(new_n321), .A3(new_n700), .ZN(new_n906));
  OAI21_X1  g705(.A(G120gat), .B1(new_n903), .B2(new_n725), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1341gat));
  INV_X1    g707(.A(new_n312), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n903), .A2(new_n909), .A3(new_n729), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n900), .A2(new_n622), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n909), .ZN(G1342gat));
  NAND3_X1  g711(.A1(new_n900), .A2(new_n310), .A3(new_n662), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n914));
  OAI21_X1  g713(.A(G134gat), .B1(new_n903), .B2(new_n663), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(G1343gat));
  AOI21_X1  g716(.A(new_n532), .B1(new_n895), .B2(new_n897), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n720), .A2(new_n751), .A3(new_n413), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n252), .B1(new_n888), .B2(KEYINPUT55), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n879), .B1(new_n923), .B2(new_n890), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n663), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n886), .A2(new_n887), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT55), .B1(new_n926), .B2(new_n859), .ZN(new_n927));
  OR3_X1    g726(.A1(new_n660), .A2(new_n661), .A3(new_n881), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n929), .B(new_n883), .C1(new_n872), .C2(new_n873), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n622), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n555), .B1(new_n931), .B2(new_n896), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n922), .B1(new_n932), .B2(KEYINPUT57), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n920), .A2(new_n252), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G141gat), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n918), .A2(new_n419), .A3(new_n252), .A4(new_n921), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(KEYINPUT120), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(KEYINPUT120), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n935), .A2(new_n936), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n936), .A2(KEYINPUT119), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n918), .A2(new_n921), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n942), .A2(new_n943), .A3(new_n419), .A4(new_n252), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n935), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n945), .B2(new_n937), .ZN(G1344gat));
  NOR4_X1   g745(.A1(new_n725), .A2(G148gat), .A3(new_n532), .A4(new_n413), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n898), .A2(new_n365), .A3(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n920), .A2(new_n933), .ZN(new_n949));
  AOI211_X1 g748(.A(KEYINPUT59), .B(new_n417), .C1(new_n949), .C2(new_n700), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n870), .A2(new_n252), .A3(new_n693), .A4(new_n871), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n662), .B1(new_n953), .B2(new_n879), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n954), .B2(new_n894), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n925), .A2(KEYINPUT121), .A3(new_n930), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n956), .A3(new_n621), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n897), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n957), .A2(KEYINPUT122), .A3(new_n897), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n960), .A2(new_n919), .A3(new_n555), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n902), .A2(new_n555), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT57), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n962), .A2(new_n964), .A3(new_n700), .A4(new_n921), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n951), .B1(new_n965), .B2(G148gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n948), .B1(new_n950), .B2(new_n966), .ZN(G1345gat));
  NAND2_X1  g766(.A1(new_n918), .A2(new_n921), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n968), .A2(new_n621), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT123), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n729), .A2(new_n432), .ZN(new_n971));
  AOI22_X1  g770(.A1(new_n970), .A2(new_n432), .B1(new_n949), .B2(new_n971), .ZN(G1346gat));
  AOI21_X1  g771(.A(new_n425), .B1(new_n942), .B2(new_n662), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n949), .A2(new_n425), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n974), .B2(new_n662), .ZN(G1347gat));
  NOR2_X1   g774(.A1(new_n703), .A2(new_n412), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n977), .B1(new_n895), .B2(new_n897), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n978), .A2(new_n899), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n979), .A2(new_n256), .A3(new_n252), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT124), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n978), .A2(new_n588), .ZN(new_n982));
  OAI21_X1  g781(.A(G169gat), .B1(new_n982), .B2(new_n253), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1348gat));
  AOI21_X1  g783(.A(G176gat), .B1(new_n979), .B2(new_n700), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n982), .A2(new_n257), .A3(new_n725), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(G1349gat));
  NOR2_X1   g786(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n988));
  AND2_X1   g787(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n979), .A2(new_n305), .A3(new_n622), .ZN(new_n990));
  OAI21_X1  g789(.A(G183gat), .B1(new_n982), .B2(new_n729), .ZN(new_n991));
  AOI211_X1 g790(.A(new_n988), .B(new_n989), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  AND4_X1   g791(.A1(KEYINPUT125), .A2(new_n990), .A3(KEYINPUT60), .A4(new_n991), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n992), .A2(new_n993), .ZN(G1350gat));
  OAI21_X1  g793(.A(G190gat), .B1(new_n982), .B2(new_n663), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT126), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g796(.A(KEYINPUT126), .B(G190gat), .C1(new_n982), .C2(new_n663), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(KEYINPUT61), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n979), .A2(new_n280), .A3(new_n662), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n995), .A2(new_n996), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(G1351gat));
  NOR2_X1   g802(.A1(new_n977), .A2(new_n720), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n918), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1005), .A2(new_n379), .A3(new_n252), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n961), .A2(new_n555), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT57), .B1(new_n958), .B2(new_n959), .ZN(new_n1008));
  AOI22_X1  g807(.A1(new_n1007), .A2(new_n1008), .B1(new_n963), .B2(KEYINPUT57), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n1009), .A2(new_n252), .A3(new_n1004), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1006), .B1(new_n1010), .B2(new_n379), .ZN(G1352gat));
  NAND4_X1  g810(.A1(new_n962), .A2(new_n964), .A3(new_n700), .A4(new_n1004), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(KEYINPUT127), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1014));
  NAND4_X1  g813(.A1(new_n1009), .A2(new_n1014), .A3(new_n700), .A4(new_n1004), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1013), .A2(new_n1015), .A3(G204gat), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1005), .A2(new_n380), .A3(new_n700), .ZN(new_n1017));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1016), .A2(new_n1019), .ZN(G1353gat));
  NAND3_X1  g819(.A1(new_n1005), .A2(new_n371), .A3(new_n622), .ZN(new_n1021));
  NAND4_X1  g820(.A1(new_n962), .A2(new_n964), .A3(new_n622), .A4(new_n1004), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1022), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1023));
  AOI21_X1  g822(.A(KEYINPUT63), .B1(new_n1022), .B2(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(G1354gat));
  NAND3_X1  g824(.A1(new_n1005), .A2(new_n372), .A3(new_n662), .ZN(new_n1026));
  AND3_X1   g825(.A1(new_n1009), .A2(new_n662), .A3(new_n1004), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1026), .B1(new_n1027), .B2(new_n372), .ZN(G1355gat));
endmodule


