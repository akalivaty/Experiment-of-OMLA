//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  NAND2_X1  g046(.A1(new_n463), .A2(G136), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n462), .A2(new_n464), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G162));
  NOR2_X1   g053(.A1(new_n464), .A2(G114), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT65), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OR3_X1    g056(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT65), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(new_n482), .B1(new_n473), .B2(G126), .ZN(new_n483));
  OAI211_X1 g058(.A(G138), .B(new_n464), .C1(new_n460), .C2(new_n461), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G164));
  INV_X1    g062(.A(KEYINPUT5), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G543), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n490));
  INV_X1    g065(.A(G543), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT5), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(KEYINPUT67), .A3(G543), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT6), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G651), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(KEYINPUT66), .A3(KEYINPUT6), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n501), .A3(G88), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(G50), .A3(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(G75), .A2(G543), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n494), .B2(G62), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n502), .B(new_n503), .C1(new_n505), .C2(new_n495), .ZN(G303));
  INV_X1    g081(.A(G303), .ZN(G166));
  NAND2_X1  g082(.A1(new_n491), .A2(KEYINPUT5), .ZN(new_n508));
  AND2_X1   g083(.A1(G63), .A2(G651), .ZN(new_n509));
  AND3_X1   g084(.A1(new_n488), .A2(KEYINPUT67), .A3(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(KEYINPUT67), .B1(new_n488), .B2(G543), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT68), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n494), .A2(new_n514), .A3(new_n509), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT69), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n519), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n494), .A2(new_n501), .A3(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n501), .A2(G51), .A3(G543), .ZN(new_n524));
  AND4_X1   g099(.A1(new_n516), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(G168));
  NAND3_X1  g100(.A1(new_n494), .A2(new_n501), .A3(G90), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n501), .A2(G52), .A3(G543), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n528), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  INV_X1    g105(.A(G77), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n491), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(new_n494), .B2(G64), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n534));
  OAI21_X1  g109(.A(G651), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI211_X1 g110(.A(KEYINPUT70), .B(new_n532), .C1(new_n494), .C2(G64), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n529), .A2(new_n530), .B1(new_n535), .B2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND3_X1  g113(.A1(new_n494), .A2(new_n501), .A3(G81), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n501), .A2(G43), .A3(G543), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g116(.A(G56), .B(new_n508), .C1(new_n510), .C2(new_n511), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n495), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(KEYINPUT72), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n539), .A2(new_n540), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n548));
  NOR3_X1   g123(.A1(new_n547), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g127(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n553));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT74), .Z(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT76), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n560));
  XNOR2_X1  g135(.A(KEYINPUT77), .B(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n494), .A2(new_n501), .ZN(new_n563));
  AOI22_X1  g138(.A1(G651), .A2(new_n562), .B1(new_n563), .B2(G91), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n501), .A2(G53), .A3(G543), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(KEYINPUT75), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n567), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n501), .A2(G53), .A3(G543), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n564), .A2(new_n571), .ZN(G299));
  NAND4_X1  g147(.A1(new_n516), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(G286));
  NAND3_X1  g148(.A1(new_n501), .A2(G49), .A3(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT78), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n501), .A2(new_n576), .A3(G49), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n494), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n494), .A2(new_n501), .A3(G87), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n494), .A2(new_n501), .A3(G86), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n501), .A2(G48), .A3(G543), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g160(.A(G61), .B(new_n508), .C1(new_n510), .C2(new_n511), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(KEYINPUT79), .B1(new_n588), .B2(G651), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n590));
  AOI211_X1 g165(.A(new_n590), .B(new_n495), .C1(new_n586), .C2(new_n587), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n585), .B1(new_n589), .B2(new_n591), .ZN(G305));
  NAND3_X1  g167(.A1(new_n494), .A2(new_n501), .A3(G85), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n501), .A2(G47), .A3(G543), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n494), .B2(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n598), .B2(KEYINPUT80), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  AOI211_X1 g175(.A(new_n600), .B(new_n597), .C1(new_n494), .C2(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n599), .B2(new_n601), .ZN(G290));
  NAND3_X1  g177(.A1(new_n563), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n494), .A2(new_n501), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT81), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n560), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n501), .A2(G543), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n612), .A2(G651), .B1(new_n613), .B2(G54), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n615), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g191(.A(new_n615), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(new_n615), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n550), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n626), .A2(new_n625), .A3(G868), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n628), .A2(new_n629), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g206(.A(new_n462), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(new_n465), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n463), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n473), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n464), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n637), .A2(new_n638), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT83), .Z(G156));
  XOR2_X1   g221(.A(KEYINPUT15), .B(G2435), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2438), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT85), .B(KEYINPUT14), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT86), .Z(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n666), .A2(new_n667), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n671), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n682), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(KEYINPUT20), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n683), .B1(new_n680), .B2(new_n684), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G23), .ZN(new_n700));
  INV_X1    g275(.A(G288), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n699), .A2(KEYINPUT89), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(KEYINPUT89), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G22), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n699), .A2(G6), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G305), .B2(G16), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n704), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n713), .A2(new_n714), .ZN(new_n717));
  OR3_X1    g292(.A1(new_n716), .A2(KEYINPUT34), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(KEYINPUT34), .B1(new_n716), .B2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n463), .A2(G131), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n473), .A2(G119), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n464), .A2(G107), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G25), .B(new_n724), .S(G29), .Z(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT35), .B(G1991), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n725), .B(new_n726), .Z(new_n727));
  MUX2_X1   g302(.A(G24), .B(G290), .S(new_n707), .Z(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(G1986), .Z(new_n729));
  NAND4_X1  g304(.A1(new_n718), .A2(new_n719), .A3(new_n727), .A4(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT36), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(G168), .A2(G16), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n734), .B(new_n735), .C1(G16), .C2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT96), .B(G1966), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT97), .Z(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n742), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT29), .Z(new_n745));
  INV_X1    g320(.A(G2090), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G4), .A2(G16), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n622), .B2(G16), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n747), .A2(KEYINPUT100), .B1(G1348), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(KEYINPUT100), .B2(new_n747), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n737), .A2(new_n739), .ZN(new_n752));
  INV_X1    g327(.A(new_n707), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G20), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT23), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n619), .B2(new_n699), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT101), .B(G1956), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G5), .A2(G16), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT99), .Z(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G301), .B2(new_n699), .ZN(new_n761));
  INV_X1    g336(.A(G1961), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n752), .A2(new_n758), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n742), .A2(G33), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n632), .A2(G127), .ZN(new_n767));
  AND2_X1   g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(G2105), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n770));
  NAND2_X1  g345(.A1(G103), .A2(G2104), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G2105), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n463), .A2(G139), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n766), .B1(new_n775), .B2(G29), .ZN(new_n776));
  INV_X1    g351(.A(G2072), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n742), .B1(new_n779), .B2(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n779), .B2(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G160), .B2(G29), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n782), .A2(G2084), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(G2084), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n778), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n742), .A2(G27), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G164), .B2(new_n742), .ZN(new_n787));
  INV_X1    g362(.A(G2078), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n785), .B(new_n789), .C1(new_n745), .C2(new_n746), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n742), .A2(G32), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n465), .A2(G105), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n463), .A2(G141), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n473), .A2(G129), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n791), .B1(new_n800), .B2(new_n742), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT27), .B(G1996), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT94), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT93), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n801), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n742), .A2(G26), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT28), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n463), .A2(G140), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n473), .A2(G128), .ZN(new_n809));
  OR2_X1    g384(.A1(G104), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(new_n742), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G2067), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n749), .A2(G1348), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT31), .B(G11), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT30), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n742), .B1(new_n818), .B2(G28), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(KEYINPUT98), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(G28), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n819), .B2(KEYINPUT98), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n817), .B1(new_n820), .B2(new_n822), .C1(new_n643), .C2(new_n742), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n776), .B2(new_n777), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n805), .A2(new_n815), .A3(new_n816), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n753), .A2(G19), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n550), .B2(new_n753), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT91), .B(G1341), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n790), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n741), .A2(new_n751), .A3(new_n765), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n733), .A2(new_n831), .ZN(G311));
  INV_X1    g407(.A(G311), .ZN(G150));
  NAND2_X1  g408(.A1(new_n494), .A2(G67), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n495), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n501), .A2(G55), .A3(G543), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n605), .B2(new_n838), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n546), .A2(new_n549), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n836), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(new_n545), .A3(new_n541), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n615), .A2(new_n623), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  INV_X1    g422(.A(G860), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n841), .A2(new_n848), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(G145));
  XNOR2_X1  g430(.A(new_n800), .B(new_n812), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(new_n486), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n486), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n775), .A2(KEYINPUT103), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n775), .A2(KEYINPUT103), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n857), .A2(new_n860), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n473), .A2(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n464), .A2(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G142), .B2(new_n463), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n634), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(new_n724), .Z(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n863), .A2(new_n872), .A3(new_n864), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(KEYINPUT104), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n865), .A2(new_n877), .A3(new_n873), .ZN(new_n878));
  XOR2_X1   g453(.A(G160), .B(new_n643), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n477), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n872), .A2(KEYINPUT105), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n865), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n880), .B1(new_n865), .B2(new_n882), .ZN(new_n884));
  AOI21_X1  g459(.A(G37), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g462(.A1(G290), .A2(G288), .ZN(new_n888));
  INV_X1    g463(.A(G60), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n596), .B1(new_n560), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n600), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n598), .A2(KEYINPUT80), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(G651), .A3(new_n892), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n893), .A2(new_n595), .B1(new_n578), .B2(new_n581), .ZN(new_n894));
  OAI211_X1 g469(.A(G303), .B(new_n585), .C1(new_n589), .C2(new_n591), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n587), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n494), .B2(G61), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n590), .B1(new_n898), .B2(new_n495), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n588), .A2(KEYINPUT79), .A3(G651), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G303), .B1(new_n901), .B2(new_n585), .ZN(new_n902));
  OAI22_X1  g477(.A1(new_n888), .A2(new_n894), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(G305), .A2(G166), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n893), .A2(new_n578), .A3(new_n581), .A4(new_n595), .ZN(new_n905));
  NAND2_X1  g480(.A1(G290), .A2(G288), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n895), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT107), .B1(new_n903), .B2(new_n907), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT108), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n843), .B(new_n626), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n608), .A2(new_n564), .A3(new_n614), .A4(new_n571), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n608), .A2(new_n614), .B1(new_n564), .B2(new_n571), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n615), .A2(G299), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(KEYINPUT41), .A3(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OR3_X1    g496(.A1(new_n913), .A2(KEYINPUT106), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT106), .B1(new_n913), .B2(new_n921), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n915), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n913), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n928));
  INV_X1    g503(.A(new_n907), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n906), .A2(new_n905), .B1(new_n904), .B2(new_n895), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n912), .A2(new_n927), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n927), .B1(new_n912), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g510(.A(new_n934), .B1(G868), .B2(new_n841), .ZN(G331));
  NOR2_X1   g511(.A1(G301), .A2(G168), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n526), .A2(new_n527), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT71), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G64), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n560), .A2(new_n942), .B1(new_n531), .B2(new_n491), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT70), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n533), .A2(new_n534), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(G651), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G286), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n541), .A2(new_n545), .A3(KEYINPUT72), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n548), .B1(new_n547), .B2(new_n544), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n841), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR4_X1   g525(.A1(new_n836), .A2(new_n839), .A3(new_n547), .A4(new_n544), .ZN(new_n951));
  OAI22_X1  g526(.A1(new_n937), .A2(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(G301), .A2(G168), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n941), .A2(new_n946), .A3(G286), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n840), .A2(new_n953), .A3(new_n842), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n925), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n929), .B2(new_n930), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n952), .A2(new_n918), .A3(new_n955), .A4(new_n920), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n907), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n957), .A2(new_n959), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G37), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n924), .B1(new_n952), .B2(new_n955), .ZN(new_n966));
  INV_X1    g541(.A(new_n921), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n952), .A2(new_n955), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n965), .B1(new_n969), .B2(new_n910), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n957), .A2(new_n960), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n959), .A2(new_n961), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(KEYINPUT111), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n964), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT43), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n969), .B2(new_n910), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n969), .A2(new_n910), .A3(new_n965), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT111), .B1(new_n971), .B2(new_n972), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n975), .B(new_n977), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT113), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT112), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n984), .A2(new_n985), .A3(KEYINPUT43), .A4(new_n980), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n964), .B1(new_n972), .B2(new_n971), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n989));
  AOI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n982), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n974), .A2(new_n989), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n987), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n991), .A2(new_n995), .ZN(G397));
  AND3_X1   g571(.A1(new_n466), .A2(new_n470), .A3(G40), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n483), .B2(new_n485), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n998), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n812), .B(G2067), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT115), .Z(new_n1002));
  INV_X1    g577(.A(G1996), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n800), .B(new_n1003), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n1000), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT116), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1008), .A3(new_n1000), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n724), .A2(new_n726), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n812), .A2(G2067), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1000), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n800), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1000), .B1(new_n1002), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT46), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1000), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1018), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1015), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1021));
  XNOR2_X1  g596(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1013), .A2(new_n1022), .ZN(new_n1023));
  OR3_X1    g598(.A1(new_n1018), .A2(G1986), .A3(G290), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n1024), .B(KEYINPUT48), .Z(new_n1025));
  AND2_X1   g600(.A1(new_n724), .A2(new_n726), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1000), .B1(new_n1010), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1007), .A2(new_n1009), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT126), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1007), .A2(KEYINPUT126), .A3(new_n1009), .A4(new_n1027), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1025), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1023), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n999), .A2(new_n997), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G8), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(G305), .A2(G1981), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n585), .B1(new_n495), .B2(new_n898), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G1981), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1037), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n701), .A2(G1976), .ZN(new_n1046));
  INV_X1    g621(.A(G1976), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1037), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT119), .B1(new_n1034), .B2(G8), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1045), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n999), .A2(KEYINPUT45), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n997), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n710), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n999), .A2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT117), .B(G2090), .Z(new_n1063));
  NAND4_X1  g638(.A1(new_n1060), .A2(new_n997), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1055), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  XOR2_X1   g643(.A(new_n1068), .B(KEYINPUT55), .Z(new_n1069));
  NAND3_X1  g644(.A1(new_n1059), .A2(new_n1064), .A3(KEYINPUT118), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1055), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1072), .A2(new_n1069), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1054), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1075), .A2(KEYINPUT53), .A3(new_n788), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1062), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n997), .B1(new_n999), .B2(new_n1061), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n762), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1057), .A2(new_n1058), .A3(G2078), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1082), .A2(KEYINPUT53), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1077), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1085));
  OAI21_X1  g660(.A(G171), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1074), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n738), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1088));
  INV_X1    g663(.A(G2084), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1060), .A2(new_n1089), .A3(new_n997), .A4(new_n1062), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1090), .A3(G168), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(G168), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT51), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(G8), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1097), .B2(KEYINPUT62), .ZN(new_n1102));
  AOI211_X1 g677(.A(KEYINPUT124), .B(new_n1099), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1087), .B(new_n1100), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1074), .A2(new_n1098), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1058), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1056), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G299), .B(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(G1348), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1034), .A2(G2067), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1115), .B1(new_n1119), .B2(new_n615), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1108), .A2(new_n1113), .A3(new_n1110), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1121), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1113), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1115), .A2(KEYINPUT61), .A3(new_n1121), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1119), .A2(KEYINPUT60), .ZN(new_n1128));
  OAI221_X1 g703(.A(KEYINPUT60), .B1(G2067), .B2(new_n1034), .C1(new_n1116), .C2(G1348), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n622), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1126), .B(new_n1127), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1057), .A2(new_n1058), .A3(G1996), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT58), .B(G1341), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1133), .B1(new_n999), .B2(new_n997), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n550), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(KEYINPUT59), .B(new_n550), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1137), .B(new_n1138), .C1(new_n622), .C2(new_n1129), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1122), .B1(new_n1131), .B2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1106), .A2(KEYINPUT122), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1106), .A2(KEYINPUT122), .ZN(new_n1142));
  NAND2_X1  g717(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1143));
  OR2_X1    g718(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1144));
  AND4_X1   g719(.A1(KEYINPUT53), .A2(new_n1056), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1083), .A2(new_n1146), .A3(G301), .A4(new_n1080), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1086), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1083), .A2(new_n1146), .A3(new_n1080), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1149), .B1(new_n1151), .B2(G171), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1153), .B2(G171), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1105), .A2(new_n1140), .A3(new_n1150), .A4(new_n1154), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1055), .B(G286), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1156), .B(new_n1157), .C1(new_n1069), .C2(new_n1072), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1071), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1054), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1045), .A2(new_n1047), .A3(new_n701), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1038), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1037), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1045), .A2(new_n1049), .A3(new_n1156), .A4(new_n1053), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1069), .A2(KEYINPUT120), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1067), .A2(KEYINPUT120), .A3(new_n1070), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1157), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1104), .A2(new_n1155), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1000), .A2(G1986), .A3(G290), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1024), .A2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT114), .Z(new_n1175));
  OR2_X1    g750(.A1(new_n1028), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1033), .B1(new_n1172), .B2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g752(.A1(G227), .A2(new_n458), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n1179), .A2(new_n663), .ZN(new_n1180));
  INV_X1    g754(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g755(.A(KEYINPUT127), .B1(new_n697), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n1183));
  AOI211_X1 g757(.A(new_n1183), .B(new_n1180), .C1(new_n695), .C2(new_n696), .ZN(new_n1184));
  OAI211_X1 g758(.A(new_n994), .B(new_n886), .C1(new_n1182), .C2(new_n1184), .ZN(G225));
  INV_X1    g759(.A(G225), .ZN(G308));
endmodule


