//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT68), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT69), .ZN(new_n204));
  XOR2_X1   g003(.A(G71gat), .B(G99gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n208), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n212), .B(new_n215), .C1(new_n211), .C2(new_n210), .ZN(new_n216));
  NOR2_X1   g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  NOR3_X1   g016(.A1(new_n213), .A2(new_n217), .A3(new_n214), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT64), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT27), .B(G183gat), .ZN(new_n221));
  INV_X1    g020(.A(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n210), .B1(new_n209), .B2(KEYINPUT26), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n210), .A2(KEYINPUT26), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n213), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n219), .A2(new_n220), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(new_n220), .B2(new_n219), .ZN(new_n230));
  XNOR2_X1  g029(.A(G113gat), .B(G120gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  INV_X1    g031(.A(G127gat), .ZN(new_n233));
  INV_X1    g032(.A(G134gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G127gat), .A2(G134gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n235), .B(new_n236), .C1(KEYINPUT66), .C2(KEYINPUT1), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n232), .B(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G227gat), .ZN(new_n242));
  INV_X1    g041(.A(G233gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n206), .B1(new_n245), .B2(KEYINPUT32), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT33), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(KEYINPUT67), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249));
  INV_X1    g048(.A(new_n244), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n239), .B2(new_n240), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n249), .B1(new_n251), .B2(KEYINPUT33), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n206), .B(KEYINPUT70), .Z(new_n254));
  OAI211_X1 g053(.A(KEYINPUT32), .B(new_n245), .C1(new_n254), .C2(new_n247), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n250), .A3(new_n240), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(KEYINPUT34), .Z(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n253), .A2(new_n258), .A3(new_n255), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT36), .ZN(new_n263));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G155gat), .B(G162gat), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G141gat), .B(G148gat), .Z(new_n268));
  INV_X1    g067(.A(G155gat), .ZN(new_n269));
  INV_X1    g068(.A(G162gat), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT2), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n266), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G197gat), .B(G204gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT72), .B(G218gat), .ZN(new_n281));
  INV_X1    g080(.A(G211gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n279), .A2(new_n280), .B1(new_n283), .B2(KEYINPUT22), .ZN(new_n284));
  XOR2_X1   g083(.A(G211gat), .B(G218gat), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n277), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n284), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT29), .B1(new_n277), .B2(new_n289), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G228gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(new_n243), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n294), .B2(new_n295), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n289), .B1(new_n293), .B2(KEYINPUT29), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n301), .B1(new_n276), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(G22gat), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n300), .A2(new_n303), .A3(G22gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n265), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n306), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n304), .A3(new_n264), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT31), .B(G50gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n311), .B(KEYINPUT79), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n307), .A2(new_n309), .A3(new_n312), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT36), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n260), .A2(new_n317), .A3(new_n261), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n263), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT74), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(new_n230), .B2(new_n287), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n320), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n322), .A2(new_n323), .B1(new_n230), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n294), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n325), .B1(new_n230), .B2(new_n287), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n230), .B2(new_n321), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n294), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT30), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n324), .A2(new_n326), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n293), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n294), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n338), .A4(new_n334), .ZN(new_n339));
  INV_X1    g138(.A(new_n338), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n333), .B1(new_n340), .B2(new_n327), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n277), .A2(new_n289), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n238), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n238), .A2(new_n276), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT4), .ZN(new_n350));
  OR3_X1    g149(.A1(new_n238), .A2(new_n276), .A3(KEYINPUT4), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT78), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n354), .A3(new_n351), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n348), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357));
  OR3_X1    g156(.A1(new_n356), .A2(KEYINPUT39), .A3(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT0), .ZN(new_n360));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  XNOR2_X1  g161(.A(new_n277), .B(new_n238), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n357), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT39), .B(new_n364), .C1(new_n356), .C2(new_n357), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n358), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT40), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT80), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n369), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n373));
  INV_X1    g172(.A(new_n351), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n347), .A2(new_n357), .ZN(new_n376));
  OAI221_X1 g175(.A(KEYINPUT5), .B1(new_n357), .B2(new_n363), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT5), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n356), .A2(new_n378), .A3(new_n357), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n362), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n371), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n343), .A2(new_n344), .A3(new_n370), .A4(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n335), .A2(new_n342), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n382), .A3(new_n371), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT81), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT37), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n334), .B1(new_n330), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n389), .B2(new_n330), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT38), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n362), .A3(new_n379), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n382), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT6), .A3(new_n381), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n336), .A2(new_n294), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n389), .B1(new_n329), .B2(new_n293), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT38), .B1(new_n401), .B2(KEYINPUT82), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n402), .B(new_n390), .C1(KEYINPUT82), .C2(new_n401), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n330), .A2(new_n334), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n392), .A2(new_n398), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n319), .B1(new_n388), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n262), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n407), .A2(new_n316), .A3(new_n397), .A4(new_n385), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT35), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n411), .A2(new_n397), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n263), .A2(new_n318), .A3(new_n315), .A4(new_n314), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n407), .A2(new_n316), .A3(KEYINPUT35), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OR3_X1    g217(.A1(new_n406), .A2(new_n410), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT91), .ZN(new_n420));
  AND2_X1   g219(.A1(G71gat), .A2(G78gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(KEYINPUT9), .ZN(new_n422));
  XNOR2_X1  g221(.A(G57gat), .B(G64gat), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(G71gat), .A2(G78gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  OAI221_X1 g226(.A(new_n420), .B1(new_n421), .B2(new_n425), .C1(new_n422), .C2(new_n423), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT21), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G231gat), .A2(G233gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G127gat), .B(G155gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G183gat), .B(G211gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT16), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(G1gat), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(KEYINPUT87), .C1(G1gat), .C2(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(G8gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n431), .B2(new_n430), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT92), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(KEYINPUT93), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n440), .B(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G134gat), .B(G162gat), .Z(new_n451));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n452));
  AND2_X1   g251(.A1(G43gat), .A2(G50gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(G43gat), .A2(G50gat), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT15), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G43gat), .ZN(new_n456));
  INV_X1    g255(.A(G50gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT15), .ZN(new_n459));
  NAND2_X1  g258(.A1(G43gat), .A2(G50gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G29gat), .A2(G36gat), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NOR3_X1   g264(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n452), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n463), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT14), .ZN(new_n470));
  INV_X1    g269(.A(G29gat), .ZN(new_n471));
  INV_X1    g270(.A(G36gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n469), .B1(new_n473), .B2(new_n464), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(KEYINPUT85), .A3(new_n455), .A4(new_n461), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n476));
  INV_X1    g275(.A(new_n455), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n474), .A2(KEYINPUT84), .A3(new_n455), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n468), .B(new_n475), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G99gat), .A2(G106gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT8), .ZN(new_n483));
  NAND2_X1  g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G85gat), .ZN(new_n487));
  INV_X1    g286(.A(G92gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n483), .A2(new_n486), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G99gat), .B(G106gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g293(.A1(KEYINPUT8), .A2(new_n482), .B1(new_n487), .B2(new_n488), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n495), .A2(new_n492), .A3(new_n486), .A4(new_n490), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT41), .ZN(new_n498));
  NAND2_X1  g297(.A1(G232gat), .A2(G233gat), .ZN(new_n499));
  OAI22_X1  g298(.A1(new_n481), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n480), .A2(KEYINPUT88), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT88), .B1(new_n480), .B2(new_n501), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n500), .B1(new_n509), .B2(new_n497), .ZN(new_n510));
  XOR2_X1   g309(.A(G190gat), .B(G218gat), .Z(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT94), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n499), .A2(new_n498), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n512), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n451), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n518), .ZN(new_n520));
  INV_X1    g319(.A(new_n451), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n450), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n446), .A2(new_n481), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(new_n509), .B2(new_n446), .ZN(new_n526));
  NAND2_X1  g325(.A1(G229gat), .A2(G233gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n525), .A2(KEYINPUT90), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(new_n446), .B2(new_n481), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n527), .B(KEYINPUT13), .Z(new_n534));
  AOI22_X1  g333(.A1(new_n528), .A2(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n527), .ZN(new_n536));
  AOI211_X1 g335(.A(new_n536), .B(new_n525), .C1(new_n509), .C2(new_n446), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT89), .B1(new_n537), .B2(KEYINPUT18), .ZN(new_n538));
  AND4_X1   g337(.A1(KEYINPUT89), .A2(new_n526), .A3(KEYINPUT18), .A4(new_n527), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT11), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(new_n207), .ZN(new_n543));
  INV_X1    g342(.A(G197gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n535), .B(new_n547), .C1(new_n538), .C2(new_n539), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n491), .A2(KEYINPUT95), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n495), .A2(new_n555), .A3(new_n486), .A4(new_n490), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT96), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n557), .A2(new_n493), .B1(new_n558), .B2(new_n496), .ZN(new_n559));
  AOI211_X1 g358(.A(KEYINPUT96), .B(new_n492), .C1(new_n554), .C2(new_n556), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n429), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n429), .A2(new_n497), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT10), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n497), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(new_n429), .A3(KEYINPUT10), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n553), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n557), .A2(new_n558), .A3(new_n493), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n492), .B1(new_n554), .B2(new_n556), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n496), .A2(new_n558), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n562), .B1(new_n573), .B2(new_n429), .ZN(new_n574));
  INV_X1    g373(.A(new_n553), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(G176gat), .B(G204gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  OR3_X1    g378(.A1(new_n569), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n569), .B2(new_n576), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n552), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n524), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n419), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n398), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g387(.A1(new_n419), .A2(new_n343), .A3(new_n585), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(new_n445), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT97), .ZN(new_n591));
  XOR2_X1   g390(.A(KEYINPUT16), .B(G8gat), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT42), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(G1325gat));
  INV_X1    g394(.A(G15gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n586), .A2(new_n596), .A3(new_n407), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n263), .A2(new_n318), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n586), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n597), .B1(new_n600), .B2(new_n596), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(G1326gat));
  INV_X1    g402(.A(new_n316), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n605), .A2(KEYINPUT99), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(KEYINPUT99), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT43), .B(G22gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(G1327gat));
  INV_X1    g412(.A(KEYINPUT45), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n406), .A2(new_n410), .A3(new_n418), .ZN(new_n615));
  INV_X1    g414(.A(new_n523), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n450), .A2(new_n584), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n397), .A2(G29gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n614), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(KEYINPUT45), .A3(new_n621), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT44), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n615), .B2(new_n616), .ZN(new_n628));
  INV_X1    g427(.A(new_n617), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n408), .A2(new_n409), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n416), .A2(new_n417), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n630), .B1(new_n631), .B2(new_n415), .ZN(new_n632));
  OAI211_X1 g431(.A(KEYINPUT44), .B(new_n523), .C1(new_n632), .C2(new_n406), .ZN(new_n633));
  AND4_X1   g432(.A1(new_n398), .A2(new_n628), .A3(new_n629), .A4(new_n633), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n624), .B(new_n626), .C1(new_n471), .C2(new_n634), .ZN(G1328gat));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n615), .A2(new_n616), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n385), .A2(G36gat), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n629), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n618), .A2(KEYINPUT101), .A3(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n636), .B1(new_n643), .B2(KEYINPUT46), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT46), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n641), .A2(KEYINPUT102), .A3(new_n645), .A4(new_n642), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n628), .A2(new_n633), .A3(new_n343), .A4(new_n629), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n643), .A2(KEYINPUT46), .B1(G36gat), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(G1329gat));
  NAND4_X1  g449(.A1(new_n628), .A2(new_n633), .A3(new_n599), .A4(new_n629), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(G43gat), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT47), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n618), .A2(new_n456), .A3(new_n407), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n654), .B(new_n656), .ZN(G1330gat));
  NAND4_X1  g456(.A1(new_n628), .A2(new_n633), .A3(new_n604), .A4(new_n629), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n316), .A2(G50gat), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n658), .A2(G50gat), .B1(new_n618), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT105), .B(KEYINPUT48), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OR3_X1    g462(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n663), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(G1331gat));
  NAND3_X1  g465(.A1(new_n524), .A2(new_n552), .A3(new_n583), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT106), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n419), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n397), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT107), .B(G57gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1332gat));
  INV_X1    g471(.A(new_n669), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n385), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(G1333gat));
  NAND3_X1  g476(.A1(new_n673), .A2(G71gat), .A3(new_n599), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n262), .B(KEYINPUT108), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n669), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(G71gat), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g481(.A1(new_n673), .A2(new_n604), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g483(.A1(new_n450), .A2(new_n552), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT51), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(KEYINPUT110), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT51), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n637), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n523), .B(new_n687), .C1(new_n632), .C2(new_n406), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(new_n688), .A3(KEYINPUT51), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n397), .A2(G85gat), .A3(new_n582), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n685), .A2(new_n582), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n628), .A2(new_n633), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT109), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n628), .A2(new_n633), .A3(new_n698), .A4(new_n695), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n697), .A2(new_n398), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n694), .B1(new_n700), .B2(new_n487), .ZN(G1336gat));
  NOR3_X1   g500(.A1(new_n385), .A2(G92gat), .A3(new_n582), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n690), .A2(new_n692), .A3(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n628), .A2(new_n633), .A3(new_n343), .A4(new_n695), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT52), .B1(new_n704), .B2(G92gat), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n703), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  AND4_X1   g508(.A1(new_n706), .A2(new_n690), .A3(new_n692), .A4(new_n702), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n697), .A2(new_n343), .A3(new_n699), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(G92gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n712), .B2(new_n707), .ZN(G1337gat));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n599), .A3(new_n699), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT112), .B(G99gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n262), .A2(new_n582), .A3(new_n715), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n690), .A2(new_n692), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(G1338gat));
  NOR3_X1   g518(.A1(new_n316), .A2(G106gat), .A3(new_n582), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n690), .A2(new_n692), .A3(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n628), .A2(new_n633), .A3(new_n604), .A4(new_n695), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT53), .B1(new_n722), .B2(G106gat), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n721), .B1(new_n723), .B2(new_n726), .ZN(new_n727));
  AND4_X1   g526(.A1(new_n724), .A2(new_n690), .A3(new_n692), .A4(new_n720), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n697), .A2(new_n604), .A3(new_n699), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(G106gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n730), .B2(new_n725), .ZN(G1339gat));
  OAI211_X1 g530(.A(new_n566), .B(new_n575), .C1(new_n574), .C2(KEYINPUT10), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n568), .A2(KEYINPUT54), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT114), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n568), .A2(new_n732), .A3(new_n735), .A4(KEYINPUT54), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n737), .B(new_n553), .C1(new_n564), .C2(new_n567), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n738), .A2(new_n739), .A3(new_n579), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n738), .B2(new_n579), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n734), .B(new_n736), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n580), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT116), .B(new_n580), .C1(new_n742), .C2(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n742), .A2(new_n743), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n551), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  OAI22_X1  g548(.A1(new_n526), .A2(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n750));
  INV_X1    g549(.A(new_n545), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n550), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n583), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n616), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n523), .A2(new_n753), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(KEYINPUT117), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT117), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n523), .B1(new_n749), .B2(new_n754), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n757), .A2(new_n758), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n450), .A3(new_n764), .ZN(new_n765));
  NOR4_X1   g564(.A1(new_n450), .A2(new_n523), .A3(new_n551), .A4(new_n583), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n397), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n604), .A2(new_n262), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n385), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n552), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT118), .B(G113gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1340gat));
  NOR2_X1   g573(.A1(new_n771), .A2(new_n582), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g575(.A1(new_n771), .A2(new_n450), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n233), .ZN(G1342gat));
  NOR2_X1   g577(.A1(new_n343), .A2(new_n616), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n770), .A2(new_n234), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT56), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n780), .A2(new_n781), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n779), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G134gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n783), .A2(new_n787), .A3(new_n789), .ZN(G1343gat));
  INV_X1    g589(.A(new_n450), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n551), .A2(new_n748), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n754), .B1(new_n792), .B2(new_n744), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n616), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n794), .B2(new_n759), .ZN(new_n795));
  OAI211_X1 g594(.A(KEYINPUT57), .B(new_n604), .C1(new_n795), .C2(new_n766), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n316), .B1(new_n765), .B2(new_n767), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(KEYINPUT57), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n598), .A2(new_n398), .A3(new_n385), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G141gat), .B1(new_n801), .B2(new_n552), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803));
  INV_X1    g602(.A(new_n416), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n768), .A2(KEYINPUT121), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n806));
  AOI211_X1 g605(.A(new_n806), .B(new_n397), .C1(new_n765), .C2(new_n767), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n385), .B(new_n804), .C1(new_n805), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n552), .A2(G141gat), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n802), .B(new_n803), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n808), .A2(new_n810), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n801), .A2(KEYINPUT120), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n814), .A3(new_n800), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n551), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n812), .B1(new_n816), .B2(G141gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n811), .B1(new_n817), .B2(new_n803), .ZN(G1344gat));
  OR3_X1    g617(.A1(new_n808), .A2(G148gat), .A3(new_n582), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(new_n604), .C1(new_n795), .C2(new_n766), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n583), .B(new_n821), .C1(new_n797), .C2(new_n820), .ZN(new_n822));
  OAI21_X1  g621(.A(G148gat), .B1(new_n822), .B2(new_n799), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT59), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(KEYINPUT122), .A3(KEYINPUT59), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(G148gat), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n798), .A2(new_n814), .A3(new_n800), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n814), .B1(new_n798), .B2(new_n800), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n833), .B2(new_n583), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n819), .B1(new_n828), .B2(new_n834), .ZN(G1345gat));
  NOR2_X1   g634(.A1(new_n808), .A2(new_n450), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n836), .A2(KEYINPUT123), .ZN(new_n837));
  AOI21_X1  g636(.A(G155gat), .B1(new_n836), .B2(KEYINPUT123), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n450), .A2(new_n269), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n837), .A2(new_n838), .B1(new_n833), .B2(new_n839), .ZN(G1346gat));
  NOR3_X1   g639(.A1(new_n343), .A2(new_n616), .A3(G162gat), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n804), .B(new_n841), .C1(new_n805), .C2(new_n807), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT124), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n831), .A2(new_n832), .A3(new_n616), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n270), .B2(new_n844), .ZN(G1347gat));
  AOI211_X1 g644(.A(new_n398), .B(new_n385), .C1(new_n765), .C2(new_n767), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n846), .A2(new_n769), .ZN(new_n847));
  AOI21_X1  g646(.A(G169gat), .B1(new_n847), .B2(new_n551), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n679), .A2(new_n604), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(new_n207), .A3(new_n552), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n848), .A2(new_n851), .ZN(G1348gat));
  NAND3_X1  g651(.A1(new_n847), .A2(new_n208), .A3(new_n583), .ZN(new_n853));
  OAI21_X1  g652(.A(G176gat), .B1(new_n850), .B2(new_n582), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1349gat));
  NAND3_X1  g654(.A1(new_n847), .A2(new_n221), .A3(new_n791), .ZN(new_n856));
  OAI21_X1  g655(.A(G183gat), .B1(new_n850), .B2(new_n450), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g659(.A(G190gat), .B1(new_n850), .B2(new_n616), .ZN(new_n861));
  XNOR2_X1  g660(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n222), .A3(new_n523), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G1351gat));
  NAND2_X1  g665(.A1(new_n846), .A2(new_n804), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n544), .B1(new_n867), .B2(new_n552), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n398), .A2(new_n385), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n598), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n821), .B(new_n871), .C1(new_n797), .C2(new_n820), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n551), .A2(G197gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n868), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(G1352gat));
  OAI21_X1  g674(.A(G204gat), .B1(new_n822), .B2(new_n870), .ZN(new_n876));
  OR3_X1    g675(.A1(new_n867), .A2(G204gat), .A3(new_n582), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT62), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n877), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT127), .B1(new_n877), .B2(KEYINPUT62), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n876), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(G1353gat));
  OR2_X1    g680(.A1(new_n872), .A2(new_n450), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT63), .B1(new_n882), .B2(G211gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n791), .A2(new_n282), .ZN(new_n886));
  OAI22_X1  g685(.A1(new_n884), .A2(new_n885), .B1(new_n867), .B2(new_n886), .ZN(G1354gat));
  NOR2_X1   g686(.A1(new_n867), .A2(new_n616), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n616), .A2(new_n281), .ZN(new_n889));
  OAI22_X1  g688(.A1(new_n888), .A2(G218gat), .B1(new_n872), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(G1355gat));
endmodule


