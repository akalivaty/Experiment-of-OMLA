

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n680), .A2(n679), .ZN(n687) );
  AND2_X1 U550 ( .A1(n723), .A2(n722), .ZN(n513) );
  NOR2_X1 U551 ( .A1(n684), .A2(G1966), .ZN(n581) );
  NAND2_X1 U552 ( .A1(G8), .A2(n627), .ZN(n684) );
  NOR2_X1 U553 ( .A1(n721), .A2(n727), .ZN(n722) );
  NOR2_X1 U554 ( .A1(G2104), .A2(G2105), .ZN(n514) );
  XOR2_X1 U555 ( .A(KEYINPUT64), .B(n514), .Z(n515) );
  NOR2_X1 U556 ( .A1(n553), .A2(G651), .ZN(n779) );
  XNOR2_X2 U557 ( .A(KEYINPUT17), .B(n515), .ZN(n877) );
  NAND2_X1 U558 ( .A1(G138), .A2(n877), .ZN(n518) );
  INV_X1 U559 ( .A(G2105), .ZN(n519) );
  AND2_X1 U560 ( .A1(n519), .A2(G2104), .ZN(n869) );
  NAND2_X1 U561 ( .A1(G102), .A2(n869), .ZN(n516) );
  XOR2_X1 U562 ( .A(KEYINPUT85), .B(n516), .Z(n517) );
  NAND2_X1 U563 ( .A1(n518), .A2(n517), .ZN(n523) );
  NOR2_X1 U564 ( .A1(G2104), .A2(n519), .ZN(n871) );
  NAND2_X1 U565 ( .A1(G126), .A2(n871), .ZN(n521) );
  AND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n872) );
  NAND2_X1 U567 ( .A1(G114), .A2(n872), .ZN(n520) );
  NAND2_X1 U568 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U569 ( .A1(n523), .A2(n522), .ZN(G164) );
  NOR2_X1 U570 ( .A1(G543), .A2(G651), .ZN(n775) );
  NAND2_X1 U571 ( .A1(n775), .A2(G89), .ZN(n524) );
  XNOR2_X1 U572 ( .A(n524), .B(KEYINPUT4), .ZN(n526) );
  XOR2_X1 U573 ( .A(KEYINPUT0), .B(G543), .Z(n553) );
  XNOR2_X1 U574 ( .A(KEYINPUT67), .B(G651), .ZN(n528) );
  NOR2_X1 U575 ( .A1(n553), .A2(n528), .ZN(n776) );
  NAND2_X1 U576 ( .A1(G76), .A2(n776), .ZN(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U578 ( .A(KEYINPUT5), .B(n527), .ZN(n535) );
  NAND2_X1 U579 ( .A1(n779), .A2(G51), .ZN(n531) );
  NOR2_X1 U580 ( .A1(G543), .A2(n528), .ZN(n529) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n529), .Z(n783) );
  NAND2_X1 U582 ( .A1(G63), .A2(n783), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n533) );
  XOR2_X1 U584 ( .A(KEYINPUT72), .B(KEYINPUT6), .Z(n532) );
  XNOR2_X1 U585 ( .A(n533), .B(n532), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U587 ( .A(KEYINPUT7), .B(n536), .ZN(G168) );
  NAND2_X1 U588 ( .A1(n779), .A2(G52), .ZN(n538) );
  NAND2_X1 U589 ( .A1(G64), .A2(n783), .ZN(n537) );
  NAND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n544) );
  NAND2_X1 U591 ( .A1(n775), .A2(G90), .ZN(n539) );
  XNOR2_X1 U592 ( .A(n539), .B(KEYINPUT68), .ZN(n541) );
  NAND2_X1 U593 ( .A1(G77), .A2(n776), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U595 ( .A(KEYINPUT9), .B(n542), .Z(n543) );
  NOR2_X1 U596 ( .A1(n544), .A2(n543), .ZN(G171) );
  XNOR2_X1 U597 ( .A(G168), .B(KEYINPUT8), .ZN(n545) );
  XNOR2_X1 U598 ( .A(n545), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U599 ( .A1(n775), .A2(G88), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G75), .A2(n776), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n779), .A2(G50), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G62), .A2(n783), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(G166) );
  XOR2_X1 U606 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NAND2_X1 U607 ( .A1(G49), .A2(n779), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT78), .ZN(n558) );
  NAND2_X1 U609 ( .A1(G74), .A2(G651), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G87), .A2(n553), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n783), .A2(n556), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n558), .A2(n557), .ZN(G288) );
  NAND2_X1 U614 ( .A1(n775), .A2(G86), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G61), .A2(n783), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n776), .A2(G73), .ZN(n561) );
  XOR2_X1 U618 ( .A(KEYINPUT2), .B(n561), .Z(n562) );
  NOR2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U620 ( .A1(n779), .A2(G48), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n565), .A2(n564), .ZN(G305) );
  NAND2_X1 U622 ( .A1(G72), .A2(n776), .ZN(n567) );
  NAND2_X1 U623 ( .A1(G60), .A2(n783), .ZN(n566) );
  NAND2_X1 U624 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n775), .A2(G85), .ZN(n568) );
  XOR2_X1 U626 ( .A(KEYINPUT66), .B(n568), .Z(n569) );
  NOR2_X1 U627 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U628 ( .A1(n779), .A2(G47), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(G290) );
  NOR2_X1 U630 ( .A1(G164), .A2(G1384), .ZN(n690) );
  NAND2_X1 U631 ( .A1(G101), .A2(n869), .ZN(n573) );
  XOR2_X1 U632 ( .A(KEYINPUT23), .B(n573), .Z(n576) );
  NAND2_X1 U633 ( .A1(n877), .A2(G137), .ZN(n574) );
  XOR2_X1 U634 ( .A(n574), .B(KEYINPUT65), .Z(n575) );
  NAND2_X1 U635 ( .A1(n576), .A2(n575), .ZN(n750) );
  NAND2_X1 U636 ( .A1(G125), .A2(n871), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G113), .A2(n872), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n749) );
  INV_X1 U639 ( .A(G40), .ZN(n579) );
  OR2_X1 U640 ( .A1(n749), .A2(n579), .ZN(n580) );
  NOR2_X1 U641 ( .A1(n750), .A2(n580), .ZN(n688) );
  NAND2_X1 U642 ( .A1(n690), .A2(n688), .ZN(n627) );
  INV_X1 U643 ( .A(n627), .ZN(n628) );
  INV_X1 U644 ( .A(n628), .ZN(n645) );
  NOR2_X1 U645 ( .A1(G2084), .A2(n645), .ZN(n653) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT92), .ZN(n655) );
  NOR2_X1 U647 ( .A1(n653), .A2(n655), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT94), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n583), .A2(G8), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n584), .B(KEYINPUT30), .ZN(n585) );
  NOR2_X1 U651 ( .A1(n585), .A2(G168), .ZN(n590) );
  XOR2_X1 U652 ( .A(G2078), .B(KEYINPUT93), .Z(n586) );
  XNOR2_X1 U653 ( .A(KEYINPUT25), .B(n586), .ZN(n911) );
  NOR2_X1 U654 ( .A1(n645), .A2(n911), .ZN(n588) );
  AND2_X1 U655 ( .A1(n645), .A2(G1961), .ZN(n587) );
  NOR2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n593) );
  NOR2_X1 U657 ( .A1(G171), .A2(n593), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U659 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n592), .B(n591), .ZN(n644) );
  NAND2_X1 U661 ( .A1(G171), .A2(n593), .ZN(n642) );
  NAND2_X1 U662 ( .A1(n775), .A2(G91), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G78), .A2(n776), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n779), .A2(G53), .ZN(n597) );
  NAND2_X1 U666 ( .A1(G65), .A2(n783), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U669 ( .A(KEYINPUT69), .B(n600), .Z(n928) );
  NAND2_X1 U670 ( .A1(n628), .A2(G2072), .ZN(n601) );
  XNOR2_X1 U671 ( .A(n601), .B(KEYINPUT27), .ZN(n603) );
  INV_X1 U672 ( .A(G1956), .ZN(n949) );
  NOR2_X1 U673 ( .A1(n949), .A2(n628), .ZN(n602) );
  NOR2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n605) );
  NOR2_X1 U675 ( .A1(n928), .A2(n605), .ZN(n604) );
  XOR2_X1 U676 ( .A(n604), .B(KEYINPUT28), .Z(n639) );
  NAND2_X1 U677 ( .A1(n928), .A2(n605), .ZN(n637) );
  NAND2_X1 U678 ( .A1(n775), .A2(G81), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT12), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G68), .A2(n776), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U682 ( .A(KEYINPUT13), .B(n609), .ZN(n615) );
  NAND2_X1 U683 ( .A1(n783), .A2(G56), .ZN(n610) );
  XOR2_X1 U684 ( .A(KEYINPUT14), .B(n610), .Z(n613) );
  NAND2_X1 U685 ( .A1(G43), .A2(n779), .ZN(n611) );
  XNOR2_X1 U686 ( .A(KEYINPUT71), .B(n611), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n941) );
  AND2_X1 U689 ( .A1(n628), .A2(G1996), .ZN(n616) );
  XOR2_X1 U690 ( .A(n616), .B(KEYINPUT26), .Z(n618) );
  NAND2_X1 U691 ( .A1(n627), .A2(G1341), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U693 ( .A1(n941), .A2(n619), .ZN(n632) );
  NAND2_X1 U694 ( .A1(n779), .A2(G54), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G66), .A2(n783), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n775), .A2(G92), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G79), .A2(n776), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(KEYINPUT15), .ZN(n924) );
  NAND2_X1 U702 ( .A1(G1348), .A2(n627), .ZN(n630) );
  NAND2_X1 U703 ( .A1(G2067), .A2(n628), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n633) );
  NOR2_X1 U705 ( .A1(n924), .A2(n633), .ZN(n631) );
  OR2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n924), .A2(n633), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U711 ( .A(KEYINPUT29), .B(n640), .Z(n641) );
  NAND2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n654) );
  NAND2_X1 U714 ( .A1(n654), .A2(G286), .ZN(n650) );
  NOR2_X1 U715 ( .A1(G1971), .A2(n684), .ZN(n647) );
  NOR2_X1 U716 ( .A1(G2090), .A2(n645), .ZN(n646) );
  NOR2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U718 ( .A1(G303), .A2(n648), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U720 ( .A1(n651), .A2(G8), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n652), .B(KEYINPUT32), .ZN(n660) );
  NAND2_X1 U722 ( .A1(G8), .A2(n653), .ZN(n658) );
  INV_X1 U723 ( .A(n654), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n683) );
  NOR2_X1 U727 ( .A1(G1976), .A2(G288), .ZN(n668) );
  NOR2_X1 U728 ( .A1(G303), .A2(G1971), .ZN(n661) );
  NOR2_X1 U729 ( .A1(n668), .A2(n661), .ZN(n935) );
  NAND2_X1 U730 ( .A1(n683), .A2(n935), .ZN(n663) );
  NAND2_X1 U731 ( .A1(G288), .A2(G1976), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n662), .B(KEYINPUT96), .ZN(n931) );
  NAND2_X1 U733 ( .A1(n663), .A2(n931), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT97), .ZN(n665) );
  INV_X1 U735 ( .A(n684), .ZN(n669) );
  NAND2_X1 U736 ( .A1(n665), .A2(n669), .ZN(n666) );
  INV_X1 U737 ( .A(KEYINPUT33), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n666), .A2(n671), .ZN(n676) );
  OR2_X1 U739 ( .A1(G1981), .A2(G305), .ZN(n677) );
  NAND2_X1 U740 ( .A1(G1981), .A2(G305), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n677), .A2(n667), .ZN(n921) );
  INV_X1 U742 ( .A(n921), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U744 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U745 ( .A(n672), .B(KEYINPUT98), .Z(n673) );
  AND2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n675) );
  AND2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n680) );
  XNOR2_X1 U748 ( .A(n677), .B(KEYINPUT24), .ZN(n678) );
  NOR2_X1 U749 ( .A1(n684), .A2(n678), .ZN(n679) );
  NOR2_X1 U750 ( .A1(G2090), .A2(G303), .ZN(n681) );
  NAND2_X1 U751 ( .A1(G8), .A2(n681), .ZN(n682) );
  NAND2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n723) );
  INV_X1 U755 ( .A(n688), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n690), .A2(n689), .ZN(n734) );
  NAND2_X1 U757 ( .A1(G140), .A2(n877), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n869), .A2(G104), .ZN(n691) );
  XOR2_X1 U759 ( .A(KEYINPUT87), .B(n691), .Z(n692) );
  NAND2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n696) );
  XOR2_X1 U761 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n694) );
  XNOR2_X1 U762 ( .A(KEYINPUT34), .B(n694), .ZN(n695) );
  XNOR2_X1 U763 ( .A(n696), .B(n695), .ZN(n702) );
  NAND2_X1 U764 ( .A1(G128), .A2(n871), .ZN(n698) );
  NAND2_X1 U765 ( .A1(G116), .A2(n872), .ZN(n697) );
  NAND2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U767 ( .A(KEYINPUT90), .B(n699), .Z(n700) );
  XNOR2_X1 U768 ( .A(KEYINPUT35), .B(n700), .ZN(n701) );
  NOR2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U770 ( .A(KEYINPUT36), .B(n703), .ZN(n888) );
  XNOR2_X1 U771 ( .A(G2067), .B(KEYINPUT37), .ZN(n732) );
  NOR2_X1 U772 ( .A1(n888), .A2(n732), .ZN(n1000) );
  NAND2_X1 U773 ( .A1(n734), .A2(n1000), .ZN(n704) );
  XOR2_X1 U774 ( .A(KEYINPUT91), .B(n704), .Z(n730) );
  INV_X1 U775 ( .A(n730), .ZN(n721) );
  NAND2_X1 U776 ( .A1(G95), .A2(n869), .ZN(n706) );
  NAND2_X1 U777 ( .A1(G131), .A2(n877), .ZN(n705) );
  NAND2_X1 U778 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U779 ( .A1(G119), .A2(n871), .ZN(n708) );
  NAND2_X1 U780 ( .A1(G107), .A2(n872), .ZN(n707) );
  NAND2_X1 U781 ( .A1(n708), .A2(n707), .ZN(n709) );
  OR2_X1 U782 ( .A1(n710), .A2(n709), .ZN(n864) );
  AND2_X1 U783 ( .A1(n864), .A2(G1991), .ZN(n719) );
  NAND2_X1 U784 ( .A1(G129), .A2(n871), .ZN(n712) );
  NAND2_X1 U785 ( .A1(G117), .A2(n872), .ZN(n711) );
  NAND2_X1 U786 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U787 ( .A1(n869), .A2(G105), .ZN(n713) );
  XOR2_X1 U788 ( .A(KEYINPUT38), .B(n713), .Z(n714) );
  NOR2_X1 U789 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U790 ( .A1(G141), .A2(n877), .ZN(n716) );
  NAND2_X1 U791 ( .A1(n717), .A2(n716), .ZN(n885) );
  AND2_X1 U792 ( .A1(G1996), .A2(n885), .ZN(n718) );
  NOR2_X1 U793 ( .A1(n719), .A2(n718), .ZN(n985) );
  INV_X1 U794 ( .A(n734), .ZN(n720) );
  NOR2_X1 U795 ( .A1(n985), .A2(n720), .ZN(n727) );
  XNOR2_X1 U796 ( .A(G1986), .B(G290), .ZN(n932) );
  NAND2_X1 U797 ( .A1(n932), .A2(n734), .ZN(n724) );
  NAND2_X1 U798 ( .A1(n513), .A2(n724), .ZN(n737) );
  NOR2_X1 U799 ( .A1(G1996), .A2(n885), .ZN(n980) );
  NOR2_X1 U800 ( .A1(G1986), .A2(G290), .ZN(n725) );
  NOR2_X1 U801 ( .A1(G1991), .A2(n864), .ZN(n983) );
  NOR2_X1 U802 ( .A1(n725), .A2(n983), .ZN(n726) );
  NOR2_X1 U803 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U804 ( .A1(n980), .A2(n728), .ZN(n729) );
  XNOR2_X1 U805 ( .A(n729), .B(KEYINPUT39), .ZN(n731) );
  NAND2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n733) );
  NAND2_X1 U807 ( .A1(n888), .A2(n732), .ZN(n989) );
  NAND2_X1 U808 ( .A1(n733), .A2(n989), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U810 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U811 ( .A(n738), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U812 ( .A(G2430), .B(G2451), .Z(n740) );
  XNOR2_X1 U813 ( .A(KEYINPUT99), .B(G2443), .ZN(n739) );
  XNOR2_X1 U814 ( .A(n740), .B(n739), .ZN(n747) );
  XOR2_X1 U815 ( .A(G2435), .B(G2446), .Z(n742) );
  XNOR2_X1 U816 ( .A(G2427), .B(G2454), .ZN(n741) );
  XNOR2_X1 U817 ( .A(n742), .B(n741), .ZN(n743) );
  XOR2_X1 U818 ( .A(n743), .B(G2438), .Z(n745) );
  XNOR2_X1 U819 ( .A(G1341), .B(G1348), .ZN(n744) );
  XNOR2_X1 U820 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U821 ( .A(n747), .B(n746), .ZN(n748) );
  AND2_X1 U822 ( .A1(n748), .A2(G14), .ZN(G401) );
  INV_X1 U823 ( .A(G171), .ZN(G301) );
  AND2_X1 U824 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U825 ( .A(G57), .ZN(G237) );
  INV_X1 U826 ( .A(G120), .ZN(G236) );
  NOR2_X1 U827 ( .A1(n750), .A2(n749), .ZN(G160) );
  NAND2_X1 U828 ( .A1(G7), .A2(G661), .ZN(n751) );
  XNOR2_X1 U829 ( .A(n751), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U830 ( .A(G223), .ZN(n819) );
  NAND2_X1 U831 ( .A1(n819), .A2(G567), .ZN(n752) );
  XOR2_X1 U832 ( .A(KEYINPUT11), .B(n752), .Z(G234) );
  INV_X1 U833 ( .A(G860), .ZN(n757) );
  OR2_X1 U834 ( .A1(n941), .A2(n757), .ZN(G153) );
  NAND2_X1 U835 ( .A1(G868), .A2(G301), .ZN(n754) );
  INV_X1 U836 ( .A(G868), .ZN(n798) );
  NAND2_X1 U837 ( .A1(n924), .A2(n798), .ZN(n753) );
  NAND2_X1 U838 ( .A1(n754), .A2(n753), .ZN(G284) );
  XOR2_X1 U839 ( .A(n928), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U840 ( .A1(G868), .A2(G299), .ZN(n756) );
  NOR2_X1 U841 ( .A1(G286), .A2(n798), .ZN(n755) );
  NOR2_X1 U842 ( .A1(n756), .A2(n755), .ZN(G297) );
  NAND2_X1 U843 ( .A1(G559), .A2(n757), .ZN(n758) );
  XNOR2_X1 U844 ( .A(KEYINPUT74), .B(n758), .ZN(n759) );
  INV_X1 U845 ( .A(n924), .ZN(n786) );
  NAND2_X1 U846 ( .A1(n759), .A2(n786), .ZN(n760) );
  XNOR2_X1 U847 ( .A(KEYINPUT16), .B(n760), .ZN(G148) );
  NOR2_X1 U848 ( .A1(G868), .A2(n941), .ZN(n763) );
  NAND2_X1 U849 ( .A1(G868), .A2(n786), .ZN(n761) );
  NOR2_X1 U850 ( .A1(G559), .A2(n761), .ZN(n762) );
  NOR2_X1 U851 ( .A1(n763), .A2(n762), .ZN(G282) );
  NAND2_X1 U852 ( .A1(G111), .A2(n872), .ZN(n764) );
  XNOR2_X1 U853 ( .A(n764), .B(KEYINPUT76), .ZN(n768) );
  XOR2_X1 U854 ( .A(KEYINPUT75), .B(KEYINPUT18), .Z(n766) );
  NAND2_X1 U855 ( .A1(G123), .A2(n871), .ZN(n765) );
  XNOR2_X1 U856 ( .A(n766), .B(n765), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n772) );
  NAND2_X1 U858 ( .A1(G99), .A2(n869), .ZN(n770) );
  NAND2_X1 U859 ( .A1(G135), .A2(n877), .ZN(n769) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n982) );
  XNOR2_X1 U862 ( .A(n982), .B(G2096), .ZN(n774) );
  INV_X1 U863 ( .A(G2100), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(G156) );
  NAND2_X1 U865 ( .A1(n775), .A2(G93), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G80), .A2(n776), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G55), .A2(n779), .ZN(n780) );
  XNOR2_X1 U869 ( .A(KEYINPUT77), .B(n780), .ZN(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G67), .A2(n783), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n799) );
  NAND2_X1 U873 ( .A1(n786), .A2(G559), .ZN(n796) );
  XNOR2_X1 U874 ( .A(n941), .B(n796), .ZN(n787) );
  NOR2_X1 U875 ( .A1(G860), .A2(n787), .ZN(n788) );
  XOR2_X1 U876 ( .A(n799), .B(n788), .Z(G145) );
  XNOR2_X1 U877 ( .A(G305), .B(n799), .ZN(n793) );
  XNOR2_X1 U878 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n790) );
  XNOR2_X1 U879 ( .A(G290), .B(G166), .ZN(n789) );
  XNOR2_X1 U880 ( .A(n790), .B(n789), .ZN(n791) );
  XNOR2_X1 U881 ( .A(n791), .B(G288), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n793), .B(n792), .ZN(n794) );
  XNOR2_X1 U883 ( .A(G299), .B(n794), .ZN(n795) );
  XNOR2_X1 U884 ( .A(n795), .B(n941), .ZN(n891) );
  XOR2_X1 U885 ( .A(n891), .B(n796), .Z(n797) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n801) );
  NOR2_X1 U887 ( .A1(G868), .A2(n799), .ZN(n800) );
  NOR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(G295) );
  XOR2_X1 U889 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n803) );
  NAND2_X1 U890 ( .A1(G2084), .A2(G2078), .ZN(n802) );
  XNOR2_X1 U891 ( .A(n803), .B(n802), .ZN(n804) );
  NAND2_X1 U892 ( .A1(G2090), .A2(n804), .ZN(n805) );
  XNOR2_X1 U893 ( .A(KEYINPUT21), .B(n805), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n806), .A2(G2072), .ZN(G158) );
  XOR2_X1 U895 ( .A(KEYINPUT81), .B(G44), .Z(n807) );
  XNOR2_X1 U896 ( .A(KEYINPUT3), .B(n807), .ZN(G218) );
  NOR2_X1 U897 ( .A1(G236), .A2(G237), .ZN(n808) );
  NAND2_X1 U898 ( .A1(G69), .A2(n808), .ZN(n809) );
  XNOR2_X1 U899 ( .A(KEYINPUT83), .B(n809), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n810), .A2(G108), .ZN(n823) );
  NAND2_X1 U901 ( .A1(G567), .A2(n823), .ZN(n811) );
  XNOR2_X1 U902 ( .A(n811), .B(KEYINPUT84), .ZN(n817) );
  NAND2_X1 U903 ( .A1(G132), .A2(G82), .ZN(n812) );
  XNOR2_X1 U904 ( .A(n812), .B(KEYINPUT22), .ZN(n813) );
  XNOR2_X1 U905 ( .A(n813), .B(KEYINPUT82), .ZN(n814) );
  NOR2_X1 U906 ( .A1(G218), .A2(n814), .ZN(n815) );
  NAND2_X1 U907 ( .A1(G96), .A2(n815), .ZN(n824) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n824), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n895) );
  NAND2_X1 U910 ( .A1(G661), .A2(G483), .ZN(n818) );
  NOR2_X1 U911 ( .A1(n895), .A2(n818), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n822), .A2(G36), .ZN(G176) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U915 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(G188) );
  XOR2_X1 U918 ( .A(G96), .B(KEYINPUT100), .Z(G221) );
  NOR2_X1 U919 ( .A1(n824), .A2(n823), .ZN(G325) );
  XNOR2_X1 U920 ( .A(KEYINPUT101), .B(G325), .ZN(G261) );
  INV_X1 U922 ( .A(G132), .ZN(G219) );
  INV_X1 U923 ( .A(G108), .ZN(G238) );
  INV_X1 U924 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U925 ( .A(G2067), .B(G2072), .ZN(n825) );
  XNOR2_X1 U926 ( .A(n825), .B(KEYINPUT42), .ZN(n835) );
  XOR2_X1 U927 ( .A(KEYINPUT103), .B(G2100), .Z(n827) );
  XNOR2_X1 U928 ( .A(G2678), .B(KEYINPUT104), .ZN(n826) );
  XNOR2_X1 U929 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U930 ( .A(G2096), .B(G2090), .Z(n829) );
  XNOR2_X1 U931 ( .A(G2078), .B(G2084), .ZN(n828) );
  XNOR2_X1 U932 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U933 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U934 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(G227) );
  XOR2_X1 U937 ( .A(G1976), .B(G1981), .Z(n837) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1971), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n847) );
  XOR2_X1 U940 ( .A(KEYINPUT106), .B(KEYINPUT41), .Z(n839) );
  XNOR2_X1 U941 ( .A(G1991), .B(KEYINPUT107), .ZN(n838) );
  XNOR2_X1 U942 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U943 ( .A(G1956), .B(G1961), .Z(n841) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1986), .ZN(n840) );
  XNOR2_X1 U945 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U946 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U947 ( .A(KEYINPUT108), .B(G2474), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G112), .A2(n872), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G100), .A2(n869), .ZN(n849) );
  NAND2_X1 U952 ( .A1(G136), .A2(n877), .ZN(n848) );
  NAND2_X1 U953 ( .A1(n849), .A2(n848), .ZN(n852) );
  NAND2_X1 U954 ( .A1(n871), .A2(G124), .ZN(n850) );
  XOR2_X1 U955 ( .A(KEYINPUT44), .B(n850), .Z(n851) );
  NOR2_X1 U956 ( .A1(n852), .A2(n851), .ZN(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n855), .B(KEYINPUT109), .ZN(G162) );
  NAND2_X1 U959 ( .A1(G130), .A2(n871), .ZN(n857) );
  NAND2_X1 U960 ( .A1(G118), .A2(n872), .ZN(n856) );
  NAND2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n863) );
  NAND2_X1 U962 ( .A1(n869), .A2(G106), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n858), .B(KEYINPUT110), .ZN(n860) );
  NAND2_X1 U964 ( .A1(G142), .A2(n877), .ZN(n859) );
  NAND2_X1 U965 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U966 ( .A(KEYINPUT45), .B(n861), .Z(n862) );
  NOR2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n868) );
  XOR2_X1 U968 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n866) );
  XOR2_X1 U969 ( .A(G160), .B(n864), .Z(n865) );
  XNOR2_X1 U970 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(n868), .B(n867), .Z(n883) );
  NAND2_X1 U972 ( .A1(n869), .A2(G103), .ZN(n870) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n870), .ZN(n881) );
  NAND2_X1 U974 ( .A1(G127), .A2(n871), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G115), .A2(n872), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n875), .B(KEYINPUT112), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT47), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G139), .A2(n877), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n991) );
  XNOR2_X1 U982 ( .A(n991), .B(n982), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(n884), .B(G162), .Z(n887) );
  XOR2_X1 U985 ( .A(G164), .B(n885), .Z(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n889) );
  XOR2_X1 U987 ( .A(n889), .B(n888), .Z(n890) );
  NOR2_X1 U988 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U989 ( .A(G286), .B(n924), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n893), .B(G301), .ZN(n894) );
  NOR2_X1 U992 ( .A1(G37), .A2(n894), .ZN(G397) );
  XOR2_X1 U993 ( .A(KEYINPUT102), .B(n895), .Z(G319) );
  NOR2_X1 U994 ( .A1(G227), .A2(G229), .ZN(n896) );
  XNOR2_X1 U995 ( .A(KEYINPUT49), .B(n896), .ZN(n897) );
  NOR2_X1 U996 ( .A1(G401), .A2(n897), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G395), .A2(G397), .ZN(n898) );
  AND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U999 ( .A1(n900), .A2(G319), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1002 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n1011) );
  XOR2_X1 U1003 ( .A(G2090), .B(G35), .Z(n903) );
  XOR2_X1 U1004 ( .A(G34), .B(KEYINPUT54), .Z(n901) );
  XNOR2_X1 U1005 ( .A(G2084), .B(n901), .ZN(n902) );
  NAND2_X1 U1006 ( .A1(n903), .A2(n902), .ZN(n916) );
  XNOR2_X1 U1007 ( .A(G1996), .B(G32), .ZN(n905) );
  XNOR2_X1 U1008 ( .A(G33), .B(G2072), .ZN(n904) );
  NOR2_X1 U1009 ( .A1(n905), .A2(n904), .ZN(n910) );
  XOR2_X1 U1010 ( .A(G25), .B(G1991), .Z(n906) );
  NAND2_X1 U1011 ( .A1(n906), .A2(G28), .ZN(n908) );
  XNOR2_X1 U1012 ( .A(G26), .B(G2067), .ZN(n907) );
  NOR2_X1 U1013 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1014 ( .A1(n910), .A2(n909), .ZN(n913) );
  XOR2_X1 U1015 ( .A(G27), .B(n911), .Z(n912) );
  NOR2_X1 U1016 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1017 ( .A(n914), .B(KEYINPUT53), .ZN(n915) );
  NOR2_X1 U1018 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(KEYINPUT55), .B(n917), .ZN(n918) );
  XNOR2_X1 U1020 ( .A(KEYINPUT115), .B(n918), .ZN(n919) );
  NOR2_X1 U1021 ( .A1(G29), .A2(n919), .ZN(n1008) );
  XNOR2_X1 U1022 ( .A(KEYINPUT56), .B(G16), .ZN(n948) );
  XOR2_X1 U1023 ( .A(G168), .B(G1966), .Z(n920) );
  NOR2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1025 ( .A(KEYINPUT116), .B(n922), .Z(n923) );
  XNOR2_X1 U1026 ( .A(KEYINPUT57), .B(n923), .ZN(n946) );
  XNOR2_X1 U1027 ( .A(G301), .B(G1961), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(n924), .B(G1348), .ZN(n925) );
  NOR2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1030 ( .A(KEYINPUT117), .B(n927), .Z(n940) );
  XNOR2_X1 U1031 ( .A(n928), .B(G1956), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(G1971), .A2(G303), .ZN(n929) );
  NAND2_X1 U1033 ( .A1(n930), .A2(n929), .ZN(n937) );
  INV_X1 U1034 ( .A(n931), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT118), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n944) );
  XOR2_X1 U1040 ( .A(G1341), .B(n941), .Z(n942) );
  XNOR2_X1 U1041 ( .A(KEYINPUT119), .B(n942), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n977) );
  XNOR2_X1 U1045 ( .A(G20), .B(n949), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G19), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(G1981), .B(G6), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1050 ( .A(KEYINPUT59), .B(G1348), .Z(n954) );
  XNOR2_X1 U1051 ( .A(G4), .B(n954), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(KEYINPUT120), .B(n957), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(n958), .B(KEYINPUT60), .ZN(n970) );
  XOR2_X1 U1055 ( .A(G1986), .B(KEYINPUT123), .Z(n959) );
  XNOR2_X1 U1056 ( .A(G24), .B(n959), .ZN(n965) );
  XOR2_X1 U1057 ( .A(G1976), .B(KEYINPUT121), .Z(n960) );
  XNOR2_X1 U1058 ( .A(G23), .B(n960), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(G22), .B(G1971), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1061 ( .A(KEYINPUT122), .B(n963), .Z(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1063 ( .A(KEYINPUT58), .B(n966), .Z(n968) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G21), .ZN(n967) );
  NOR2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G5), .B(G1961), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1069 ( .A(KEYINPUT61), .B(n973), .Z(n974) );
  NOR2_X1 U1070 ( .A1(G16), .A2(n974), .ZN(n975) );
  XOR2_X1 U1071 ( .A(KEYINPUT124), .B(n975), .Z(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT125), .B(n978), .ZN(n1006) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n981), .Z(n998) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(G2084), .B(G160), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(KEYINPUT113), .B(n986), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n996) );
  XOR2_X1 U1083 ( .A(G2072), .B(n991), .Z(n993) );
  XOR2_X1 U1084 ( .A(G164), .B(G2078), .Z(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1086 ( .A(KEYINPUT50), .B(n994), .Z(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1090 ( .A(KEYINPUT52), .B(n1001), .Z(n1002) );
  NOR2_X1 U1091 ( .A1(KEYINPUT55), .A2(n1002), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT114), .B(n1003), .Z(n1004) );
  NAND2_X1 U1093 ( .A1(G29), .A2(n1004), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(G11), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(n1011), .B(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(KEYINPUT62), .B(n1012), .ZN(G150) );
  INV_X1 U1099 ( .A(G150), .ZN(G311) );
endmodule

