//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n597,
    new_n599, new_n600, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n464), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n466), .B(new_n467), .C1(new_n461), .C2(new_n460), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  XOR2_X1   g045(.A(new_n470), .B(KEYINPUT69), .Z(new_n471));
  AND3_X1   g046(.A1(new_n469), .A2(KEYINPUT70), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT70), .B1(new_n469), .B2(new_n471), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n462), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n462), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n462), .A2(new_n463), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n463), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  XOR2_X1   g062(.A(new_n487), .B(KEYINPUT71), .Z(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND2_X1  g064(.A1(KEYINPUT4), .A2(G138), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT3), .ZN(new_n491));
  INV_X1    g066(.A(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n463), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n493), .B2(new_n494), .ZN(new_n499));
  AND2_X1   g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  OAI21_X1  g075(.A(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n463), .C1(new_n460), .C2(new_n461), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n497), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(G543), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT72), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI221_X1 g104(.A(new_n527), .B1(new_n528), .B2(new_n515), .C1(new_n512), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  INV_X1    g106(.A(new_n512), .ZN(new_n532));
  INV_X1    g107(.A(new_n515), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(G90), .B1(G52), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n517), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G171));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n512), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n517), .ZN(new_n541));
  AOI211_X1 g116(.A(new_n539), .B(new_n541), .C1(G43), .C2(new_n533), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n548));
  INV_X1    g123(.A(G91), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n512), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n510), .A2(KEYINPUT74), .A3(G91), .A4(new_n511), .ZN(new_n551));
  INV_X1    g126(.A(G78), .ZN(new_n552));
  INV_X1    g127(.A(G543), .ZN(new_n553));
  OR3_X1    g128(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT75), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT75), .B1(new_n552), .B2(new_n553), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n509), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n550), .A2(new_n551), .B1(G651), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n515), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n515), .B2(new_n559), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  XNOR2_X1  g138(.A(G171), .B(KEYINPUT76), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  NAND2_X1  g141(.A1(new_n533), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n568));
  INV_X1    g143(.A(G87), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n512), .ZN(G288));
  AOI22_X1  g145(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n517), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT77), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n571), .A2(KEYINPUT77), .A3(new_n517), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  INV_X1    g150(.A(G48), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n512), .A2(new_n575), .B1(new_n576), .B2(new_n515), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n574), .A3(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n532), .A2(G85), .B1(G47), .B2(new_n533), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n517), .B2(new_n581), .ZN(G290));
  AND3_X1   g157(.A1(new_n510), .A2(G92), .A3(new_n511), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT10), .ZN(new_n584));
  NAND2_X1  g159(.A1(G79), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G66), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n509), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(G54), .A2(new_n533), .B1(new_n587), .B2(G651), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(G301), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G284));
  AOI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G321));
  MUX2_X1   g169(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g170(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n589), .B1(new_n597), .B2(G860), .ZN(G148));
  NAND2_X1  g173(.A1(new_n589), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g176(.A(KEYINPUT78), .B(KEYINPUT11), .ZN(new_n602));
  XNOR2_X1  g177(.A(G323), .B(new_n602), .ZN(G282));
  XNOR2_X1  g178(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT13), .Z(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(G2100), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n481), .A2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n483), .A2(G123), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n463), .A2(G111), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2096), .Z(new_n615));
  NAND3_X1  g190(.A1(new_n608), .A2(new_n609), .A3(new_n615), .ZN(G156));
  XNOR2_X1  g191(.A(KEYINPUT15), .B(G2435), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2438), .Z(new_n618));
  XNOR2_X1  g193(.A(G2427), .B(G2430), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(KEYINPUT14), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT81), .Z(new_n622));
  INV_X1    g197(.A(new_n618), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n619), .ZN(new_n624));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n631));
  OAI21_X1  g206(.A(G14), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(G401));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT18), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(KEYINPUT17), .ZN(new_n640));
  INV_X1    g215(.A(new_n634), .ZN(new_n641));
  INV_X1    g216(.A(new_n635), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n641), .A2(new_n637), .A3(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(new_n636), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n639), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XNOR2_X1  g223(.A(G1956), .B(G2474), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1961), .B(G1966), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n651), .A2(KEYINPUT83), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n653));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(KEYINPUT83), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n652), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT20), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n649), .A3(new_n650), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n649), .B(new_n650), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n658), .B(new_n659), .C1(new_n655), .C2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G229));
  INV_X1    g242(.A(G305), .ZN(new_n668));
  INV_X1    g243(.A(G16), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(G6), .B2(new_n669), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT32), .B(G1981), .Z(new_n672));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n673));
  MUX2_X1   g248(.A(G23), .B(G288), .S(G16), .Z(new_n674));
  XOR2_X1   g249(.A(KEYINPUT33), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT84), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  AOI22_X1  g252(.A1(new_n671), .A2(new_n672), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n669), .A2(G22), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G166), .B2(new_n669), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1971), .ZN(new_n681));
  INV_X1    g256(.A(new_n677), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(KEYINPUT85), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n678), .B(new_n683), .C1(new_n672), .C2(new_n671), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n686));
  MUX2_X1   g261(.A(G24), .B(G290), .S(G16), .Z(new_n687));
  INV_X1    g262(.A(G1986), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n481), .A2(G131), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n483), .A2(G119), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n463), .A2(G107), .ZN(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT35), .B(G1991), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n685), .A2(new_n686), .A3(new_n689), .A4(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT36), .Z(new_n699));
  NOR2_X1   g274(.A1(G29), .A2(G35), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G162), .B2(G29), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT29), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(G2090), .ZN(new_n703));
  NOR3_X1   g278(.A1(KEYINPUT89), .A2(G5), .A3(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(KEYINPUT89), .B1(G5), .B2(G16), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI211_X1 g281(.A(new_n704), .B(new_n706), .C1(G171), .C2(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G1961), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT90), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n669), .A2(G4), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n589), .B2(new_n669), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1348), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n702), .A2(G2090), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n669), .A2(G20), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT23), .Z(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G299), .B2(G16), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1956), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n703), .A2(new_n713), .A3(new_n714), .A4(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G168), .A2(new_n669), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n669), .B2(G21), .ZN(new_n721));
  INV_X1    g296(.A(G1966), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT88), .Z(new_n724));
  INV_X1    g299(.A(G2084), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(KEYINPUT24), .B2(G34), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(KEYINPUT24), .B2(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n479), .B2(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n483), .A2(G129), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  AND3_X1   g307(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT26), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n733), .B(new_n735), .C1(G141), .C2(new_n481), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT87), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(KEYINPUT87), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(new_n726), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n726), .B2(G32), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT27), .B(G1996), .ZN(new_n744));
  OAI221_X1 g319(.A(new_n724), .B1(new_n725), .B2(new_n729), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n669), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n542), .B2(new_n669), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1341), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n707), .A2(G1961), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT25), .ZN(new_n751));
  OAI21_X1  g326(.A(G127), .B1(new_n460), .B2(new_n461), .ZN(new_n752));
  NAND2_X1  g327(.A1(G115), .A2(G2104), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n463), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n751), .B(new_n754), .C1(G139), .C2(new_n481), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(new_n726), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n726), .B2(G33), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n614), .A2(new_n726), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT30), .B(G28), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n760), .B(new_n761), .C1(new_n726), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n757), .A2(new_n758), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n749), .A2(new_n759), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G2078), .ZN(new_n766));
  NAND2_X1  g341(.A1(G164), .A2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G27), .B2(G29), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n748), .B(new_n765), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n726), .A2(G26), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT28), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n481), .A2(G140), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n483), .A2(G128), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n463), .A2(G116), .ZN(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n772), .B(new_n773), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n771), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2067), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n766), .B2(new_n768), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n722), .B2(new_n721), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n729), .A2(new_n725), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n743), .A2(new_n744), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n769), .A2(new_n780), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n699), .A2(new_n719), .A3(new_n745), .A4(new_n783), .ZN(G311));
  INV_X1    g359(.A(G311), .ZN(G150));
  NAND2_X1  g360(.A1(new_n589), .A2(G559), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT92), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT38), .Z(new_n788));
  AND2_X1   g363(.A1(new_n510), .A2(G67), .ZN(new_n789));
  AND2_X1   g364(.A1(G80), .A2(G543), .ZN(new_n790));
  OAI21_X1  g365(.A(G651), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT91), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n532), .A2(G93), .B1(G55), .B2(new_n533), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(KEYINPUT91), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(new_n542), .Z(new_n797));
  XOR2_X1   g372(.A(new_n788), .B(new_n797), .Z(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(KEYINPUT39), .ZN(new_n799));
  INV_X1    g374(.A(G860), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(KEYINPUT39), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n796), .A2(new_n800), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT93), .B(KEYINPUT37), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n805), .ZN(G145));
  XNOR2_X1  g381(.A(new_n479), .B(new_n614), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(new_n488), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n740), .B(new_n505), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(new_n776), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(new_n755), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n483), .A2(G130), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n463), .A2(G118), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G142), .B2(new_n481), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(new_n694), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n606), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT94), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n811), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n811), .A2(new_n819), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n808), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g399(.A(KEYINPUT95), .B(new_n808), .C1(new_n820), .C2(new_n821), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n820), .A2(new_n808), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n810), .B(new_n755), .Z(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(new_n818), .ZN(new_n829));
  AOI21_X1  g404(.A(G37), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g407(.A1(new_n589), .A2(G299), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT96), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n589), .A2(G299), .ZN(new_n835));
  AOI21_X1  g410(.A(KEYINPUT41), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n833), .A2(KEYINPUT41), .A3(new_n835), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n797), .B(new_n599), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n833), .A2(new_n835), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(G305), .B(G290), .ZN(new_n843));
  XOR2_X1   g418(.A(G166), .B(G288), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT97), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT42), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n845), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n842), .B1(new_n849), .B2(KEYINPUT98), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(KEYINPUT98), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n849), .A2(new_n842), .A3(KEYINPUT98), .ZN(new_n853));
  OAI21_X1  g428(.A(G868), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n796), .A2(G868), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G295));
  XNOR2_X1  g432(.A(G295), .B(KEYINPUT99), .ZN(G331));
  NOR2_X1   g433(.A1(G168), .A2(G171), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n592), .B2(G168), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n797), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT100), .Z(new_n862));
  OR2_X1    g437(.A1(new_n860), .A2(new_n797), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n841), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n863), .A2(new_n861), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n862), .A2(new_n864), .B1(new_n838), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n846), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n866), .A2(new_n867), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT43), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n834), .A2(KEYINPUT41), .A3(new_n835), .ZN(new_n873));
  INV_X1    g448(.A(new_n841), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(KEYINPUT41), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n863), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n862), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n863), .A2(new_n841), .A3(new_n861), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(new_n867), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n880), .A2(new_n868), .A3(new_n881), .A4(new_n869), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(KEYINPUT44), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n868), .A3(new_n869), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT43), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT101), .ZN(new_n887));
  OR3_X1    g462(.A1(new_n870), .A2(KEYINPUT43), .A3(new_n871), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n889), .A3(KEYINPUT43), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n884), .B1(new_n891), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g467(.A1(new_n469), .A2(new_n471), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT70), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT70), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n478), .A2(G40), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G1384), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n505), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n696), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n694), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G1996), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n740), .B(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G2067), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n776), .B(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n906), .B1(new_n911), .B2(new_n904), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n776), .A2(G2067), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n904), .B1(new_n914), .B2(KEYINPUT125), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(KEYINPUT125), .B2(new_n914), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n903), .A2(KEYINPUT46), .A3(new_n907), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n904), .B2(G1996), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n741), .A2(new_n910), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n917), .B(new_n919), .C1(new_n920), .C2(new_n904), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT47), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n904), .A2(G1986), .A3(G290), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(KEYINPUT48), .Z(new_n924));
  XNOR2_X1  g499(.A(new_n694), .B(new_n696), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n911), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n926), .B2(new_n904), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n916), .A2(new_n922), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT126), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT126), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n916), .A2(new_n930), .A3(new_n922), .A4(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G1976), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT52), .B1(G288), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n898), .A2(new_n900), .ZN(new_n935));
  INV_X1    g510(.A(G8), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n933), .B2(G288), .ZN(new_n938));
  MUX2_X1   g513(.A(new_n934), .B(KEYINPUT52), .S(new_n938), .Z(new_n939));
  NOR2_X1   g514(.A1(G305), .A2(G1981), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n577), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n572), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n577), .A2(new_n941), .ZN(new_n944));
  OAI21_X1  g519(.A(G1981), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n940), .B1(new_n945), .B2(KEYINPUT108), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n945), .A2(KEYINPUT108), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(KEYINPUT49), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT49), .B1(new_n946), .B2(new_n947), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n951), .A2(new_n936), .A3(new_n935), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n939), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(G303), .A2(G8), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT106), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n954), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(KEYINPUT55), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n954), .A2(new_n955), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n901), .A2(G1384), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n505), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n505), .A2(KEYINPUT102), .A3(new_n962), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n902), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT103), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n902), .A2(new_n965), .A3(new_n966), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n970), .A2(new_n971), .A3(new_n898), .ZN(new_n972));
  OR3_X1    g547(.A1(new_n969), .A2(new_n972), .A3(G1971), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n505), .A2(new_n974), .A3(new_n899), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n974), .B1(new_n505), .B2(new_n899), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n900), .A2(KEYINPUT105), .A3(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n968), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI22_X1  g557(.A1(new_n973), .A2(KEYINPUT104), .B1(G2090), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n973), .A2(KEYINPUT104), .ZN(new_n984));
  OAI211_X1 g559(.A(G8), .B(new_n961), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n900), .A2(KEYINPUT50), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n474), .A2(new_n986), .A3(new_n897), .A4(new_n975), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n973), .B1(G2090), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G8), .ZN(new_n989));
  INV_X1    g564(.A(new_n961), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND4_X1   g566(.A1(new_n895), .A2(new_n963), .A3(new_n896), .A4(new_n897), .ZN(new_n992));
  AOI21_X1  g567(.A(G1966), .B1(new_n992), .B2(new_n902), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n725), .B(new_n968), .C1(new_n979), .C2(new_n981), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(KEYINPUT110), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n895), .A2(new_n725), .A3(new_n897), .A4(new_n896), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n986), .A2(new_n976), .A3(new_n975), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(new_n980), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n936), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G168), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n953), .A2(new_n985), .A3(new_n991), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT63), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(G8), .B1(new_n983), .B2(new_n984), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n990), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n985), .A3(new_n953), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n985), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n953), .ZN(new_n1013));
  AOI211_X1 g588(.A(G1976), .B(G288), .C1(new_n950), .C2(new_n952), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n937), .B1(new_n1014), .B2(new_n940), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G286), .A2(G8), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n998), .A2(new_n999), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n968), .A2(new_n963), .A3(new_n902), .ZN(new_n1022));
  OAI22_X1  g597(.A1(new_n999), .A2(new_n998), .B1(new_n1022), .B2(G1966), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1020), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1019), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1001), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1023), .B2(new_n1021), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1029), .A2(KEYINPUT120), .A3(new_n1026), .A4(new_n1019), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1026), .B1(new_n1029), .B2(new_n1019), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1028), .B(new_n1030), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1024), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT62), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(G2078), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1022), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n997), .A2(new_n980), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT114), .B1(new_n1041), .B2(new_n968), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n1043));
  AOI211_X1 g618(.A(new_n1043), .B(new_n898), .C1(new_n997), .C2(new_n980), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1961), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1040), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n766), .B1(new_n969), .B2(new_n972), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(new_n1037), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n971), .B1(new_n970), .B2(new_n898), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n964), .A2(new_n963), .B1(new_n900), .B2(new_n901), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(new_n968), .A3(KEYINPUT103), .A4(new_n966), .ZN(new_n1053));
  AOI21_X1  g628(.A(G2078), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1054), .A2(KEYINPUT121), .A3(KEYINPUT53), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1047), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n592), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n1024), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1036), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT124), .B1(new_n1056), .B2(new_n592), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n897), .A2(new_n1038), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n474), .B2(KEYINPUT122), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n970), .B(new_n1065), .C1(KEYINPUT122), .C2(new_n474), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1063), .B1(new_n1068), .B2(G171), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n982), .A2(new_n1043), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1041), .A2(KEYINPUT114), .A3(new_n968), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1046), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1039), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT121), .B1(new_n1054), .B2(KEYINPUT53), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1049), .A2(new_n1048), .A3(new_n1037), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1077), .A3(G301), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1062), .A2(new_n1069), .A3(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1067), .B(G301), .C1(new_n1050), .C2(new_n1055), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT123), .B(KEYINPUT54), .C1(new_n1057), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1076), .B2(G301), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(new_n1063), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1035), .B(new_n1079), .C1(new_n1081), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1348), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1070), .A2(new_n1086), .A3(new_n1071), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n935), .A2(new_n909), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n589), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1087), .A2(KEYINPUT60), .A3(new_n590), .A4(new_n1088), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1091), .A2(new_n1092), .B1(new_n1090), .B2(new_n1089), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n970), .A2(new_n898), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n907), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT58), .B(G1341), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n935), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n542), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT59), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1100), .A3(new_n542), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n558), .A2(KEYINPUT57), .A3(new_n562), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n558), .A2(KEYINPUT113), .A3(KEYINPUT57), .A4(new_n562), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT112), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n562), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n558), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n562), .A2(new_n1109), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1107), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1094), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n987), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n987), .B2(new_n1118), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1114), .B(new_n1116), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT116), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n987), .A2(new_n1118), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT111), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n987), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1114), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1122), .A2(new_n1128), .A3(KEYINPUT61), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1121), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1114), .B1(new_n1126), .B2(new_n1116), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1129), .A2(KEYINPUT115), .A3(new_n1130), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1102), .B(new_n1132), .C1(new_n1136), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1093), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1143), .A2(KEYINPUT117), .A3(new_n1132), .A4(new_n1102), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1089), .A2(new_n589), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1131), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1142), .A2(new_n1144), .B1(new_n1146), .B2(new_n1121), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1061), .B1(new_n1085), .B2(new_n1147), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n953), .A2(new_n985), .A3(new_n991), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1016), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(G290), .B(new_n688), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n904), .B1(new_n926), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n932), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT127), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1155), .B(new_n932), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g732(.A(G319), .ZN(new_n1159));
  NOR4_X1   g733(.A1(G401), .A2(new_n1159), .A3(G229), .A4(G227), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n831), .A2(new_n883), .A3(new_n1160), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


