//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n192), .B1(new_n189), .B2(new_n191), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT0), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT64), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(KEYINPUT0), .B2(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n198), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n187), .B1(new_n197), .B2(new_n205), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n190), .A2(KEYINPUT1), .A3(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n189), .A2(new_n191), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(new_n200), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n189), .A3(new_n191), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n187), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G224), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G953), .ZN(new_n216));
  XOR2_X1   g030(.A(new_n214), .B(new_n216), .Z(new_n217));
  XNOR2_X1  g031(.A(G116), .B(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT5), .ZN(new_n219));
  INV_X1    g033(.A(G113), .ZN(new_n220));
  INV_X1    g034(.A(G116), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(G119), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT5), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(KEYINPUT2), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G113), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n229), .A2(new_n218), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n229), .B2(new_n218), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n225), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT3), .B1(new_n234), .B2(G107), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n236));
  INV_X1    g050(.A(G107), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G104), .ZN(new_n238));
  INV_X1    g052(.A(G101), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(G107), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n235), .A2(new_n238), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT83), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(G104), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n240), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n244), .B2(G101), .ZN(new_n245));
  AOI211_X1 g059(.A(KEYINPUT83), .B(new_n239), .C1(new_n243), .C2(new_n240), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT86), .B1(new_n233), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G116), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n221), .A2(G119), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT2), .B(G113), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n229), .A2(new_n218), .A3(new_n230), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n254), .A2(new_n255), .B1(new_n219), .B2(new_n224), .ZN(new_n256));
  XNOR2_X1  g070(.A(G104), .B(G107), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT83), .B1(new_n257), .B2(new_n239), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n244), .A2(new_n242), .A3(G101), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n235), .A2(new_n238), .A3(new_n240), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n258), .A2(new_n259), .B1(new_n260), .B2(new_n239), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT86), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n256), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n252), .A2(new_n253), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n231), .B2(new_n232), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n235), .A2(new_n238), .A3(new_n240), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G101), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT4), .A3(new_n241), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n269), .A3(G101), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G122), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n248), .A2(new_n263), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n248), .A2(new_n271), .A3(new_n263), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n272), .A2(KEYINPUT87), .ZN(new_n275));
  AOI22_X1  g089(.A1(KEYINPUT6), .A2(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n274), .A2(KEYINPUT6), .A3(new_n275), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n217), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT7), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n216), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n206), .B2(new_n213), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n194), .A2(new_n196), .B1(new_n204), .B2(new_n198), .ZN(new_n282));
  OAI221_X1 g096(.A(new_n212), .B1(new_n279), .B2(new_n216), .C1(new_n282), .C2(new_n187), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n272), .B(KEYINPUT8), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n233), .A2(new_n247), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n254), .A2(new_n255), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n258), .A2(new_n259), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n287), .A2(new_n225), .B1(new_n288), .B2(new_n241), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n285), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n273), .A2(new_n284), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n278), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT89), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n278), .B(new_n297), .C1(new_n294), .C2(new_n295), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n301), .A2(new_n300), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT21), .B(G898), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n304), .B(KEYINPUT96), .ZN(new_n305));
  INV_X1    g119(.A(G953), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n293), .B(new_n306), .C1(G234), .C2(G237), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G952), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n309), .A2(KEYINPUT95), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(KEYINPUT95), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(G234), .B2(G237), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT97), .Z(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G214), .B1(G237), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n302), .A2(new_n303), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G221), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT9), .B(G234), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n325), .B2(new_n293), .ZN(new_n326));
  INV_X1    g140(.A(G469), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n293), .ZN(new_n328));
  XNOR2_X1  g142(.A(G110), .B(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n306), .A2(G227), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n211), .A2(KEYINPUT84), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n210), .A2(new_n189), .A3(new_n191), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n209), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n241), .A3(new_n288), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(new_n209), .B2(new_n211), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n339), .A2(new_n340), .B1(new_n261), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT11), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G137), .ZN(new_n344));
  AND2_X1   g158(.A1(KEYINPUT67), .A2(G134), .ZN(new_n345));
  NOR2_X1   g159(.A1(KEYINPUT67), .A2(G134), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G137), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT11), .A3(G134), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(G137), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G131), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n351), .ZN(new_n353));
  OR2_X1    g167(.A1(KEYINPUT67), .A2(G134), .ZN(new_n354));
  NAND2_X1  g168(.A1(KEYINPUT67), .A2(G134), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n354), .B(new_n355), .C1(new_n343), .C2(G137), .ZN(new_n356));
  INV_X1    g170(.A(G131), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n352), .A2(new_n358), .A3(KEYINPUT70), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT70), .B1(new_n352), .B2(new_n358), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n197), .A2(new_n205), .A3(new_n270), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(new_n268), .ZN(new_n364));
  AND4_X1   g178(.A1(new_n362), .A2(new_n268), .A3(new_n282), .A4(new_n270), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n342), .B(new_n361), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n268), .A2(new_n282), .A3(new_n270), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT82), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n268), .A2(new_n282), .A3(new_n362), .A4(new_n270), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n361), .B1(new_n371), .B2(new_n342), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n334), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n209), .A2(new_n211), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n261), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n209), .A2(new_n211), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n247), .A2(new_n377), .A3(KEYINPUT85), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n376), .A2(new_n378), .B1(new_n261), .B2(new_n338), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n352), .A2(new_n358), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT12), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n261), .A2(new_n374), .A3(new_n375), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT85), .B1(new_n247), .B2(new_n377), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n339), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT70), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n347), .A2(G131), .A3(new_n351), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n357), .B1(new_n353), .B2(new_n356), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n352), .A2(new_n358), .A3(KEYINPUT70), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT12), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n382), .A2(new_n366), .A3(new_n333), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(G902), .B1(new_n373), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n328), .B1(new_n394), .B2(new_n327), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n366), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT12), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n385), .B2(new_n380), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n334), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n372), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n366), .A3(new_n333), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n401), .A3(G469), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n326), .B1(new_n395), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G116), .B(G122), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n237), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT94), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n345), .A2(new_n346), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n190), .A2(G128), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n200), .A2(G143), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n354), .A2(new_n355), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n410), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT14), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n404), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n221), .A2(KEYINPUT14), .A3(G122), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n417), .A2(G107), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n411), .A2(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n412), .A2(new_n413), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n404), .A2(new_n237), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n420), .B1(new_n421), .B2(new_n405), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT13), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n409), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n410), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n409), .A2(new_n423), .ZN(new_n426));
  OAI21_X1  g240(.A(G134), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n407), .A2(new_n419), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G217), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n324), .A2(new_n429), .A3(G953), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n428), .A2(new_n430), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n293), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G478), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT15), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n434), .B(new_n436), .Z(new_n437));
  XNOR2_X1  g251(.A(G113), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(new_n234), .ZN(new_n439));
  OR3_X1    g253(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT75), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n443));
  XNOR2_X1  g257(.A(G125), .B(G140), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(KEYINPUT16), .ZN(new_n445));
  OAI211_X1 g259(.A(G146), .B(new_n442), .C1(new_n445), .C2(new_n441), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(KEYINPUT91), .A2(KEYINPUT19), .ZN(new_n449));
  INV_X1    g263(.A(G140), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G125), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n187), .A2(G140), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n444), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(G237), .A2(G953), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(G143), .A3(G214), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G143), .B1(new_n456), .B2(G214), .ZN(new_n459));
  OAI21_X1  g273(.A(G131), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G237), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n306), .A3(G214), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n190), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n357), .A3(new_n457), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n455), .A2(new_n188), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT16), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n441), .B1(new_n466), .B2(new_n440), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(KEYINPUT76), .A3(G146), .A4(new_n442), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n448), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n457), .ZN(new_n471));
  AND2_X1   g285(.A1(KEYINPUT18), .A2(G131), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n451), .A2(new_n452), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G146), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n444), .A2(new_n188), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n471), .A2(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n458), .A2(new_n459), .ZN(new_n477));
  INV_X1    g291(.A(new_n472), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT90), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n471), .A2(new_n480), .A3(new_n472), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n476), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n439), .B1(new_n470), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n439), .B(KEYINPUT92), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n460), .A2(new_n485), .A3(new_n464), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n443), .A2(KEYINPUT75), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n188), .B1(new_n467), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n471), .A2(KEYINPUT17), .A3(G131), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n486), .A2(new_n488), .A3(new_n446), .A4(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n484), .A2(new_n490), .A3(new_n482), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n493));
  NOR2_X1   g307(.A1(G475), .A2(G902), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n492), .A2(KEYINPUT93), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n493), .B(new_n494), .C1(new_n483), .C2(new_n491), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n483), .A2(new_n491), .ZN(new_n499));
  INV_X1    g313(.A(new_n494), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT20), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n439), .B1(new_n490), .B2(new_n482), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n293), .B1(new_n491), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G475), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n437), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n322), .A2(KEYINPUT98), .A3(new_n403), .A4(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT32), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT68), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n412), .A2(new_n509), .A3(new_n348), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n408), .A2(G137), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT68), .B1(new_n348), .B2(G134), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(G131), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n358), .A3(new_n375), .ZN(new_n514));
  OAI22_X1  g328(.A1(new_n282), .A2(KEYINPUT66), .B1(new_n387), .B2(new_n388), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n197), .A2(KEYINPUT66), .A3(new_n205), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n282), .B1(new_n359), .B2(new_n360), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT30), .A3(new_n514), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n521), .A3(new_n265), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n523));
  NAND2_X1  g337(.A1(new_n456), .A2(G210), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT26), .B(G101), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n513), .A2(new_n358), .A3(new_n375), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n389), .A2(new_n390), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n529), .B1(new_n530), .B2(new_n282), .ZN(new_n531));
  INV_X1    g345(.A(new_n265), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n522), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n522), .A2(new_n533), .A3(KEYINPUT31), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n517), .A2(new_n265), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT28), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n531), .B2(new_n532), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n539), .A2(new_n520), .A3(new_n532), .A4(new_n514), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n536), .A2(new_n537), .B1(new_n528), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G472), .A2(G902), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n508), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n522), .A2(KEYINPUT31), .A3(new_n533), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT31), .B1(new_n522), .B2(new_n533), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n531), .A2(new_n539), .A3(new_n532), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n520), .A2(new_n532), .A3(new_n514), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT28), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n549), .A2(new_n551), .B1(new_n265), .B2(new_n517), .ZN(new_n552));
  OAI22_X1  g366(.A1(new_n547), .A2(new_n548), .B1(new_n552), .B2(new_n527), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT32), .A3(new_n544), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n554), .A3(KEYINPUT72), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n544), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT72), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n508), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G472), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT73), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n542), .B2(new_n528), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n552), .A2(KEYINPUT73), .A3(new_n527), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT29), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n522), .A2(new_n550), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n528), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n562), .A2(new_n563), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n531), .A2(new_n532), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n551), .B2(new_n549), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n528), .A2(new_n564), .ZN(new_n570));
  AOI21_X1  g384(.A(G902), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n560), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n559), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n403), .A2(new_n506), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n575), .B1(new_n576), .B2(new_n321), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n429), .B1(G234), .B2(new_n293), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT22), .B(G137), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n306), .A2(G221), .A3(G234), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n581), .B(new_n582), .Z(new_n583));
  INV_X1    g397(.A(KEYINPUT78), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT74), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n200), .A2(G119), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n200), .A2(G119), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT23), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G110), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n585), .B1(new_n249), .B2(G128), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n249), .A2(G128), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(KEYINPUT23), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n586), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT24), .B(G110), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n594), .A2(new_n597), .B1(new_n188), .B2(new_n444), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n448), .A2(new_n469), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT77), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n448), .A2(new_n469), .A3(KEYINPUT77), .A4(new_n598), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n589), .A2(new_n593), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n604), .A2(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n446), .B2(new_n488), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n584), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  AOI211_X1 g422(.A(KEYINPUT78), .B(new_n606), .C1(new_n601), .C2(new_n602), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n583), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n583), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n603), .A2(new_n607), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n611), .B1(new_n612), .B2(KEYINPUT78), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n580), .B1(new_n614), .B2(G902), .ZN(new_n615));
  INV_X1    g429(.A(new_n580), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n610), .A2(new_n293), .A3(new_n616), .A4(new_n613), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n579), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n614), .A2(G902), .A3(new_n578), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n507), .A2(new_n574), .A3(new_n577), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  INV_X1    g436(.A(new_n403), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n623), .A2(new_n618), .A3(new_n619), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n560), .B1(new_n553), .B2(new_n293), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n625), .A2(KEYINPUT99), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n556), .B1(new_n625), .B2(KEYINPUT99), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n319), .B1(new_n299), .B2(new_n301), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n434), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT101), .B(G478), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n428), .B2(new_n430), .ZN(new_n636));
  OAI211_X1 g450(.A(KEYINPUT33), .B(new_n636), .C1(new_n432), .C2(new_n433), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n428), .A2(new_n430), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n638), .B(new_n431), .C1(new_n635), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n435), .A2(G902), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n502), .A2(new_n505), .B1(new_n634), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n631), .A2(new_n645), .A3(new_n317), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n629), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NAND2_X1  g463(.A1(new_n501), .A2(new_n496), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n505), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n631), .A2(new_n317), .A3(new_n437), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n629), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G107), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT102), .B(KEYINPUT35), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NAND2_X1  g470(.A1(new_n507), .A2(new_n577), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n615), .A2(new_n617), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n578), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n611), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n612), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n578), .A2(G902), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n659), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n664), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT103), .B1(new_n618), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(new_n628), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n657), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT37), .B(G110), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G12));
  NAND2_X1  g485(.A1(new_n403), .A2(new_n630), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n559), .B2(new_n573), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n313), .B1(new_n674), .B2(new_n307), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n651), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n437), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n673), .A2(new_n667), .A3(new_n665), .A4(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT104), .B(G128), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G30));
  XOR2_X1   g496(.A(new_n675), .B(KEYINPUT39), .Z(new_n683));
  NAND2_X1  g497(.A1(new_n403), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT40), .Z(new_n685));
  NAND2_X1  g499(.A1(new_n302), .A2(new_n303), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n319), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n502), .A2(new_n505), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n677), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n618), .A2(new_n666), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n528), .B1(new_n522), .B2(new_n550), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n550), .A2(new_n528), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n293), .B1(new_n694), .B2(new_n568), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n559), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n685), .A2(new_n689), .A3(new_n692), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  INV_X1    g513(.A(new_n675), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n644), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT106), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n673), .A2(new_n667), .A3(new_n665), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  INV_X1    g518(.A(new_n620), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n572), .B1(new_n555), .B2(new_n558), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n394), .A2(new_n327), .ZN(new_n708));
  INV_X1    g522(.A(new_n326), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n394), .A2(new_n327), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n707), .A2(new_n646), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT107), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n713), .B(new_n715), .ZN(G15));
  NAND3_X1  g530(.A1(new_n707), .A2(new_n652), .A3(new_n712), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  AND2_X1   g532(.A1(new_n665), .A2(new_n667), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n631), .A2(new_n711), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n720), .A2(new_n316), .A3(new_n506), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n574), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  OAI22_X1  g537(.A1(new_n547), .A2(new_n548), .B1(new_n569), .B2(new_n527), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(new_n544), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n625), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n620), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n631), .A2(new_n691), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n316), .A3(new_n712), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NOR2_X1   g545(.A1(new_n618), .A2(new_n666), .ZN(new_n732));
  INV_X1    g546(.A(new_n726), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n702), .A3(new_n720), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  AOI21_X1  g550(.A(new_n319), .B1(new_n302), .B2(new_n303), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n399), .A2(new_n401), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT108), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n401), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(G469), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n326), .B1(new_n742), .B2(new_n395), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n737), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n744), .B1(new_n737), .B2(new_n743), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n702), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n574), .A2(new_n620), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT110), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n737), .A2(new_n743), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT109), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n737), .A2(new_n743), .A3(new_n744), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n707), .A3(new_n755), .A4(new_n702), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n749), .A2(new_n750), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n554), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n553), .A2(KEYINPUT111), .A3(KEYINPUT32), .A4(new_n544), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n573), .A2(new_n760), .A3(new_n546), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n620), .A3(KEYINPUT42), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n758), .B1(new_n747), .B2(new_n763), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n762), .A2(new_n620), .A3(KEYINPUT42), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n754), .A3(KEYINPUT112), .A4(new_n702), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n757), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G131), .ZN(G33));
  NOR3_X1   g583(.A1(new_n705), .A2(new_n706), .A3(new_n678), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n754), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  NAND2_X1  g586(.A1(new_n634), .A2(new_n643), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n505), .A3(new_n502), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT43), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n628), .A2(new_n732), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT115), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT115), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n737), .B1(new_n779), .B2(KEYINPUT44), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(KEYINPUT44), .B2(new_n779), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n327), .B1(new_n738), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT113), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n739), .A2(KEYINPUT45), .A3(new_n741), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(KEYINPUT113), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n328), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(KEYINPUT114), .A3(new_n710), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n787), .A2(new_n788), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n790), .B1(KEYINPUT46), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT114), .B1(new_n789), .B2(new_n710), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n709), .B(new_n683), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n781), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  OAI21_X1  g611(.A(new_n709), .B1(new_n792), .B2(new_n793), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT47), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(KEYINPUT47), .B(new_n709), .C1(new_n792), .C2(new_n793), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n737), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n574), .A2(new_n620), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n702), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  NAND2_X1  g620(.A1(new_n712), .A2(new_n737), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n775), .A2(KEYINPUT119), .A3(new_n314), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT119), .B1(new_n775), .B2(new_n314), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n762), .A2(new_n620), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT48), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n727), .B1(new_n808), .B2(new_n809), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n720), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n697), .A2(new_n705), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n313), .A3(new_n712), .A4(new_n737), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n645), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n312), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n813), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n817), .A2(new_n690), .A3(new_n773), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n810), .A2(new_n734), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n688), .A2(new_n319), .A3(new_n712), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n814), .A2(KEYINPUT50), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT50), .B1(new_n814), .B2(new_n823), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n821), .B(new_n822), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n708), .A2(new_n710), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n326), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n800), .A2(new_n801), .A3(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n814), .A2(new_n737), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n826), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n820), .B1(new_n831), .B2(KEYINPUT51), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(KEYINPUT51), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(KEYINPUT120), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n831), .A2(new_n835), .A3(KEYINPUT51), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n832), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n713), .A2(new_n722), .A3(new_n717), .A4(new_n730), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n734), .B(new_n702), .C1(new_n745), .C2(new_n746), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n403), .A2(new_n437), .A3(new_n676), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n706), .A2(new_n841), .A3(new_n803), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n719), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n771), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n302), .A2(new_n644), .A3(new_n303), .A4(new_n320), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n677), .A2(new_n505), .A3(new_n502), .ZN(new_n847));
  OAI22_X1  g661(.A1(new_n845), .A2(new_n846), .B1(new_n321), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n628), .B(new_n624), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n850), .B(new_n621), .C1(new_n657), .C2(new_n668), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n768), .A2(new_n839), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n631), .A2(new_n675), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n697), .A2(new_n692), .A3(new_n743), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n680), .A2(new_n703), .A3(new_n735), .A4(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT52), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT53), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n680), .A2(new_n735), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(KEYINPUT52), .A3(new_n703), .A4(new_n855), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n838), .B1(new_n757), .B2(new_n767), .ZN(new_n864));
  XOR2_X1   g678(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n852), .A4(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n858), .A2(KEYINPUT54), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n865), .B1(new_n853), .B2(new_n857), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n754), .A2(new_n770), .B1(new_n719), .B2(new_n842), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n665), .A2(new_n628), .A3(new_n667), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n577), .B(new_n507), .C1(new_n871), .C2(new_n707), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n870), .A2(new_n872), .A3(new_n850), .A4(new_n840), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n869), .B1(new_n873), .B2(KEYINPUT118), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n852), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n874), .A2(new_n863), .A3(new_n876), .A4(new_n864), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n868), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n837), .A2(new_n880), .B1(G952), .B2(G953), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n774), .A2(new_n319), .A3(new_n326), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n827), .B(KEYINPUT49), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n816), .A2(new_n688), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n306), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n293), .B1(new_n868), .B2(new_n877), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(G210), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n276), .A2(new_n277), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n217), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n887), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n892), .B(KEYINPUT121), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n868), .A2(new_n877), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(G902), .ZN(new_n897));
  INV_X1    g711(.A(G210), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n894), .B(new_n895), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(KEYINPUT122), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(KEYINPUT122), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n893), .B1(new_n900), .B2(new_n901), .ZN(G51));
  NAND2_X1  g716(.A1(new_n896), .A2(KEYINPUT54), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n904), .A3(new_n879), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n896), .A2(KEYINPUT123), .A3(KEYINPUT54), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n328), .B(KEYINPUT57), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n373), .A2(new_n393), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n897), .A2(new_n787), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n886), .B1(new_n910), .B2(new_n911), .ZN(G54));
  AND3_X1   g726(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n887), .B1(new_n913), .B2(new_n492), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n492), .B2(new_n913), .ZN(G60));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT59), .Z(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n867), .B2(new_n879), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n887), .B1(new_n918), .B2(new_n641), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n905), .A2(new_n906), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n917), .B1(new_n637), .B2(new_n640), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G63));
  XNOR2_X1  g736(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n429), .A2(new_n293), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n896), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n614), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n896), .A2(new_n662), .A3(new_n925), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n887), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT61), .B1(new_n928), .B2(KEYINPUT125), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G66));
  OAI21_X1  g745(.A(G953), .B1(new_n305), .B2(new_n215), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n838), .A2(new_n851), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n890), .B1(G898), .B2(new_n306), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G69));
  NAND2_X1  g750(.A1(new_n519), .A2(new_n521), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n455), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n684), .B(new_n803), .C1(new_n645), .C2(new_n847), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n707), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT126), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n781), .B2(new_n795), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n859), .A2(new_n698), .A3(new_n703), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT62), .Z(new_n944));
  AND3_X1   g758(.A1(new_n942), .A2(new_n805), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n938), .B1(new_n945), .B2(G953), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n938), .B1(G900), .B2(G953), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n811), .A2(new_n729), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n795), .B1(new_n781), .B2(new_n948), .ZN(new_n949));
  AND4_X1   g763(.A1(new_n703), .A2(new_n768), .A3(new_n771), .A4(new_n859), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n949), .A2(new_n805), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n951), .B2(G953), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n306), .B1(G227), .B2(G900), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n954), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n946), .A2(new_n956), .A3(new_n952), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(G72));
  NAND4_X1  g772(.A1(new_n942), .A2(new_n805), .A3(new_n933), .A4(new_n944), .ZN(new_n959));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT63), .Z(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(KEYINPUT127), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n693), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT127), .B1(new_n959), .B2(new_n961), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n566), .A2(new_n534), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n858), .A2(new_n866), .A3(new_n961), .A4(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n949), .A2(new_n805), .A3(new_n933), .A4(new_n950), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n968), .A2(new_n961), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n522), .A2(new_n528), .A3(new_n550), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n887), .B(new_n967), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n965), .A2(new_n971), .ZN(G57));
endmodule


