//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G107), .A2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n209), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g0019(.A1(G58), .A2(G232), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NOR2_X1   g0022(.A1(G58), .A2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT66), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AND2_X1   g0028(.A1(KEYINPUT65), .A2(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(KEYINPUT65), .A2(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n226), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  OR3_X1    g0032(.A1(new_n208), .A2(KEYINPUT64), .A3(G13), .ZN(new_n233));
  OAI21_X1  g0033(.A(KEYINPUT64), .B1(new_n208), .B2(G13), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n235), .B(G250), .C1(G257), .C2(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT0), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n222), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G264), .ZN(new_n246));
  INV_X1    g0046(.A(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n244), .B(new_n248), .Z(G358));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n227), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n205), .A2(G20), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n260), .A2(G50), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G50), .B2(new_n261), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT71), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n263), .B(KEYINPUT71), .C1(G50), .C2(new_n261), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g0068(.A(KEYINPUT69), .B(G58), .Z(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT8), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT65), .B(G20), .ZN(new_n271));
  OR2_X1    g0071(.A1(KEYINPUT8), .A2(G58), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n270), .A2(G33), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G150), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n206), .B1(new_n223), .B2(new_n215), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n273), .A2(KEYINPUT70), .A3(new_n275), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n268), .B(KEYINPUT9), .C1(new_n283), .C2(new_n260), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G1), .A3(G13), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n291), .B2(new_n217), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G222), .ZN(new_n294));
  INV_X1    g0094(.A(G223), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n290), .B(new_n294), .C1(new_n295), .C2(new_n293), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n287), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n289), .A2(new_n285), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G190), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT74), .B(G200), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n284), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n260), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n282), .A2(new_n308), .B1(new_n266), .B2(new_n267), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT10), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n309), .A2(KEYINPUT9), .B1(new_n301), .B2(new_n305), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n268), .B1(new_n283), .B2(new_n260), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n312), .A2(new_n315), .A3(new_n316), .A4(new_n303), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n302), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT72), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n301), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n313), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT69), .B(G58), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n224), .B1(new_n326), .B2(new_n211), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(G20), .B1(G159), .B2(new_n274), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT79), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(G33), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(KEYINPUT3), .A2(G33), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n206), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT7), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n333), .A2(new_n271), .A3(new_n338), .A4(new_n335), .ZN(new_n339));
  AND4_X1   g0139(.A1(KEYINPUT80), .A2(new_n337), .A3(G68), .A4(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n211), .B1(new_n336), .B2(KEYINPUT7), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT80), .B1(new_n341), .B2(new_n339), .ZN(new_n342));
  OAI211_X1 g0142(.A(KEYINPUT16), .B(new_n328), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n258), .ZN(new_n344));
  INV_X1    g0144(.A(G33), .ZN(new_n345));
  AND2_X1   g0145(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(KEYINPUT3), .A2(G33), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n348), .A2(new_n271), .A3(KEYINPUT7), .A4(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n338), .B1(new_n290), .B2(G20), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G68), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n328), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n344), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n343), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n289), .A2(G232), .A3(new_n285), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT81), .ZN(new_n360));
  INV_X1    g0160(.A(new_n287), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n293), .A2(G226), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n333), .B2(new_n335), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n295), .A2(new_n293), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n363), .A2(new_n364), .B1(G33), .B2(G87), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n360), .B(new_n361), .C1(new_n365), .C2(new_n289), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G200), .ZN(new_n367));
  INV_X1    g0167(.A(new_n362), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n346), .A2(new_n347), .A3(new_n345), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n364), .B(new_n368), .C1(new_n369), .C2(new_n334), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n289), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n287), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(G190), .A3(new_n360), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n270), .A2(new_n272), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n375), .A2(new_n261), .A3(new_n260), .A4(new_n262), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n270), .A2(new_n272), .ZN(new_n377));
  INV_X1    g0177(.A(new_n261), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n358), .A2(new_n367), .A3(new_n374), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n380), .B1(new_n343), .B2(new_n357), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n385), .A2(KEYINPUT17), .A3(new_n367), .A4(new_n374), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n373), .A2(G179), .A3(new_n360), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n366), .A2(G169), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n327), .A2(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n274), .A2(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n211), .B1(new_n351), .B2(new_n352), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n356), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n258), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n337), .A2(G68), .A3(new_n339), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT80), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n341), .A2(KEYINPUT80), .A3(new_n339), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n393), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n396), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  OAI211_X1 g0202(.A(KEYINPUT18), .B(new_n390), .C1(new_n402), .C2(new_n380), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT81), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n359), .B(new_n405), .ZN(new_n406));
  NOR4_X1   g0206(.A1(new_n372), .A2(new_n406), .A3(new_n319), .A4(new_n287), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(G169), .B2(new_n366), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n404), .B1(new_n385), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G238), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n290), .B(new_n411), .C1(new_n241), .C2(G1698), .ZN(new_n412));
  INV_X1    g0212(.A(new_n289), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n413), .C1(G107), .C2(new_n290), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n361), .C1(new_n218), .C2(new_n298), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g0217(.A(new_n417), .B(KEYINPUT73), .Z(new_n418));
  AND2_X1   g0218(.A1(new_n415), .A2(new_n305), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT8), .B(G58), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n274), .B1(new_n231), .B2(G77), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n271), .A2(G33), .ZN(new_n423));
  XOR2_X1   g0223(.A(KEYINPUT15), .B(G87), .Z(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n258), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n344), .A2(G77), .A3(new_n262), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n427), .B(new_n428), .C1(G77), .C2(new_n261), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n418), .A2(new_n419), .A3(new_n429), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n325), .A2(new_n387), .A3(new_n410), .A4(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n211), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n423), .B2(new_n217), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n308), .A2(new_n433), .ZN(new_n434));
  XOR2_X1   g0234(.A(new_n434), .B(KEYINPUT11), .Z(new_n435));
  NAND4_X1  g0235(.A1(new_n205), .A2(new_n211), .A3(G13), .A4(G20), .ZN(new_n436));
  XOR2_X1   g0236(.A(new_n436), .B(KEYINPUT12), .Z(new_n437));
  NAND3_X1  g0237(.A1(new_n344), .A2(G68), .A3(new_n262), .ZN(new_n438));
  XOR2_X1   g0238(.A(new_n438), .B(KEYINPUT77), .Z(new_n439));
  NOR3_X1   g0239(.A1(new_n435), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n361), .B1(new_n298), .B2(new_n212), .ZN(new_n442));
  OAI211_X1 g0242(.A(G226), .B(new_n293), .C1(new_n349), .C2(new_n334), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT75), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n290), .A2(KEYINPUT75), .A3(G226), .A4(new_n293), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G97), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n290), .A2(G232), .A3(G1698), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n445), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n442), .B1(new_n449), .B2(new_n413), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT13), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n441), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n445), .A2(new_n446), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n448), .A2(new_n447), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n413), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n442), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT13), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n441), .A3(KEYINPUT13), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(G200), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n450), .A2(new_n451), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n458), .A2(G190), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n440), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n459), .A2(G169), .A3(new_n460), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT14), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n459), .A2(KEYINPUT14), .A3(G169), .A4(new_n460), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n458), .A2(G179), .A3(new_n462), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT78), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT78), .ZN(new_n473));
  INV_X1    g0273(.A(new_n471), .ZN(new_n474));
  AOI211_X1 g0274(.A(new_n473), .B(new_n474), .C1(new_n468), .C2(new_n469), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n440), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n465), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n415), .A2(G179), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n415), .A2(new_n322), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n429), .A3(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n431), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n333), .A2(new_n335), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G250), .A3(new_n293), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT87), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G294), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n484), .A2(KEYINPUT87), .A3(G250), .A4(new_n293), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(G257), .A3(G1698), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G45), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n492), .A2(G1), .ZN(new_n493));
  AND2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NOR2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n289), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n491), .A2(new_n413), .B1(G264), .B2(new_n498), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n496), .A2(new_n286), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G200), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n205), .A2(G33), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n260), .A2(new_n261), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT24), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n507), .A2(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(KEYINPUT86), .ZN(new_n509));
  INV_X1    g0309(.A(G87), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n231), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT22), .B1(new_n511), .B2(new_n290), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n231), .A2(new_n513), .A3(new_n505), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT23), .A2(G107), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n345), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n206), .B1(new_n517), .B2(KEYINPUT23), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n484), .A2(new_n511), .A3(KEYINPUT22), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n509), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT22), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n271), .A2(G87), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n291), .ZN(new_n526));
  AND4_X1   g0326(.A1(new_n509), .A2(new_n523), .A3(new_n526), .A4(new_n521), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n508), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n506), .B1(new_n528), .B2(new_n258), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n499), .A2(G190), .A3(new_n500), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n261), .A2(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT25), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n502), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT85), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n484), .A2(G68), .A3(new_n271), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n271), .A2(G33), .A3(G97), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n271), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n535), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n258), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n424), .A2(new_n261), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n534), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AOI211_X1 g0347(.A(KEYINPUT85), .B(new_n545), .C1(new_n543), .C2(new_n258), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n547), .A2(new_n548), .B1(new_n425), .B2(new_n504), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n212), .A2(new_n293), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n218), .A2(G1698), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n484), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n517), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n289), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n493), .A2(G250), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n413), .B(new_n555), .C1(new_n286), .C2(new_n493), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n322), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n554), .A2(new_n556), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n319), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n549), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n558), .A2(new_n304), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(G190), .B2(new_n558), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n231), .B1(new_n333), .B2(new_n335), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n541), .B1(new_n563), .B2(G68), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n344), .B1(new_n564), .B2(new_n538), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT85), .B1(new_n565), .B2(new_n545), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n544), .A2(new_n534), .A3(new_n546), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n504), .A2(new_n510), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n562), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n533), .A2(new_n560), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G257), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n293), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n484), .B(new_n574), .C1(G264), .C2(new_n293), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n291), .A2(G303), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n289), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n500), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n497), .A2(new_n247), .ZN(new_n579));
  OR3_X1    g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n205), .A2(new_n516), .A3(G13), .A4(G20), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n344), .A2(G116), .A3(new_n261), .A4(new_n503), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n344), .B1(G20), .B2(new_n516), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G283), .ZN(new_n584));
  INV_X1    g0384(.A(G97), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n271), .B(new_n584), .C1(G33), .C2(new_n585), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n583), .A2(KEYINPUT20), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT20), .B1(new_n583), .B2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n581), .B(new_n582), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n580), .A2(G169), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR4_X1   g0392(.A1(new_n577), .A2(new_n319), .A3(new_n578), .A4(new_n579), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n589), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n580), .A2(KEYINPUT21), .A3(new_n589), .A4(G169), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n528), .A2(new_n258), .ZN(new_n597));
  INV_X1    g0397(.A(new_n506), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(new_n532), .ZN(new_n599));
  AOI21_X1  g0399(.A(G169), .B1(new_n499), .B2(new_n500), .ZN(new_n600));
  INV_X1    g0400(.A(new_n501), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n319), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n596), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n378), .A2(new_n585), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n504), .B2(new_n585), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n585), .A2(new_n505), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n202), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n608), .B2(KEYINPUT6), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n353), .A2(G107), .B1(new_n231), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n274), .A2(G77), .ZN(new_n611));
  XOR2_X1   g0411(.A(new_n611), .B(KEYINPUT82), .Z(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n605), .B1(new_n613), .B2(new_n258), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n500), .B1(new_n573), .B2(new_n497), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n218), .A2(G1698), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n616), .A2(KEYINPUT4), .B1(G250), .B2(G1698), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n617), .A2(new_n291), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT4), .ZN(new_n619));
  INV_X1    g0419(.A(new_n616), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n333), .B2(new_n335), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n621), .B2(KEYINPUT83), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n484), .A2(KEYINPUT83), .A3(new_n616), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n584), .B(new_n618), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n615), .B1(new_n624), .B2(new_n413), .ZN(new_n625));
  INV_X1    g0425(.A(G200), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n614), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI211_X1 g0427(.A(new_n416), .B(new_n615), .C1(new_n624), .C2(new_n413), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT84), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n624), .A2(new_n413), .ZN(new_n630));
  INV_X1    g0430(.A(new_n615), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n322), .ZN(new_n633));
  INV_X1    g0433(.A(new_n614), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n625), .A2(new_n319), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(G200), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n625), .A2(G190), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n614), .A4(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n629), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n589), .B1(new_n642), .B2(G190), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n626), .B2(new_n642), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n572), .A2(new_n603), .A3(new_n641), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n483), .A2(new_n645), .ZN(G372));
  INV_X1    g0446(.A(KEYINPUT90), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT89), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n568), .B2(new_n570), .ZN(new_n649));
  AOI211_X1 g0449(.A(KEYINPUT89), .B(new_n569), .C1(new_n566), .C2(new_n567), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n562), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n557), .A2(KEYINPUT88), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT88), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n653), .B(new_n322), .C1(new_n554), .C2(new_n556), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n549), .A2(new_n559), .A3(new_n652), .A4(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(new_n533), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n629), .A2(new_n640), .A3(new_n636), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n647), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n504), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n566), .A2(new_n567), .B1(new_n424), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n652), .A2(new_n654), .ZN(new_n661));
  INV_X1    g0461(.A(new_n559), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n570), .B1(new_n547), .B2(new_n548), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT89), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n568), .A2(new_n648), .A3(new_n570), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n663), .B1(new_n667), .B2(new_n562), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n641), .A2(new_n668), .A3(KEYINPUT90), .A4(new_n533), .ZN(new_n669));
  INV_X1    g0469(.A(new_n603), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n658), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n636), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n560), .A3(new_n571), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT26), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n651), .A2(new_n672), .A3(new_n675), .A4(new_n655), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n674), .A2(new_n676), .A3(new_n655), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n482), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n324), .ZN(new_n680));
  INV_X1    g0480(.A(new_n410), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n465), .A2(new_n481), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n476), .B2(new_n477), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n683), .B2(new_n387), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n680), .B1(new_n684), .B2(new_n318), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n679), .A2(new_n685), .ZN(G369));
  INV_X1    g0486(.A(G13), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n231), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n205), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT27), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT92), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT92), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n689), .A2(new_n693), .A3(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G213), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT91), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n689), .B2(KEYINPUT27), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n688), .A2(KEYINPUT91), .A3(new_n691), .A4(new_n205), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n589), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n596), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n596), .A2(new_n704), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n644), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT93), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n602), .A2(new_n599), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n703), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n599), .A2(new_n703), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n712), .A2(new_n533), .B1(new_n602), .B2(new_n599), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(G330), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n703), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n596), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n711), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n711), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n715), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n235), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n539), .A2(new_n516), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT94), .Z(new_n724));
  OR2_X1    g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n722), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n725), .A2(new_n205), .B1(new_n225), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n703), .B1(new_n671), .B2(new_n677), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n729), .A2(KEYINPUT29), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n651), .A2(new_n672), .A3(new_n655), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT26), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n732), .B(new_n655), .C1(KEYINPUT26), .C2(new_n673), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n603), .A2(new_n656), .A3(new_n657), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT29), .B(new_n716), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n499), .A2(new_n625), .A3(new_n593), .A4(new_n558), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n642), .A2(G179), .A3(new_n558), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(new_n501), .A3(new_n632), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n645), .B2(new_n703), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT95), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n741), .A2(new_n501), .A3(KEYINPUT95), .A4(new_n632), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n739), .A2(new_n747), .A3(new_n740), .A4(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT31), .B1(new_n749), .B2(new_n703), .ZN(new_n750));
  OAI21_X1  g0550(.A(G330), .B1(new_n745), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n736), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n728), .B1(new_n753), .B2(G1), .ZN(G364));
  AOI21_X1  g0554(.A(new_n227), .B1(G20), .B2(new_n322), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n304), .A2(G179), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(G20), .A3(G190), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT100), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G87), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n271), .A2(G190), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n756), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n762), .B(new_n290), .C1(new_n505), .C2(new_n764), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT101), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(G179), .A3(new_n626), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT97), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n767), .A2(KEYINPUT97), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n271), .A2(new_n319), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n771), .A2(G77), .B1(new_n269), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT98), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n773), .A2(new_n626), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n775), .A2(new_n776), .B1(new_n215), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT99), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n763), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G159), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n765), .A2(KEYINPUT101), .B1(new_n776), .B2(new_n775), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n781), .A2(G190), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n271), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n585), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n626), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n772), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n790), .B1(G68), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT102), .ZN(new_n795));
  AND4_X1   g0595(.A1(new_n766), .A2(new_n786), .A3(new_n787), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n789), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT103), .B(G326), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n797), .A2(G294), .B1(new_n777), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G329), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n782), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G322), .B2(new_n774), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n761), .A2(G303), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n291), .B1(new_n764), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(new_n793), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n802), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G311), .B2(new_n771), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n755), .B1(new_n796), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n721), .A2(new_n484), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n492), .B2(new_n226), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT96), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n492), .B2(new_n252), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n721), .A2(new_n291), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G355), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(G116), .C2(new_n235), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G13), .A2(G33), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(G20), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n755), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n205), .B1(new_n688), .B2(G45), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n722), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n707), .B2(new_n821), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n810), .A2(new_n823), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G330), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n708), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n826), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n709), .A2(G330), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n829), .B1(new_n833), .B2(new_n834), .ZN(G396));
  AND2_X1   g0635(.A1(new_n703), .A2(new_n429), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n430), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n481), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n481), .A2(new_n703), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n729), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(new_n751), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n827), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n755), .A2(new_n819), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n827), .B1(new_n217), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n839), .B1(new_n837), .B2(new_n481), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n761), .A2(G107), .B1(G303), .B2(new_n777), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n510), .B2(new_n764), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n790), .B(new_n849), .C1(G294), .C2(new_n774), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n290), .B1(new_n783), .B2(G311), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n771), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n852), .B1(new_n516), .B2(new_n853), .C1(new_n804), .C2(new_n792), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n764), .A2(new_n211), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n761), .B2(G50), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n783), .A2(G132), .ZN(new_n857));
  INV_X1    g0657(.A(new_n484), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n797), .B2(new_n269), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n774), .A2(G143), .B1(new_n793), .B2(G150), .ZN(new_n861));
  INV_X1    g0661(.A(G137), .ZN(new_n862));
  INV_X1    g0662(.A(G159), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n861), .B1(new_n862), .B2(new_n778), .C1(new_n853), .C2(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT34), .Z(new_n865));
  OAI21_X1  g0665(.A(new_n854), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT104), .ZN(new_n867));
  INV_X1    g0667(.A(new_n755), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n846), .B1(new_n820), .B2(new_n847), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n844), .A2(new_n869), .ZN(G384));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n477), .B(new_n703), .C1(new_n476), .C2(new_n465), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n470), .A2(new_n471), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n473), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n470), .A2(KEYINPUT78), .A3(new_n471), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n477), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n477), .A2(new_n703), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n464), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n749), .A2(new_n703), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT31), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(KEYINPUT107), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(KEYINPUT107), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n749), .A2(new_n703), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n882), .B(new_n884), .C1(new_n645), .C2(new_n703), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n879), .A2(new_n847), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n701), .A2(new_n388), .A3(new_n389), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n328), .B1(new_n340), .B2(new_n342), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n356), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n308), .A3(new_n343), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n887), .B1(new_n890), .B2(new_n381), .ZN(new_n891));
  INV_X1    g0691(.A(new_n382), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT105), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n382), .B(new_n895), .C1(new_n385), .C2(new_n887), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(KEYINPUT37), .C1(new_n891), .C2(new_n892), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n701), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n890), .A2(new_n381), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n900), .B(new_n901), .C1(new_n410), .C2(new_n387), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n899), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n871), .B1(new_n886), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n907));
  INV_X1    g0707(.A(new_n385), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n908), .B(new_n900), .C1(new_n410), .C2(new_n387), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n887), .A2(new_n385), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n892), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n896), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n871), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n841), .B1(new_n872), .B2(new_n878), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(new_n885), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n906), .A2(G330), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n482), .A2(G330), .A3(new_n885), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT108), .Z(new_n922));
  NAND2_X1  g0722(.A1(new_n899), .A2(new_n902), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n914), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n907), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n917), .A3(new_n885), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n879), .A2(new_n847), .A3(new_n885), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n871), .A2(new_n926), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n482), .A3(new_n885), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n730), .A2(new_n482), .A3(new_n735), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n931), .A2(new_n685), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n907), .A2(new_n915), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT106), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT39), .B1(new_n903), .B2(new_n904), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT106), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n907), .A2(new_n915), .A3(new_n938), .A4(new_n934), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n876), .A2(new_n703), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n678), .A2(new_n716), .A3(new_n847), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n840), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n925), .A3(new_n879), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n681), .A2(new_n900), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n942), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n933), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n205), .B2(new_n688), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n228), .B(new_n231), .C1(new_n609), .C2(KEYINPUT35), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n516), .B(new_n951), .C1(KEYINPUT35), .C2(new_n609), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT36), .Z(new_n953));
  AOI211_X1 g0753(.A(new_n217), .B(new_n225), .C1(new_n269), .C2(G68), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n211), .A2(G50), .ZN(new_n955));
  OAI211_X1 g0755(.A(G1), .B(new_n687), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n950), .A2(new_n953), .A3(new_n956), .ZN(G367));
  INV_X1    g0757(.A(new_n667), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n703), .ZN(new_n959));
  MUX2_X1   g0759(.A(new_n663), .B(new_n668), .S(new_n959), .Z(new_n960));
  INV_X1    g0760(.A(KEYINPUT109), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n960), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n821), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n792), .A2(new_n863), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n771), .A2(G50), .B1(G68), .B2(new_n797), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n782), .A2(new_n862), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n764), .A2(new_n217), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(G143), .C2(new_n777), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n761), .A2(new_n269), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n967), .A2(new_n290), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n966), .B(new_n972), .C1(G150), .C2(new_n774), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n783), .A2(G317), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n771), .A2(G283), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n793), .A2(G294), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G303), .A2(new_n774), .B1(new_n777), .B2(G311), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n484), .B1(new_n797), .B2(G107), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n761), .A2(KEYINPUT46), .A3(G116), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n585), .B2(new_n764), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT46), .B1(new_n761), .B2(G116), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n973), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT47), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n755), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n822), .B1(new_n235), .B2(new_n425), .C1(new_n812), .C2(new_n248), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n965), .A2(new_n986), .A3(new_n826), .A4(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT113), .Z(new_n989));
  NOR2_X1   g0789(.A1(new_n963), .A2(new_n964), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n641), .B1(new_n614), .B2(new_n716), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n672), .A2(new_n703), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT112), .B1(new_n715), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT112), .ZN(new_n996));
  INV_X1    g0796(.A(new_n994), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n831), .A2(new_n996), .A3(new_n714), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n991), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n995), .A2(new_n991), .A3(new_n998), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT42), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n997), .A2(KEYINPUT110), .A3(new_n718), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT110), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n718), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n1006), .B2(new_n994), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1003), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n992), .A2(new_n710), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n703), .B1(new_n1010), .B2(new_n636), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(KEYINPUT111), .A3(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1004), .A2(new_n1007), .A3(new_n1003), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT111), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1002), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n1000), .A3(new_n1018), .A4(new_n1001), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n719), .A2(new_n997), .A3(KEYINPUT44), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT44), .B1(new_n719), .B2(new_n997), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT45), .B1(new_n719), .B2(new_n997), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT45), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n994), .A2(new_n718), .A3(new_n1027), .A4(new_n711), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n831), .B(new_n714), .C1(new_n1025), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1029), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1031), .A2(new_n715), .A3(new_n1024), .A4(new_n1023), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n714), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n717), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n1006), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n831), .B(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n753), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n722), .B(KEYINPUT41), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n825), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n989), .B1(new_n1022), .B2(new_n1041), .ZN(G387));
  AOI21_X1  g0842(.A(new_n812), .B1(new_n244), .B2(G45), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n724), .B2(new_n816), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n421), .A2(new_n215), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n211), .A2(new_n217), .ZN(new_n1047));
  NOR4_X1   g0847(.A1(new_n1046), .A2(new_n724), .A3(G45), .A4(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1044), .A2(new_n1048), .B1(G107), .B2(new_n235), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n827), .B1(new_n1049), .B2(new_n822), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT114), .Z(new_n1051));
  AOI22_X1  g0851(.A1(new_n777), .A2(G322), .B1(new_n793), .B2(G311), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT116), .Z(new_n1053));
  AOI22_X1  g0853(.A1(new_n771), .A2(G303), .B1(G317), .B2(new_n774), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT48), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n761), .ZN(new_n1057));
  INV_X1    g0857(.A(G294), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1057), .A2(new_n1058), .B1(new_n789), .B2(new_n804), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1056), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  XOR2_X1   g0862(.A(KEYINPUT117), .B(KEYINPUT49), .Z(new_n1063));
  XNOR2_X1  g0863(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n783), .A2(new_n798), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n764), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n484), .B1(new_n1066), .B2(G116), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n377), .A2(new_n792), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n761), .A2(G77), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n853), .B2(new_n211), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(G97), .C2(new_n1066), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n797), .A2(new_n424), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n774), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1073), .B1(new_n215), .B2(new_n1074), .C1(new_n863), .C2(new_n778), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G150), .B2(new_n783), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1072), .A2(new_n484), .A3(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1068), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1051), .B1(new_n1078), .B2(new_n868), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1079), .A2(KEYINPUT118), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1034), .A2(new_n821), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1079), .A2(KEYINPUT118), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n722), .B1(new_n753), .B2(new_n1037), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n753), .A2(new_n1037), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1083), .B1(new_n824), .B2(new_n1038), .C1(new_n1084), .C2(new_n1086), .ZN(G393));
  NAND3_X1  g0887(.A1(new_n1030), .A2(new_n1032), .A3(new_n825), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G311), .A2(new_n774), .B1(new_n777), .B2(G317), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT52), .Z(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n505), .B2(new_n764), .C1(new_n804), .C2(new_n1057), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G294), .B2(new_n771), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n793), .A2(G303), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n797), .A2(G116), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n290), .B1(new_n783), .B2(G322), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT119), .Z(new_n1097));
  OAI22_X1  g0897(.A1(new_n789), .A2(new_n217), .B1(new_n215), .B2(new_n792), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n858), .B1(new_n783), .B2(G143), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n510), .B2(new_n764), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(new_n421), .C2(new_n771), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G150), .A2(new_n777), .B1(new_n774), .B2(G159), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G68), .B2(new_n761), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n755), .B1(new_n1097), .B2(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n822), .B1(new_n585), .B2(new_n235), .C1(new_n812), .C2(new_n255), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n827), .B1(new_n994), .B2(new_n821), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1088), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1033), .A2(new_n1085), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n722), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1033), .A2(new_n1085), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(G390));
  OAI21_X1  g0915(.A(new_n716), .B1(new_n733), .B2(new_n734), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n838), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n840), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n879), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n907), .A2(new_n915), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n941), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n879), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1125), .A2(new_n751), .A3(new_n841), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n941), .B1(new_n944), .B2(new_n879), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1124), .B(new_n1126), .C1(new_n1127), .C2(new_n940), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1122), .B1(new_n1118), .B2(new_n879), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n839), .B1(new_n729), .B2(new_n847), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1121), .B1(new_n1131), .B2(new_n1125), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n885), .A2(G330), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n1125), .A2(new_n1134), .A3(new_n841), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1128), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n931), .A2(new_n920), .A3(new_n685), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n751), .A2(new_n841), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1138), .A2(new_n879), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n944), .B1(new_n1139), .B2(new_n1135), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n879), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1118), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1125), .B1(new_n1134), .B2(new_n841), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1137), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n726), .B1(new_n1136), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n1136), .B2(new_n1145), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1130), .A2(new_n819), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n761), .A2(G150), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n291), .B(new_n1151), .C1(G132), .C2(new_n774), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n783), .A2(G125), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n777), .A2(G128), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n789), .A2(new_n863), .B1(new_n862), .B2(new_n792), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT54), .B(G143), .Z(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n771), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT120), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G50), .B2(new_n1066), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1159), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n762), .B1(new_n516), .B2(new_n1074), .C1(new_n804), .C2(new_n778), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n789), .A2(new_n217), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n291), .B1(new_n782), .B2(new_n1058), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1161), .A2(new_n855), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n585), .B2(new_n853), .C1(new_n505), .C2(new_n792), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n868), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n827), .B(new_n1166), .C1(new_n377), .C2(new_n845), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1136), .A2(new_n825), .B1(new_n1148), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1147), .A2(new_n1168), .ZN(G378));
  XOR2_X1   g0969(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1170));
  XNOR2_X1  g0970(.A(new_n325), .B(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n313), .A2(new_n900), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n928), .B2(G330), .ZN(new_n1174));
  AND4_X1   g0974(.A1(G330), .A2(new_n906), .A3(new_n918), .A4(new_n1173), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1174), .A2(new_n1175), .A3(new_n948), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1173), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n919), .A2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n906), .A2(new_n1173), .A3(G330), .A4(new_n918), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n946), .B1(new_n940), .B2(new_n941), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1178), .A2(new_n1179), .B1(new_n945), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1136), .A2(new_n1145), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1137), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1185), .A3(KEYINPUT57), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT57), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n948), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1178), .A2(new_n945), .A3(new_n1180), .A4(new_n1179), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1137), .B1(new_n1136), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1187), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1186), .A2(new_n1193), .A3(new_n722), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n853), .A2(new_n425), .B1(new_n211), .B2(new_n789), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n783), .A2(G283), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1066), .A2(new_n269), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n484), .A2(G41), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1070), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT122), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1195), .B(new_n1200), .C1(G97), .C2(new_n793), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n505), .B2(new_n1074), .C1(new_n516), .C2(new_n778), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT58), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n215), .B1(new_n369), .B2(G41), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n771), .A2(G137), .B1(G128), .B2(new_n774), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n761), .A2(new_n1156), .B1(G132), .B2(new_n793), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n797), .A2(G150), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n777), .A2(G125), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(G33), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1066), .A2(G159), .ZN(new_n1213));
  AOI21_X1  g1013(.A(G41), .B1(new_n783), .B2(G124), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1203), .A2(new_n1204), .A3(new_n1215), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1216), .A2(new_n755), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n827), .B(new_n1217), .C1(new_n215), .C2(new_n845), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1173), .A2(new_n819), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n825), .A2(new_n1182), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1194), .A2(new_n1220), .ZN(G375));
  INV_X1    g1021(.A(new_n1145), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1140), .A2(new_n1137), .A3(new_n1144), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1040), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1125), .A2(new_n819), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n783), .A2(G128), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1197), .B(new_n1226), .C1(new_n789), .C2(new_n215), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1057), .A2(new_n863), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(G150), .C2(new_n771), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n774), .A2(G137), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n793), .A2(new_n1156), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n858), .B1(new_n777), .B2(G132), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1073), .B1(new_n804), .B2(new_n1074), .C1(new_n1058), .C2(new_n778), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G107), .B2(new_n771), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n783), .A2(G303), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n761), .A2(G97), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n290), .B(new_n969), .C1(G116), .C2(new_n793), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n868), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n827), .B(new_n1240), .C1(new_n211), .C2(new_n845), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1191), .A2(new_n825), .B1(new_n1225), .B2(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1224), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G381));
  NOR2_X1   g1044(.A1(G375), .A2(G378), .ZN(new_n1245));
  INV_X1    g1045(.A(G384), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(new_n1247), .A2(G387), .A3(G396), .A4(G393), .ZN(new_n1248));
  INV_X1    g1048(.A(G390), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1245), .A2(new_n1248), .A3(new_n1249), .ZN(G407));
  AOI21_X1  g1050(.A(new_n696), .B1(new_n1245), .B2(new_n702), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(G407), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT123), .ZN(G409));
  XOR2_X1   g1053(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1254));
  NOR2_X1   g1054(.A1(new_n696), .A2(G343), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G375), .B2(G378), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT124), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT124), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1188), .A2(new_n1258), .A3(new_n1189), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n825), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT125), .ZN(new_n1263));
  INV_X1    g1063(.A(G378), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT125), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1260), .A2(new_n1265), .A3(new_n1261), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1182), .A2(new_n1185), .A3(new_n1040), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1256), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1255), .A2(G2897), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1223), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1223), .A2(new_n1272), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n722), .A3(new_n1222), .A4(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(G384), .A3(new_n1242), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1275), .B2(new_n1242), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1271), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1278), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(new_n1276), .A3(new_n1270), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1254), .B1(new_n1269), .B2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1256), .A2(new_n1268), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT62), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1256), .A2(new_n1268), .A3(new_n1287), .A4(new_n1284), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1283), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(new_n1249), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G390), .B(new_n989), .C1(new_n1041), .C2(new_n1022), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1291), .A2(KEYINPUT126), .ZN(new_n1293));
  INV_X1    g1093(.A(G396), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(G393), .B(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1292), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(G393), .B(G396), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1291), .A4(new_n1290), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1289), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(new_n1256), .B2(new_n1268), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1285), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1256), .A2(new_n1268), .A3(KEYINPUT63), .A4(new_n1284), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1307), .A2(new_n1300), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1302), .A2(new_n1310), .ZN(G405));
  XNOR2_X1  g1111(.A(G375), .B(new_n1264), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1300), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1300), .A2(new_n1312), .ZN(new_n1315));
  OAI22_X1  g1115(.A1(new_n1314), .A2(new_n1315), .B1(new_n1278), .B2(new_n1277), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1315), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(new_n1284), .A3(new_n1313), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(G402));
endmodule


