//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT80), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n190), .A2(new_n192), .A3(G128), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT64), .B1(new_n191), .B2(G146), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(new_n189), .A3(G143), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(new_n192), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT0), .B(G128), .Z(new_n198));
  AOI22_X1  g012(.A1(KEYINPUT0), .A2(new_n193), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT79), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n190), .A2(new_n192), .A3(new_n204), .A4(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT65), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n207), .A2(new_n208), .A3(new_n204), .A4(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G128), .ZN(new_n211));
  AOI22_X1  g025(.A1(new_n206), .A2(new_n209), .B1(new_n197), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n203), .B1(new_n212), .B2(new_n200), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n202), .B1(new_n213), .B2(new_n201), .ZN(new_n214));
  INV_X1    g028(.A(G224), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G953), .ZN(new_n216));
  XOR2_X1   g030(.A(new_n214), .B(new_n216), .Z(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G104), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G107), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n221), .B2(G107), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n219), .A3(G104), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n225), .A2(new_n227), .A3(new_n218), .A4(new_n222), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT74), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n224), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT76), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n219), .A2(G104), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(KEYINPUT3), .B2(new_n220), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n235), .A2(KEYINPUT74), .A3(new_n218), .A4(new_n227), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n228), .A2(new_n229), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n223), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT76), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G116), .B(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT5), .ZN(new_n242));
  INV_X1    g056(.A(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G116), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n242), .B(G113), .C1(KEYINPUT5), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT2), .ZN(new_n246));
  INV_X1    g060(.A(G113), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT66), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT2), .A3(G113), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n247), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(new_n241), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n245), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n233), .A2(new_n240), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n225), .A2(new_n227), .A3(new_n222), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT75), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(G101), .ZN(new_n261));
  OAI211_X1 g075(.A(KEYINPUT4), .B(new_n261), .C1(new_n230), .C2(new_n231), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n251), .A2(new_n252), .ZN(new_n263));
  INV_X1    g077(.A(new_n241), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n253), .A3(KEYINPUT67), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n251), .A2(new_n252), .A3(new_n241), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n241), .B1(new_n251), .B2(new_n252), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n260), .A2(new_n262), .A3(new_n266), .A4(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT78), .B1(new_n256), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  XOR2_X1   g087(.A(G110), .B(G122), .Z(new_n274));
  NAND3_X1  g088(.A1(new_n256), .A2(KEYINPUT78), .A3(new_n271), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n274), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n256), .A2(new_n271), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT6), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n273), .A2(KEYINPUT6), .A3(new_n274), .A4(new_n275), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n217), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n232), .A2(new_n254), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n256), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n274), .B(KEYINPUT8), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n278), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT7), .B1(new_n215), .B2(G953), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n214), .B(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n283), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n188), .B1(new_n282), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n256), .A2(KEYINPUT78), .A3(new_n271), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n292), .A2(new_n272), .A3(new_n277), .ZN(new_n293));
  INV_X1    g107(.A(new_n279), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n281), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n217), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n290), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n188), .A2(KEYINPUT81), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n187), .ZN(new_n301));
  AOI211_X1 g115(.A(new_n301), .B(new_n290), .C1(new_n295), .C2(new_n296), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT81), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n291), .B(new_n300), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  OR2_X1    g119(.A1(KEYINPUT97), .A2(G952), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT97), .A2(G952), .ZN(new_n307));
  AOI21_X1  g121(.A(G953), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G234), .ZN(new_n309));
  INV_X1    g123(.A(G237), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G953), .ZN(new_n312));
  AOI211_X1 g126(.A(new_n283), .B(new_n312), .C1(G234), .C2(G237), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT21), .B(G898), .Z(new_n315));
  OAI21_X1  g129(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n304), .A2(new_n305), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G472), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n270), .A2(new_n266), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT11), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(G137), .ZN(new_n324));
  INV_X1    g138(.A(G137), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT11), .A3(G134), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(G137), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G131), .ZN(new_n329));
  INV_X1    g143(.A(G131), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n324), .A2(new_n326), .A3(new_n330), .A4(new_n327), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n199), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n327), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n323), .A2(G137), .ZN(new_n335));
  OAI21_X1  g149(.A(G131), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n331), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n333), .B1(new_n212), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n320), .B1(new_n321), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(G237), .A2(G953), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G210), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(G101), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n344), .A2(KEYINPUT29), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n206), .A2(new_n209), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n211), .A2(new_n197), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n337), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n348), .A2(new_n349), .B1(new_n332), .B2(new_n199), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n270), .A2(new_n266), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT68), .B1(new_n321), .B2(new_n338), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT68), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n352), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n339), .B(new_n345), .C1(new_n356), .C2(new_n320), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT70), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n357), .A2(new_n358), .A3(new_n283), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n357), .B2(new_n283), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n344), .B(KEYINPUT69), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n363), .B(new_n339), .C1(new_n356), .C2(new_n320), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT30), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n199), .A2(new_n332), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n337), .B1(new_n346), .B2(new_n347), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n333), .B(KEYINPUT30), .C1(new_n212), .C2(new_n337), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n321), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n355), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n354), .B1(new_n350), .B2(new_n351), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n344), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT29), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n364), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n319), .B1(new_n361), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT32), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n339), .B1(new_n356), .B2(new_n320), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n344), .B(new_n370), .C1(new_n371), .C2(new_n372), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT31), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n353), .A2(new_n355), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n384), .A2(KEYINPUT31), .A3(new_n344), .A4(new_n370), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n380), .A2(new_n362), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(G472), .A2(G902), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n379), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n362), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n383), .A2(new_n385), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT32), .A3(new_n387), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n378), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n397));
  OR3_X1    g211(.A1(new_n200), .A2(KEYINPUT16), .A3(G140), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(G146), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n189), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT24), .B(G110), .Z(new_n401));
  NOR2_X1   g215(.A1(new_n243), .A2(G128), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n243), .A2(G128), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT71), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT71), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n401), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G110), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n402), .A2(KEYINPUT23), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n404), .A2(KEYINPUT23), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n410), .B(new_n411), .C1(new_n412), .C2(new_n402), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n399), .B(new_n400), .C1(new_n409), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(new_n408), .A3(new_n401), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n411), .B1(new_n412), .B2(new_n402), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G110), .ZN(new_n418));
  INV_X1    g232(.A(new_n399), .ZN(new_n419));
  AOI21_X1  g233(.A(G146), .B1(new_n397), .B2(new_n398), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n416), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT22), .B(G137), .ZN(new_n423));
  INV_X1    g237(.A(G221), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n424), .A2(new_n309), .A3(G953), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n423), .B(new_n425), .Z(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n415), .A2(new_n421), .A3(new_n426), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT72), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT25), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n432), .A2(KEYINPUT25), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n431), .A2(new_n283), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G217), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(G234), .B2(new_n283), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n432), .B(KEYINPUT25), .C1(new_n430), .C2(G902), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n437), .A2(G902), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n431), .A2(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n395), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n340), .A2(G143), .A3(G214), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT84), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n447));
  AND4_X1   g261(.A1(KEYINPUT82), .A2(new_n310), .A3(new_n312), .A4(G214), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT82), .B1(new_n340), .B2(G214), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(new_n450), .B2(new_n191), .ZN(new_n451));
  NOR4_X1   g265(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT83), .A4(G143), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G131), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT17), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n446), .B(new_n330), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n419), .A2(new_n420), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(KEYINPUT17), .A3(G131), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT85), .B(G104), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n445), .B(KEYINPUT84), .Z(new_n464));
  NAND3_X1  g278(.A1(new_n450), .A2(new_n447), .A3(new_n191), .ZN(new_n465));
  INV_X1    g279(.A(new_n449), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n340), .A2(KEYINPUT82), .A3(G214), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n191), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT83), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT18), .A2(G131), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n396), .A2(new_n189), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n470), .A2(new_n471), .B1(new_n400), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n453), .A2(KEYINPUT18), .A3(G131), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n460), .A2(new_n463), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n460), .A2(new_n475), .A3(new_n478), .A4(new_n463), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n454), .A2(new_n456), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n396), .B(KEYINPUT19), .Z(new_n482));
  OAI21_X1  g296(.A(new_n399), .B1(new_n482), .B2(G146), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n481), .A2(new_n484), .B1(new_n473), .B2(new_n474), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT86), .B1(new_n485), .B2(new_n463), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n487));
  INV_X1    g301(.A(new_n463), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n473), .A2(new_n474), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n483), .B1(new_n454), .B2(new_n456), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n480), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G475), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT20), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(KEYINPUT88), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n493), .A2(new_n494), .A3(new_n283), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n463), .B1(new_n460), .B2(new_n475), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n477), .B2(new_n479), .ZN(new_n499));
  OAI21_X1  g313(.A(G475), .B1(new_n499), .B2(G902), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n477), .A2(new_n479), .B1(new_n486), .B2(new_n491), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n501), .A2(G475), .A3(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n496), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n495), .A2(KEYINPUT88), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n497), .B(new_n500), .C1(new_n502), .C2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  NOR2_X1   g321(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT94), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT9), .B(G234), .Z(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n514), .A2(new_n436), .A3(G953), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT90), .B1(new_n191), .B2(G128), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n518));
  INV_X1    g332(.A(G128), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n519), .A3(G143), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n191), .A2(G128), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n191), .A2(KEYINPUT13), .A3(G128), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G134), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT91), .ZN(new_n528));
  INV_X1    g342(.A(G116), .ZN(new_n529));
  OR2_X1    g343(.A1(KEYINPUT89), .A2(G122), .ZN(new_n530));
  NAND2_X1  g344(.A1(KEYINPUT89), .A2(G122), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(G122), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n219), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n534), .ZN(new_n536));
  OAI21_X1  g350(.A(G107), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n526), .A2(new_n539), .A3(G134), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n528), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n521), .A2(new_n323), .A3(new_n522), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n521), .A2(new_n544), .A3(new_n323), .A4(new_n522), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n532), .A2(new_n536), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n219), .A2(KEYINPUT14), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT14), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n532), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n551), .B1(new_n553), .B2(new_n537), .ZN(new_n554));
  INV_X1    g368(.A(new_n542), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n323), .B1(new_n521), .B2(new_n522), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT93), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n556), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n542), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n554), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n516), .B1(new_n547), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n560), .ZN(new_n563));
  INV_X1    g377(.A(new_n554), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n546), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n566), .A2(new_n528), .A3(new_n540), .A4(new_n538), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n567), .A3(new_n515), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n512), .B1(new_n569), .B2(new_n283), .ZN(new_n570));
  AOI211_X1 g384(.A(KEYINPUT94), .B(G902), .C1(new_n562), .C2(new_n568), .ZN(new_n571));
  OAI211_X1 g385(.A(KEYINPUT96), .B(new_n511), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n511), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n547), .A2(new_n561), .A3(new_n516), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n515), .B1(new_n565), .B2(new_n567), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT94), .B1(new_n576), .B2(G902), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n569), .A2(new_n512), .A3(new_n283), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n576), .A2(G902), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n573), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n572), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n506), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n348), .B1(new_n233), .B2(new_n240), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n207), .B1(G128), .B2(new_n210), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n209), .B2(new_n206), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n232), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n332), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT12), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT12), .B(new_n332), .C1(new_n585), .C2(new_n588), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(KEYINPUT77), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n233), .A2(new_n240), .A3(KEYINPUT10), .A4(new_n348), .ZN(new_n594));
  INV_X1    g408(.A(new_n332), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n260), .A2(new_n262), .A3(new_n199), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n232), .B2(new_n587), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(G110), .B(G140), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n312), .A2(G227), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT77), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n589), .A2(new_n603), .A3(new_n590), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n593), .A2(new_n599), .A3(new_n602), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n594), .A2(new_n596), .A3(new_n598), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n332), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n599), .ZN(new_n608));
  INV_X1    g422(.A(new_n602), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G469), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n612), .A3(new_n283), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n283), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n593), .A2(new_n599), .A3(new_n604), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n602), .B(KEYINPUT73), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n607), .A2(new_n599), .A3(new_n602), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(G469), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n613), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n424), .B1(new_n513), .B2(new_n283), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n318), .A2(new_n444), .A3(new_n584), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  AOI21_X1  g441(.A(new_n319), .B1(new_n392), .B2(new_n283), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n386), .A2(new_n388), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND4_X1   g444(.A1(new_n442), .A2(new_n621), .A3(new_n623), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n576), .A2(KEYINPUT33), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n569), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(G478), .A3(new_n283), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n507), .B1(new_n570), .B2(new_n571), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n635), .A2(KEYINPUT98), .A3(G478), .A4(new_n283), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n506), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n305), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n301), .B1(new_n282), .B2(new_n290), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n297), .A2(new_n187), .A3(new_n298), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n647), .A2(new_n316), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n631), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT34), .B(G104), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  NAND3_X1  g465(.A1(new_n493), .A2(new_n494), .A3(new_n283), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n504), .A3(new_n503), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n500), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g469(.A(KEYINPUT99), .B(G475), .C1(new_n499), .C2(G902), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n653), .A2(new_n497), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n583), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n631), .A2(new_n659), .A3(new_n648), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n317), .A2(new_n624), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n427), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n422), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n440), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n439), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT100), .B1(new_n630), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n667), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n670));
  NOR4_X1   g484(.A1(new_n628), .A2(new_n669), .A3(new_n629), .A4(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n663), .A2(new_n584), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NOR3_X1   g489(.A1(new_n359), .A2(new_n376), .A3(new_n360), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n389), .B(new_n393), .C1(new_n676), .C2(new_n319), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n677), .A2(new_n623), .A3(new_n621), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n655), .A2(new_n656), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n497), .B1(new_n502), .B2(new_n505), .ZN(new_n680));
  INV_X1    g494(.A(new_n311), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n681), .B1(new_n682), .B2(new_n313), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n647), .A2(new_n667), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n678), .A2(new_n583), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  XNOR2_X1  g502(.A(new_n683), .B(KEYINPUT39), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n621), .A2(new_n623), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n644), .B1(new_n691), .B2(KEYINPUT40), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n381), .B1(new_n363), .B2(new_n356), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n283), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G472), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n389), .A2(new_n393), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n667), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n506), .A2(new_n583), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT38), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n304), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n297), .A2(new_n298), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n646), .A2(KEYINPUT81), .B1(new_n704), .B2(new_n188), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(KEYINPUT38), .A3(new_n300), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT40), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n621), .A2(new_n707), .A3(new_n623), .A4(new_n690), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n701), .A2(new_n703), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n699), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n191), .ZN(G45));
  INV_X1    g525(.A(new_n683), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n506), .A2(new_n641), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n678), .A2(new_n686), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  NAND2_X1  g529(.A1(new_n611), .A2(new_n283), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n612), .A2(KEYINPUT101), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n611), .B(new_n283), .C1(KEYINPUT101), .C2(new_n612), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n623), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n444), .A2(new_n643), .A3(new_n648), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND2_X1  g538(.A1(new_n645), .A2(new_n646), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n305), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n720), .A2(new_n395), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(new_n442), .A3(new_n316), .A4(new_n659), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G116), .ZN(G18));
  NAND4_X1  g543(.A1(new_n727), .A2(new_n584), .A3(new_n316), .A4(new_n667), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n380), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(KEYINPUT102), .B(new_n339), .C1(new_n356), .C2(new_n320), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n362), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n388), .B1(new_n735), .B2(new_n391), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n628), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n442), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n720), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n506), .A2(new_n741), .A3(new_n583), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n741), .B1(new_n506), .B2(new_n583), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n740), .B(new_n648), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n700), .A2(KEYINPUT103), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n506), .A2(new_n741), .A3(new_n583), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n648), .A4(new_n740), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  NOR3_X1   g566(.A1(new_n736), .A2(new_n628), .A3(new_n669), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n506), .A2(new_n753), .A3(new_n641), .A4(new_n712), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n720), .A2(new_n726), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(KEYINPUT42), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n619), .A2(KEYINPUT105), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n607), .A2(new_n762), .A3(new_n599), .A4(new_n602), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n618), .A2(G469), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n613), .A2(new_n615), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n623), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n304), .B2(new_n644), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n705), .A2(KEYINPUT107), .A3(new_n305), .A4(new_n300), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n766), .A2(KEYINPUT106), .A3(new_n623), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n769), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n444), .ZN(new_n775));
  INV_X1    g589(.A(new_n713), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n758), .A2(KEYINPUT42), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n760), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n771), .A2(new_n772), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n766), .A2(KEYINPUT106), .A3(new_n623), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT106), .B1(new_n766), .B2(new_n623), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n781), .A2(new_n784), .A3(new_n444), .A4(new_n713), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n759), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n780), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G131), .ZN(G33));
  NOR3_X1   g602(.A1(new_n657), .A2(new_n658), .A3(new_n683), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n781), .A2(new_n784), .A3(new_n444), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  INV_X1    g605(.A(new_n781), .ZN(new_n792));
  INV_X1    g606(.A(new_n641), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT43), .B1(new_n793), .B2(new_n506), .ZN(new_n794));
  INV_X1    g608(.A(new_n680), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT43), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n500), .A4(new_n641), .ZN(new_n797));
  INV_X1    g611(.A(new_n630), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n794), .A2(new_n797), .A3(new_n798), .A4(new_n667), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n799), .A2(KEYINPUT110), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT110), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n792), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n800), .ZN(new_n804));
  INV_X1    g618(.A(new_n613), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n618), .A2(KEYINPUT45), .A3(new_n764), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(G469), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT45), .B1(new_n618), .B2(new_n619), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT109), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n616), .A2(new_n617), .B1(new_n761), .B2(new_n763), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n612), .B1(new_n810), .B2(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n618), .A2(new_n619), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n614), .B1(new_n809), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n805), .B1(new_n817), .B2(KEYINPUT46), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n807), .A2(KEYINPUT109), .A3(new_n808), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n815), .B1(new_n811), .B2(new_n814), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n615), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT46), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n622), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n803), .A2(new_n690), .A3(new_n804), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G137), .ZN(G39));
  INV_X1    g640(.A(KEYINPUT47), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  AOI211_X1 g642(.A(KEYINPUT47), .B(new_n622), .C1(new_n818), .C2(new_n823), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n792), .A2(new_n677), .A3(new_n442), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(KEYINPUT111), .A3(new_n713), .A4(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n613), .B1(new_n821), .B2(new_n822), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n817), .A2(KEYINPUT46), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n623), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT47), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n824), .A2(new_n827), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n713), .A4(new_n831), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n751), .A2(new_n722), .A3(new_n728), .A4(new_n730), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n684), .A2(new_n771), .A3(new_n772), .A4(new_n667), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n583), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n678), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT113), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n677), .A2(new_n848), .A3(new_n623), .A4(new_n621), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n657), .A2(new_n669), .A3(new_n683), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n781), .A2(new_n851), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n781), .A2(new_n784), .A3(new_n754), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n663), .B(new_n584), .C1(new_n444), .C2(new_n672), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n642), .B1(new_n848), .B2(new_n506), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n318), .A3(new_n631), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n790), .A2(new_n856), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n696), .A2(new_n669), .A3(new_n712), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n767), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n863), .B(new_n647), .C1(new_n742), .C2(new_n743), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n687), .A3(new_n714), .A4(new_n756), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n624), .A2(new_n685), .A3(new_n395), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n868), .A2(new_n789), .B1(new_n754), .B2(new_n755), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT52), .A3(new_n714), .A4(new_n864), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n845), .A2(new_n861), .A3(new_n787), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n873));
  INV_X1    g687(.A(new_n860), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n850), .A2(new_n854), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n871), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n872), .A2(KEYINPUT53), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n872), .B1(KEYINPUT53), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n843), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n794), .A2(new_n797), .A3(new_n681), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n739), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n755), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT116), .ZN(new_n884));
  NAND2_X1  g698(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n308), .A3(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n792), .A2(new_n720), .A3(new_n881), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT48), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n887), .B(new_n444), .C1(KEYINPUT117), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(KEYINPUT48), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n887), .A2(KEYINPUT117), .A3(new_n888), .A4(new_n444), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n792), .A2(new_n696), .A3(new_n720), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n442), .A3(new_n681), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(new_n642), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n867), .A2(new_n870), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n673), .A2(new_n859), .A3(new_n626), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n875), .A2(new_n898), .A3(new_n790), .A4(new_n856), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n897), .A2(new_n899), .A3(new_n844), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n787), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n872), .A2(KEYINPUT53), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(KEYINPUT54), .A3(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n880), .A2(new_n893), .A3(new_n896), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n718), .A2(new_n719), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(new_n623), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n781), .B(new_n882), .C1(new_n830), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n706), .A2(new_n703), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n882), .A2(new_n644), .A3(new_n909), .A4(new_n721), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT50), .Z(new_n911));
  OR3_X1    g725(.A1(new_n895), .A2(new_n506), .A3(new_n641), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n887), .A2(new_n753), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n908), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n905), .A2(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n506), .B(new_n793), .C1(new_n706), .C2(new_n703), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n305), .A3(new_n697), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n906), .A2(KEYINPUT49), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n906), .A2(KEYINPUT49), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(new_n442), .A3(new_n623), .A4(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n917), .B1(new_n919), .B2(new_n922), .ZN(G75));
  NAND2_X1  g737(.A1(new_n876), .A2(KEYINPUT53), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n787), .A3(new_n900), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(G210), .A3(G902), .A4(new_n877), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n295), .A2(new_n296), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(new_n282), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n929), .B(new_n930), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n926), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n926), .B2(new_n927), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n312), .A2(G952), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(G51));
  XOR2_X1   g750(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n614), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n937), .A2(new_n614), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n925), .A2(KEYINPUT54), .A3(new_n877), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT54), .B1(new_n925), .B2(new_n877), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n611), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n878), .A2(new_n879), .A3(new_n283), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n816), .A3(new_n809), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n935), .B1(new_n943), .B2(new_n945), .ZN(G54));
  NAND3_X1  g760(.A1(new_n944), .A2(KEYINPUT58), .A3(G475), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n501), .ZN(new_n948));
  INV_X1    g762(.A(new_n935), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n944), .A2(KEYINPUT58), .A3(G475), .A4(new_n493), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(G60));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT59), .Z(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n635), .B(new_n954), .C1(new_n940), .C2(new_n941), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n949), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT120), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n953), .B1(new_n880), .B2(new_n904), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(new_n635), .ZN(new_n959));
  INV_X1    g773(.A(new_n904), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n954), .B1(new_n960), .B2(new_n941), .ZN(new_n961));
  INV_X1    g775(.A(new_n635), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(KEYINPUT120), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n956), .B1(new_n959), .B2(new_n963), .ZN(G63));
  XNOR2_X1  g778(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n436), .A2(new_n283), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n925), .A2(new_n877), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n430), .B(KEYINPUT123), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n935), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT122), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT61), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n925), .A2(new_n665), .A3(new_n877), .A4(new_n967), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n970), .B(new_n973), .C1(new_n971), .C2(KEYINPUT61), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G66));
  NAND2_X1  g791(.A1(new_n845), .A2(new_n898), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n312), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n315), .A2(G224), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n979), .B(KEYINPUT124), .C1(new_n312), .C2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(KEYINPUT124), .B2(new_n979), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n280), .B(new_n281), .C1(G898), .C2(new_n312), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n982), .B(new_n983), .Z(G69));
  INV_X1    g798(.A(new_n786), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n759), .B1(new_n785), .B2(new_n778), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n790), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n748), .A2(new_n647), .ZN(new_n988));
  NOR4_X1   g802(.A1(new_n835), .A2(new_n775), .A3(new_n689), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n869), .A2(new_n714), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n841), .A2(new_n312), .A3(new_n825), .A4(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n682), .B2(new_n312), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n368), .A2(new_n369), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(new_n482), .Z(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(G227), .A2(G900), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(G953), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT62), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n999), .A2(KEYINPUT125), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n990), .B2(new_n710), .ZN(new_n1001));
  INV_X1    g815(.A(new_n691), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n781), .A2(new_n1002), .A3(new_n444), .A4(new_n858), .ZN(new_n1003));
  INV_X1    g817(.A(new_n710), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n687), .A2(new_n714), .A3(new_n756), .ZN(new_n1005));
  AOI22_X1  g819(.A1(new_n1004), .A2(new_n1005), .B1(KEYINPUT125), .B2(new_n999), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1001), .B(new_n1003), .C1(new_n1006), .C2(new_n1000), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n841), .A2(new_n825), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n995), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1009), .A2(new_n312), .A3(new_n1010), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n996), .A2(new_n998), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n998), .B1(new_n996), .B2(new_n1011), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(G72));
  INV_X1    g828(.A(new_n978), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n841), .A2(new_n825), .A3(new_n1015), .A4(new_n991), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n373), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n374), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1023), .A2(KEYINPUT127), .A3(new_n949), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT127), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1021), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n1026), .B2(new_n935), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n902), .A2(new_n903), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1020), .A2(new_n374), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1029), .A2(new_n1018), .A3(new_n1031), .A4(new_n1021), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT126), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n841), .A2(new_n825), .A3(new_n1015), .A4(new_n1008), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n1018), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(new_n1035), .B2(new_n1030), .ZN(new_n1036));
  AOI211_X1 g850(.A(KEYINPUT126), .B(new_n1031), .C1(new_n1034), .C2(new_n1018), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1032), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1028), .A2(new_n1038), .ZN(G57));
endmodule


