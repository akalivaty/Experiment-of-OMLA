

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n1024, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U551 ( .A(n1024), .Z(G160) );
  NOR2_X1 U552 ( .A1(n708), .A2(n707), .ZN(n691) );
  XNOR2_X1 U553 ( .A(n723), .B(n722), .ZN(n725) );
  AND2_X1 U554 ( .A1(n725), .A2(n724), .ZN(n518) );
  XNOR2_X1 U555 ( .A(KEYINPUT101), .B(KEYINPUT30), .ZN(n722) );
  INV_X1 U556 ( .A(G168), .ZN(n724) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n715) );
  XNOR2_X1 U558 ( .A(n716), .B(n715), .ZN(n720) );
  AND2_X1 U559 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U560 ( .A1(G8), .A2(n694), .ZN(n763) );
  INV_X1 U561 ( .A(G651), .ZN(n537) );
  XNOR2_X1 U562 ( .A(KEYINPUT15), .B(n599), .ZN(n966) );
  NOR2_X2 U563 ( .A1(G2104), .A2(n522), .ZN(n878) );
  XOR2_X1 U564 ( .A(KEYINPUT65), .B(n536), .Z(n640) );
  INV_X1 U565 ( .A(KEYINPUT66), .ZN(n529) );
  XNOR2_X1 U566 ( .A(n530), .B(n529), .ZN(n1024) );
  XNOR2_X1 U567 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n520) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XNOR2_X2 U569 ( .A(n520), .B(n519), .ZN(n882) );
  NAND2_X1 U570 ( .A1(n882), .A2(G137), .ZN(n528) );
  INV_X1 U571 ( .A(G2105), .ZN(n522) );
  AND2_X2 U572 ( .A1(n522), .A2(G2104), .ZN(n881) );
  NAND2_X1 U573 ( .A1(G101), .A2(n881), .ZN(n521) );
  XNOR2_X1 U574 ( .A(n521), .B(KEYINPUT23), .ZN(n526) );
  AND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U576 ( .A1(G113), .A2(n877), .ZN(n524) );
  NAND2_X1 U577 ( .A1(G125), .A2(n878), .ZN(n523) );
  NAND2_X1 U578 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n530) );
  NOR2_X1 U581 ( .A1(G543), .A2(G651), .ZN(n636) );
  NAND2_X1 U582 ( .A1(G89), .A2(n636), .ZN(n531) );
  XNOR2_X1 U583 ( .A(n531), .B(KEYINPUT4), .ZN(n532) );
  XNOR2_X1 U584 ( .A(n532), .B(KEYINPUT76), .ZN(n534) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  NOR2_X1 U586 ( .A1(n623), .A2(n537), .ZN(n637) );
  NAND2_X1 U587 ( .A1(G76), .A2(n637), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U589 ( .A(n535), .B(KEYINPUT5), .ZN(n544) );
  NOR2_X1 U590 ( .A1(n623), .A2(G651), .ZN(n536) );
  NAND2_X1 U591 ( .A1(n640), .A2(G51), .ZN(n541) );
  NOR2_X1 U592 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U593 ( .A(KEYINPUT68), .B(n538), .Z(n539) );
  XNOR2_X2 U594 ( .A(KEYINPUT1), .B(n539), .ZN(n641) );
  NAND2_X1 U595 ( .A1(G63), .A2(n641), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U597 ( .A(KEYINPUT6), .B(n542), .Z(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U599 ( .A(n545), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U600 ( .A1(G85), .A2(n636), .ZN(n547) );
  NAND2_X1 U601 ( .A1(G72), .A2(n637), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U603 ( .A1(n640), .A2(G47), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G60), .A2(n641), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U606 ( .A1(n551), .A2(n550), .ZN(G290) );
  NAND2_X1 U607 ( .A1(G99), .A2(n881), .ZN(n553) );
  NAND2_X1 U608 ( .A1(G111), .A2(n877), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U610 ( .A(KEYINPUT82), .B(n554), .Z(n561) );
  XOR2_X1 U611 ( .A(KEYINPUT80), .B(KEYINPUT18), .Z(n556) );
  NAND2_X1 U612 ( .A1(G123), .A2(n878), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n556), .B(n555), .ZN(n559) );
  NAND2_X1 U614 ( .A1(G135), .A2(n882), .ZN(n557) );
  XNOR2_X1 U615 ( .A(KEYINPUT81), .B(n557), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n919) );
  XNOR2_X1 U618 ( .A(G2096), .B(n919), .ZN(n562) );
  OR2_X1 U619 ( .A1(G2100), .A2(n562), .ZN(G156) );
  NAND2_X1 U620 ( .A1(n640), .A2(G53), .ZN(n564) );
  NAND2_X1 U621 ( .A1(G65), .A2(n641), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G91), .A2(n636), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G78), .A2(n637), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n971) );
  INV_X1 U627 ( .A(n971), .ZN(G299) );
  INV_X1 U628 ( .A(G132), .ZN(G219) );
  INV_X1 U629 ( .A(G82), .ZN(G220) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G94), .A2(G452), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT70), .B(n569), .Z(G173) );
  XOR2_X1 U633 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n571) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U636 ( .A(KEYINPUT72), .B(n572), .Z(n824) );
  NAND2_X1 U637 ( .A1(n824), .A2(G567), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  NAND2_X1 U639 ( .A1(n641), .A2(G56), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n574), .Z(n581) );
  NAND2_X1 U641 ( .A1(G81), .A2(n636), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT12), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n576), .B(KEYINPUT74), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G68), .A2(n637), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(n579), .Z(n580) );
  NOR2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n640), .A2(G43), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n965) );
  INV_X1 U650 ( .A(G860), .ZN(n606) );
  OR2_X1 U651 ( .A1(n965), .A2(n606), .ZN(G153) );
  NAND2_X1 U652 ( .A1(n640), .A2(G52), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G64), .A2(n641), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U655 ( .A1(G90), .A2(n636), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G77), .A2(n637), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U658 ( .A(KEYINPUT9), .B(n588), .Z(n589) );
  NOR2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U660 ( .A(KEYINPUT69), .B(n591), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U662 ( .A1(n640), .A2(G54), .ZN(n598) );
  NAND2_X1 U663 ( .A1(G92), .A2(n636), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G79), .A2(n637), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G66), .A2(n641), .ZN(n594) );
  XNOR2_X1 U667 ( .A(KEYINPUT75), .B(n594), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  INV_X1 U670 ( .A(n966), .ZN(n708) );
  INV_X1 U671 ( .A(G868), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n708), .A2(n602), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(G284) );
  NOR2_X1 U674 ( .A1(G286), .A2(n602), .ZN(n604) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U677 ( .A(KEYINPUT77), .B(n605), .Z(G297) );
  NAND2_X1 U678 ( .A1(n606), .A2(G559), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n607), .A2(n966), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT16), .ZN(n610) );
  XOR2_X1 U681 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n609) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n965), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n966), .A2(G868), .ZN(n611) );
  NOR2_X1 U685 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U687 ( .A1(n966), .A2(G559), .ZN(n653) );
  XNOR2_X1 U688 ( .A(n965), .B(n653), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n614), .A2(G860), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n640), .A2(G55), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G67), .A2(n641), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G93), .A2(n636), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G80), .A2(n637), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U696 ( .A(KEYINPUT83), .B(n619), .Z(n620) );
  NOR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n656) );
  XNOR2_X1 U698 ( .A(n622), .B(n656), .ZN(G145) );
  NAND2_X1 U699 ( .A1(G49), .A2(n640), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G87), .A2(n623), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U702 ( .A1(n641), .A2(n626), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G651), .A2(G74), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(G288) );
  NAND2_X1 U705 ( .A1(n636), .A2(G86), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G61), .A2(n641), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n637), .A2(G73), .ZN(n631) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n631), .Z(n632) );
  NOR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n640), .A2(G48), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G88), .A2(n636), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G75), .A2(n637), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n640), .A2(G50), .ZN(n643) );
  NAND2_X1 U717 ( .A1(G62), .A2(n641), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n645), .A2(n644), .ZN(G166) );
  INV_X1 U720 ( .A(G166), .ZN(G303) );
  XOR2_X1 U721 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n646) );
  XNOR2_X1 U722 ( .A(G288), .B(n646), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n647), .B(G290), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n648), .B(G305), .ZN(n652) );
  XOR2_X1 U725 ( .A(G303), .B(n656), .Z(n650) );
  XOR2_X1 U726 ( .A(n965), .B(G299), .Z(n649) );
  XNOR2_X1 U727 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(n893) );
  XNOR2_X1 U729 ( .A(KEYINPUT85), .B(n653), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n893), .B(n654), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n655), .A2(G868), .ZN(n658) );
  OR2_X1 U732 ( .A1(G868), .A2(n656), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U734 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XOR2_X1 U735 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n659) );
  XNOR2_X1 U736 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U737 ( .A1(n661), .A2(G2090), .ZN(n664) );
  XOR2_X1 U738 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n662) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  XNOR2_X1 U740 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U744 ( .A1(G69), .A2(G120), .ZN(n666) );
  NOR2_X1 U745 ( .A1(G237), .A2(n666), .ZN(n667) );
  XNOR2_X1 U746 ( .A(KEYINPUT90), .B(n667), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n668), .A2(G108), .ZN(n829) );
  NAND2_X1 U748 ( .A1(G567), .A2(n829), .ZN(n674) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n669) );
  XNOR2_X1 U750 ( .A(KEYINPUT22), .B(n669), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n670), .A2(G96), .ZN(n671) );
  NOR2_X1 U752 ( .A1(n671), .A2(G218), .ZN(n672) );
  XNOR2_X1 U753 ( .A(n672), .B(KEYINPUT89), .ZN(n830) );
  NAND2_X1 U754 ( .A1(G2106), .A2(n830), .ZN(n673) );
  NAND2_X1 U755 ( .A1(n674), .A2(n673), .ZN(n831) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U757 ( .A1(n831), .A2(n675), .ZN(n827) );
  NAND2_X1 U758 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U759 ( .A1(G102), .A2(n881), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G138), .A2(n882), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n681) );
  NAND2_X1 U762 ( .A1(G114), .A2(n877), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G126), .A2(n878), .ZN(n678) );
  NAND2_X1 U764 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n681), .A2(n680), .ZN(G164) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n770) );
  INV_X1 U767 ( .A(n770), .ZN(n682) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n769) );
  NOR2_X2 U769 ( .A1(n682), .A2(n769), .ZN(n695) );
  INV_X1 U770 ( .A(n695), .ZN(n694) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n683) );
  XOR2_X1 U772 ( .A(n683), .B(KEYINPUT98), .Z(n684) );
  XNOR2_X1 U773 ( .A(KEYINPUT24), .B(n684), .ZN(n685) );
  NOR2_X1 U774 ( .A1(n763), .A2(n685), .ZN(n768) );
  NAND2_X1 U775 ( .A1(n695), .A2(G1996), .ZN(n686) );
  XNOR2_X1 U776 ( .A(n686), .B(KEYINPUT26), .ZN(n687) );
  XNOR2_X1 U777 ( .A(n687), .B(KEYINPUT64), .ZN(n690) );
  AND2_X1 U778 ( .A1(G1341), .A2(n694), .ZN(n688) );
  NOR2_X1 U779 ( .A1(n688), .A2(n965), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n707) );
  XOR2_X1 U781 ( .A(KEYINPUT100), .B(n691), .Z(n702) );
  NOR2_X1 U782 ( .A1(n695), .A2(G1348), .ZN(n693) );
  NOR2_X1 U783 ( .A1(G2067), .A2(n694), .ZN(n692) );
  NOR2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n700) );
  NAND2_X1 U785 ( .A1(n694), .A2(G1956), .ZN(n698) );
  NAND2_X1 U786 ( .A1(n695), .A2(G2072), .ZN(n696) );
  XOR2_X1 U787 ( .A(n696), .B(KEYINPUT27), .Z(n697) );
  NAND2_X1 U788 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n699), .B(KEYINPUT99), .ZN(n703) );
  NAND2_X1 U790 ( .A1(n971), .A2(n703), .ZN(n706) );
  AND2_X1 U791 ( .A1(n700), .A2(n706), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n714) );
  NOR2_X1 U793 ( .A1(n971), .A2(n703), .ZN(n705) );
  INV_X1 U794 ( .A(KEYINPUT28), .ZN(n704) );
  XNOR2_X1 U795 ( .A(n705), .B(n704), .ZN(n712) );
  INV_X1 U796 ( .A(n706), .ZN(n710) );
  NAND2_X1 U797 ( .A1(n708), .A2(n707), .ZN(n709) );
  OR2_X1 U798 ( .A1(n710), .A2(n709), .ZN(n711) );
  AND2_X1 U799 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U800 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U801 ( .A1(G1961), .A2(n694), .ZN(n718) );
  XOR2_X1 U802 ( .A(KEYINPUT25), .B(G2078), .Z(n946) );
  NAND2_X1 U803 ( .A1(n695), .A2(n946), .ZN(n717) );
  NAND2_X1 U804 ( .A1(n718), .A2(n717), .ZN(n726) );
  OR2_X1 U805 ( .A1(G301), .A2(n726), .ZN(n719) );
  NAND2_X1 U806 ( .A1(n720), .A2(n719), .ZN(n732) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n763), .ZN(n743) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n694), .ZN(n742) );
  NOR2_X1 U809 ( .A1(n743), .A2(n742), .ZN(n721) );
  NAND2_X1 U810 ( .A1(G8), .A2(n721), .ZN(n723) );
  NAND2_X1 U811 ( .A1(G301), .A2(n726), .ZN(n727) );
  XOR2_X1 U812 ( .A(KEYINPUT102), .B(n727), .Z(n728) );
  NOR2_X1 U813 ( .A1(n518), .A2(n728), .ZN(n730) );
  INV_X1 U814 ( .A(KEYINPUT31), .ZN(n729) );
  XNOR2_X1 U815 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U816 ( .A1(n732), .A2(n731), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n744), .A2(G286), .ZN(n740) );
  INV_X1 U818 ( .A(G8), .ZN(n738) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n763), .ZN(n734) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n694), .ZN(n733) );
  NOR2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U822 ( .A(KEYINPUT103), .B(n735), .Z(n736) );
  NAND2_X1 U823 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U825 ( .A(n741), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U826 ( .A1(G8), .A2(n742), .ZN(n747) );
  INV_X1 U827 ( .A(n744), .ZN(n745) );
  NOR2_X1 U828 ( .A1(n743), .A2(n745), .ZN(n746) );
  NAND2_X1 U829 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U830 ( .A1(n749), .A2(n748), .ZN(n762) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n755) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U833 ( .A1(n755), .A2(n750), .ZN(n975) );
  NAND2_X1 U834 ( .A1(n762), .A2(n975), .ZN(n751) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n970) );
  NAND2_X1 U836 ( .A1(n751), .A2(n970), .ZN(n752) );
  XNOR2_X1 U837 ( .A(n752), .B(KEYINPUT104), .ZN(n753) );
  NOR2_X1 U838 ( .A1(n753), .A2(n763), .ZN(n754) );
  NOR2_X1 U839 ( .A1(KEYINPUT33), .A2(n754), .ZN(n758) );
  NAND2_X1 U840 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n756), .A2(n763), .ZN(n757) );
  NOR2_X1 U842 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U843 ( .A(G1981), .B(G305), .Z(n981) );
  NAND2_X1 U844 ( .A1(n759), .A2(n981), .ZN(n766) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U846 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U847 ( .A1(n762), .A2(n761), .ZN(n764) );
  NAND2_X1 U848 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U849 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U850 ( .A1(n768), .A2(n767), .ZN(n804) );
  NOR2_X1 U851 ( .A1(n770), .A2(n769), .ZN(n817) );
  XOR2_X1 U852 ( .A(G2067), .B(KEYINPUT37), .Z(n771) );
  XNOR2_X1 U853 ( .A(KEYINPUT91), .B(n771), .ZN(n815) );
  XNOR2_X1 U854 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n776) );
  NAND2_X1 U855 ( .A1(G116), .A2(n877), .ZN(n773) );
  NAND2_X1 U856 ( .A1(G128), .A2(n878), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U858 ( .A(n774), .B(KEYINPUT35), .ZN(n775) );
  XNOR2_X1 U859 ( .A(n776), .B(n775), .ZN(n782) );
  NAND2_X1 U860 ( .A1(n881), .A2(G104), .ZN(n777) );
  XNOR2_X1 U861 ( .A(n777), .B(KEYINPUT92), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G140), .A2(n882), .ZN(n778) );
  NAND2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U864 ( .A(KEYINPUT34), .B(n780), .ZN(n781) );
  NOR2_X1 U865 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U866 ( .A(KEYINPUT36), .B(n783), .ZN(n874) );
  NOR2_X1 U867 ( .A1(n815), .A2(n874), .ZN(n933) );
  NAND2_X1 U868 ( .A1(n817), .A2(n933), .ZN(n813) );
  XOR2_X1 U869 ( .A(KEYINPUT38), .B(KEYINPUT96), .Z(n785) );
  NAND2_X1 U870 ( .A1(G105), .A2(n881), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n785), .B(n784), .ZN(n790) );
  NAND2_X1 U872 ( .A1(G117), .A2(n877), .ZN(n787) );
  NAND2_X1 U873 ( .A1(G129), .A2(n878), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U875 ( .A(KEYINPUT95), .B(n788), .Z(n789) );
  NOR2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n882), .A2(G141), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n869) );
  AND2_X1 U879 ( .A1(n869), .A2(G1996), .ZN(n800) );
  NAND2_X1 U880 ( .A1(G95), .A2(n881), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G131), .A2(n882), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G107), .A2(n877), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G119), .A2(n878), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n868) );
  INV_X1 U887 ( .A(G1991), .ZN(n843) );
  NOR2_X1 U888 ( .A1(n868), .A2(n843), .ZN(n799) );
  NOR2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n924) );
  XNOR2_X1 U890 ( .A(KEYINPUT97), .B(n817), .ZN(n801) );
  NOR2_X1 U891 ( .A1(n924), .A2(n801), .ZN(n809) );
  INV_X1 U892 ( .A(n809), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n813), .A2(n802), .ZN(n803) );
  NOR2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n806) );
  XNOR2_X1 U895 ( .A(G1986), .B(G290), .ZN(n977) );
  NAND2_X1 U896 ( .A1(n977), .A2(n817), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n820) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n869), .ZN(n926) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n807) );
  AND2_X1 U900 ( .A1(n843), .A2(n868), .ZN(n922) );
  NOR2_X1 U901 ( .A1(n807), .A2(n922), .ZN(n808) );
  NOR2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U903 ( .A(KEYINPUT105), .B(n810), .Z(n811) );
  NOR2_X1 U904 ( .A1(n926), .A2(n811), .ZN(n812) );
  XNOR2_X1 U905 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U907 ( .A1(n815), .A2(n874), .ZN(n930) );
  NAND2_X1 U908 ( .A1(n816), .A2(n930), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n823) );
  XOR2_X1 U911 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n821) );
  XNOR2_X1 U912 ( .A(KEYINPUT40), .B(n821), .ZN(n822) );
  XNOR2_X1 U913 ( .A(n823), .B(n822), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n824), .ZN(G217) );
  INV_X1 U915 ( .A(n824), .ZN(G223) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U917 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n826) );
  XNOR2_X1 U919 ( .A(KEYINPUT110), .B(n826), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G108), .ZN(G238) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U928 ( .A(KEYINPUT111), .B(n831), .ZN(G319) );
  XOR2_X1 U929 ( .A(G2100), .B(G2096), .Z(n833) );
  XNOR2_X1 U930 ( .A(KEYINPUT42), .B(G2678), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U932 ( .A(KEYINPUT43), .B(G2090), .Z(n835) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U935 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(G227) );
  XOR2_X1 U938 ( .A(KEYINPUT113), .B(G1981), .Z(n841) );
  XNOR2_X1 U939 ( .A(G1966), .B(G1961), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U941 ( .A(n842), .B(KEYINPUT41), .Z(n845) );
  XOR2_X1 U942 ( .A(G1996), .B(n843), .Z(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U944 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1956), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U947 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U948 ( .A(KEYINPUT112), .B(G2474), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n878), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n852), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U952 ( .A1(G112), .A2(n877), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n853), .B(KEYINPUT114), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G100), .A2(n881), .ZN(n857) );
  NAND2_X1 U956 ( .A1(G136), .A2(n882), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U958 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U959 ( .A(G164), .B(KEYINPUT46), .Z(n860) );
  XNOR2_X1 U960 ( .A(n919), .B(n860), .ZN(n873) );
  NAND2_X1 U961 ( .A1(G103), .A2(n881), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G139), .A2(n882), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G115), .A2(n877), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G127), .A2(n878), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n865), .Z(n866) );
  NOR2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n914) );
  XOR2_X1 U969 ( .A(G162), .B(n914), .Z(n871) );
  XOR2_X1 U970 ( .A(n869), .B(n868), .Z(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n876) );
  XNOR2_X1 U973 ( .A(n874), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n891) );
  NAND2_X1 U975 ( .A1(G118), .A2(n877), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G130), .A2(n878), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U978 ( .A1(G106), .A2(n881), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G142), .A2(n882), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U981 ( .A(KEYINPUT115), .B(n885), .ZN(n886) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n886), .ZN(n887) );
  NOR2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U984 ( .A(G160), .B(n889), .Z(n890) );
  XNOR2_X1 U985 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U986 ( .A1(G37), .A2(n892), .ZN(G395) );
  INV_X1 U987 ( .A(G301), .ZN(G171) );
  XOR2_X1 U988 ( .A(G286), .B(n966), .Z(n894) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U990 ( .A(n895), .B(G171), .Z(n896) );
  NOR2_X1 U991 ( .A1(G37), .A2(n896), .ZN(G397) );
  XNOR2_X1 U992 ( .A(G2451), .B(G2446), .ZN(n906) );
  XOR2_X1 U993 ( .A(G2430), .B(KEYINPUT109), .Z(n898) );
  XNOR2_X1 U994 ( .A(G2454), .B(G2435), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U996 ( .A(G2438), .B(KEYINPUT108), .Z(n900) );
  XNOR2_X1 U997 ( .A(G1348), .B(G1341), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U999 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U1000 ( .A(G2443), .B(G2427), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(n907), .A2(G14), .ZN(n913) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(n913), .ZN(G401) );
  XOR2_X1 U1012 ( .A(G2072), .B(n914), .Z(n916) );
  XOR2_X1 U1013 ( .A(G164), .B(G2078), .Z(n915) );
  NOR2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1015 ( .A(KEYINPUT50), .B(n917), .Z(n936) );
  XNOR2_X1 U1016 ( .A(G2084), .B(KEYINPUT116), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n918), .B(G160), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n929) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n927), .B(KEYINPUT51), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n931) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(KEYINPUT117), .B(n934), .ZN(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(n937), .ZN(n939) );
  INV_X1 U1030 ( .A(KEYINPUT55), .ZN(n938) );
  NAND2_X1 U1031 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1032 ( .A1(n940), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1033 ( .A(G2084), .B(KEYINPUT54), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(G34), .ZN(n956) );
  XOR2_X1 U1035 ( .A(G25), .B(G1991), .Z(n942) );
  NAND2_X1 U1036 ( .A1(n942), .A2(G28), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(G32), .B(G1996), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(KEYINPUT120), .B(n943), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n953) );
  XNOR2_X1 U1040 ( .A(n946), .B(G27), .ZN(n951) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G2072), .B(G33), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(KEYINPUT119), .B(n949), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1047 ( .A(KEYINPUT53), .B(n954), .Z(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1049 ( .A(G2090), .B(KEYINPUT118), .Z(n957) );
  XNOR2_X1 U1050 ( .A(G35), .B(n957), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1052 ( .A(KEYINPUT55), .B(n960), .Z(n962) );
  INV_X1 U1053 ( .A(G29), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(G11), .A2(n963), .ZN(n1020) );
  INV_X1 U1056 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1057 ( .A(n1016), .B(KEYINPUT56), .Z(n990) );
  XOR2_X1 U1058 ( .A(G1961), .B(G301), .Z(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT122), .ZN(n988) );
  XNOR2_X1 U1060 ( .A(G1341), .B(n965), .ZN(n968) );
  XOR2_X1 U1061 ( .A(G1348), .B(n966), .Z(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n980) );
  NAND2_X1 U1063 ( .A1(G1971), .A2(G303), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1065 ( .A(G1956), .B(n971), .Z(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(KEYINPUT123), .B(n978), .Z(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n986) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G168), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(n983), .B(KEYINPUT57), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(n984), .B(KEYINPUT121), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n1018) );
  XOR2_X1 U1078 ( .A(G1348), .B(KEYINPUT59), .Z(n991) );
  XNOR2_X1 U1079 ( .A(G4), .B(n991), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(G20), .B(G1956), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1086 ( .A(KEYINPUT60), .B(n998), .Z(n999) );
  XNOR2_X1 U1087 ( .A(KEYINPUT124), .B(n999), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G21), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G5), .B(G1961), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1013) );
  XNOR2_X1 U1092 ( .A(G1986), .B(KEYINPUT126), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(n1004), .B(G24), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT125), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(KEYINPUT127), .B(n1010), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .ZN(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

