//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT74), .B1(new_n187), .B2(G125), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT74), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT19), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n190), .A2(G140), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT91), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n198), .A2(new_n199), .A3(new_n200), .A4(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n193), .A3(new_n197), .A4(new_n200), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT91), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n195), .A2(new_n196), .A3(new_n202), .A4(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT92), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n187), .A3(G125), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT76), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n190), .A2(G140), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(new_n188), .B2(new_n191), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n212), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT75), .B1(new_n212), .B2(KEYINPUT16), .ZN(new_n214));
  OAI211_X1 g028(.A(G146), .B(new_n210), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(G237), .A2(G953), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(G143), .A3(G214), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(G143), .B1(new_n216), .B2(G214), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n219), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n194), .A2(KEYINPUT19), .B1(KEYINPUT91), .B2(new_n203), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT92), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n196), .A4(new_n202), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n206), .A2(new_n215), .A3(new_n224), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n217), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT18), .A2(G131), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n198), .A2(new_n196), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n212), .B2(new_n196), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G113), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT93), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT17), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n220), .A2(new_n223), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT94), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n196), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n229), .A2(KEYINPUT17), .A3(G131), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n245), .A2(new_n247), .A3(new_n215), .A4(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n238), .A3(new_n234), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n235), .A2(new_n251), .A3(new_n239), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n241), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(G475), .A2(G902), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT20), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n241), .A2(new_n250), .A3(new_n252), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(new_n254), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(G234), .A2(G237), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(G952), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT21), .B(G898), .Z(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(G902), .A3(G953), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G128), .B(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT13), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G128), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n268), .B(G134), .C1(KEYINPUT13), .C2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G116), .B(G122), .ZN(new_n272));
  INV_X1    g086(.A(G107), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n267), .B(new_n275), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n273), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT14), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G116), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT14), .A3(G122), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(G107), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(new_n279), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g100(.A(KEYINPUT9), .B(G234), .Z(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(G217), .A3(new_n262), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n288), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n277), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  INV_X1    g107(.A(G478), .ZN(new_n294));
  NOR2_X1   g108(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n292), .A2(new_n293), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n292), .B2(new_n293), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n303), .A2(KEYINPUT96), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(KEYINPUT96), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n249), .A2(new_n234), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n239), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n250), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n293), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G475), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n260), .A2(new_n266), .A3(new_n306), .A4(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(G110), .B(G140), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n262), .A2(G227), .ZN(new_n314));
  XOR2_X1   g128(.A(new_n313), .B(new_n314), .Z(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT79), .Z(new_n316));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT4), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n273), .A2(G104), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n237), .B2(G107), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n273), .A2(KEYINPUT3), .A3(G104), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G101), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n318), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n319), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n273), .A2(KEYINPUT3), .A3(G104), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT3), .B1(new_n273), .B2(G104), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G101), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n269), .A2(G146), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n196), .A2(G143), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT0), .ZN(new_n334));
  INV_X1    g148(.A(G128), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n332), .B(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n334), .A2(new_n335), .ZN(new_n337));
  NOR2_X1   g151(.A1(KEYINPUT0), .A2(G128), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G143), .B(G146), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n329), .A2(new_n318), .A3(G101), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n331), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT11), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n275), .B2(G137), .ZN(new_n345));
  INV_X1    g159(.A(G137), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT11), .A3(G134), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n275), .A2(G137), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G131), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n345), .A2(new_n347), .A3(new_n222), .A4(new_n348), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT80), .B1(new_n273), .B2(G104), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n237), .A3(G107), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n273), .A2(G104), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G101), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n335), .A2(KEYINPUT1), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n332), .A3(new_n333), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n335), .A2(new_n196), .A3(G143), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n269), .B(G146), .C1(new_n335), .C2(KEYINPUT1), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n326), .B(new_n324), .C1(new_n327), .C2(new_n328), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n359), .A2(new_n364), .A3(new_n365), .A4(KEYINPUT10), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n343), .A2(new_n353), .A3(new_n366), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n359), .A2(new_n365), .ZN(new_n371));
  INV_X1    g185(.A(new_n364), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n367), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT12), .B1(new_n374), .B2(new_n352), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n364), .B1(new_n365), .B2(new_n359), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT12), .B(new_n352), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n317), .B(new_n370), .C1(new_n375), .C2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n352), .B1(new_n376), .B2(new_n377), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT12), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n378), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n317), .B1(new_n385), .B2(new_n370), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n316), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n370), .A2(new_n315), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n343), .A2(new_n366), .A3(new_n369), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n352), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(G902), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G469), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n375), .A2(new_n379), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(new_n388), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n315), .B1(new_n391), .B2(new_n370), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n394), .B(new_n293), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n315), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n369), .A2(new_n366), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n353), .B1(new_n402), .B2(new_n343), .ZN(new_n403));
  INV_X1    g217(.A(new_n370), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n385), .A2(new_n370), .A3(new_n315), .ZN(new_n406));
  AOI21_X1  g220(.A(G902), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT82), .B1(new_n407), .B2(new_n394), .ZN(new_n408));
  OAI22_X1  g222(.A1(new_n393), .A2(new_n394), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G221), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n287), .B2(new_n293), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G214), .B1(G237), .B2(G902), .ZN(new_n414));
  OAI21_X1  g228(.A(G210), .B1(G237), .B2(G902), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT67), .ZN(new_n417));
  INV_X1    g231(.A(G119), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(G116), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n282), .A2(KEYINPUT67), .A3(G119), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n282), .A2(G119), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(KEYINPUT2), .A2(G113), .ZN(new_n424));
  NOR2_X1   g238(.A1(KEYINPUT2), .A2(G113), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT68), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n422), .B1(new_n419), .B2(new_n420), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT68), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n426), .ZN(new_n431));
  INV_X1    g245(.A(G113), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n422), .ZN(new_n434));
  INV_X1    g248(.A(new_n433), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n428), .A2(new_n431), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n371), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT87), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n428), .A2(new_n431), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n429), .A2(KEYINPUT5), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n434), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n436), .A2(new_n434), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n429), .A2(new_n430), .A3(new_n426), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n430), .B1(new_n429), .B2(new_n426), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n371), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n439), .A2(new_n443), .A3(new_n449), .ZN(new_n450));
  XOR2_X1   g264(.A(G110), .B(G122), .Z(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT8), .Z(new_n452));
  AND2_X1   g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n341), .B2(new_n190), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n332), .A2(new_n333), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n337), .B2(new_n338), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n457), .A2(KEYINPUT85), .A3(G125), .A4(new_n336), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(KEYINPUT86), .A3(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n372), .A2(new_n190), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n262), .A2(G224), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(new_n464), .B2(KEYINPUT89), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(KEYINPUT89), .B2(new_n464), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n455), .A2(new_n463), .A3(new_n458), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(KEYINPUT7), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT88), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n440), .A2(new_n438), .A3(new_n444), .ZN(new_n472));
  INV_X1    g286(.A(new_n451), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n429), .A2(new_n426), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n428), .B2(new_n431), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n331), .A2(new_n342), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n472), .B(new_n473), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n468), .A2(new_n478), .A3(new_n469), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n467), .A2(new_n471), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n293), .B1(new_n453), .B2(new_n480), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n476), .A2(new_n475), .B1(new_n447), .B2(new_n371), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT84), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT84), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n472), .B(new_n484), .C1(new_n475), .C2(new_n476), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n451), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n483), .A2(KEYINPUT6), .A3(new_n451), .A4(new_n485), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n477), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n464), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n416), .B(new_n481), .C1(new_n490), .C2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n486), .A2(new_n487), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n477), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n481), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n415), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n414), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n312), .A2(new_n413), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G472), .A2(G902), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT73), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n352), .A2(new_n341), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n475), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n346), .A2(KEYINPUT66), .A3(G134), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n508), .B1(new_n346), .B2(G134), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n275), .A2(G137), .ZN(new_n510));
  OAI211_X1 g324(.A(G131), .B(new_n507), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n364), .A2(new_n351), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n504), .B1(new_n506), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT65), .B1(new_n352), .B2(new_n341), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n352), .A2(KEYINPUT65), .A3(new_n341), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n512), .A3(new_n517), .ZN(new_n518));
  OAI22_X1  g332(.A1(new_n445), .A2(new_n446), .B1(new_n429), .B2(new_n426), .ZN(new_n519));
  INV_X1    g333(.A(new_n506), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n512), .B(KEYINPUT69), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n514), .B1(new_n522), .B2(new_n504), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n216), .A2(G210), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT71), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n216), .A2(new_n526), .A3(G210), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT26), .B(G101), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n528), .B1(new_n525), .B2(new_n527), .ZN(new_n533));
  OR3_X1    g347(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n532), .B1(new_n530), .B2(new_n533), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT69), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n511), .A2(new_n351), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(new_n364), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n538), .A2(new_n364), .A3(new_n351), .A4(new_n511), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT30), .B(new_n505), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n352), .A2(KEYINPUT65), .A3(new_n341), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n543), .A2(new_n515), .A3(new_n513), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n519), .B(new_n542), .C1(new_n544), .C2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n475), .B(new_n505), .C1(new_n540), .C2(new_n541), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n548), .A2(new_n549), .A3(new_n536), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n548), .B2(new_n536), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT31), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n547), .B(KEYINPUT31), .C1(new_n550), .C2(new_n551), .ZN(new_n555));
  AOI221_X4 g369(.A(new_n503), .B1(new_n523), .B2(new_n537), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n523), .A2(new_n537), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT73), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n502), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT32), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n548), .A2(new_n536), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT72), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n548), .A2(new_n536), .A3(new_n549), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT31), .B1(new_n566), .B2(new_n547), .ZN(new_n567));
  INV_X1    g381(.A(new_n555), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n558), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n503), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n557), .A2(KEYINPUT73), .A3(new_n558), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n502), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n547), .A2(new_n548), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n537), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT29), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n575), .B(new_n576), .C1(new_n523), .C2(new_n537), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n521), .A2(new_n505), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n548), .B1(new_n579), .B2(new_n475), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT28), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n514), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n536), .A2(KEYINPUT29), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n577), .B(new_n293), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G472), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n562), .A2(new_n573), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT23), .B1(new_n335), .B2(G119), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n418), .A2(G128), .ZN(new_n592));
  MUX2_X1   g406(.A(new_n591), .B(KEYINPUT23), .S(new_n592), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G110), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT24), .B(G110), .Z(new_n595));
  XNOR2_X1  g409(.A(G119), .B(G128), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n247), .B2(new_n215), .ZN(new_n599));
  OAI22_X1  g413(.A1(new_n593), .A2(G110), .B1(new_n596), .B2(new_n595), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n215), .A2(new_n232), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT77), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n598), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n192), .A2(KEYINPUT16), .A3(new_n193), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT75), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n212), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G146), .B1(new_n609), .B2(new_n210), .ZN(new_n610));
  AOI211_X1 g424(.A(new_n196), .B(new_n209), .C1(new_n607), .C2(new_n608), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n604), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n215), .A2(new_n232), .A3(new_n600), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT77), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n590), .B1(new_n603), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n599), .A2(new_n601), .A3(new_n590), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n293), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT25), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n602), .B1(new_n599), .B2(new_n601), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n612), .A2(KEYINPUT77), .A3(new_n613), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n616), .B1(new_n622), .B2(new_n590), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT25), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n293), .ZN(new_n625));
  INV_X1    g439(.A(G217), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(G234), .B2(new_n293), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n619), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  OR3_X1    g442(.A1(new_n618), .A2(KEYINPUT78), .A3(new_n627), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT78), .B1(new_n618), .B2(new_n627), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n501), .A2(new_n586), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  AOI21_X1  g447(.A(G902), .B1(new_n570), .B2(new_n571), .ZN(new_n634));
  INV_X1    g448(.A(G472), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n560), .B(new_n409), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n628), .A2(new_n629), .A3(new_n630), .A4(new_n412), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT97), .Z(new_n640));
  OAI211_X1 g454(.A(new_n414), .B(new_n266), .C1(new_n494), .C2(new_n499), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n257), .A2(new_n258), .A3(new_n254), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n258), .B1(new_n257), .B2(new_n254), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n311), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT33), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n291), .B(KEYINPUT99), .Z(new_n646));
  NAND2_X1  g460(.A1(new_n288), .A2(KEYINPUT98), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n288), .A2(KEYINPUT98), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n286), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n645), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n292), .A2(KEYINPUT33), .ZN(new_n651));
  OAI211_X1 g465(.A(G478), .B(new_n293), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n292), .A2(new_n293), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n294), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n644), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n641), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n640), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT34), .B(G104), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(G475), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n309), .B2(new_n293), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n256), .B2(new_n259), .ZN(new_n664));
  INV_X1    g478(.A(new_n306), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n640), .A2(new_n641), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT35), .B(G107), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NOR2_X1   g483(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n620), .A2(new_n621), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n671), .B1(new_n620), .B2(new_n621), .ZN(new_n674));
  OAI221_X1 g488(.A(new_n293), .B1(new_n626), .B2(G234), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n628), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n560), .B(new_n676), .C1(new_n634), .C2(new_n635), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n293), .B1(new_n556), .B2(new_n559), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G472), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(KEYINPUT100), .A3(new_n560), .A4(new_n676), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n679), .A2(new_n501), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  XOR2_X1   g499(.A(new_n263), .B(KEYINPUT101), .Z(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  INV_X1    g501(.A(new_n265), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n664), .A2(new_n665), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n500), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n673), .A2(new_n674), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(G902), .A3(new_n627), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n624), .B1(new_n623), .B2(new_n293), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n589), .B1(new_n620), .B2(new_n621), .ZN(new_n696));
  NOR4_X1   g510(.A1(new_n696), .A2(KEYINPUT25), .A3(G902), .A4(new_n616), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n694), .B1(new_n698), .B2(new_n627), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n413), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n586), .A2(new_n692), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT102), .B(G128), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G30));
  XNOR2_X1  g517(.A(new_n689), .B(KEYINPUT39), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n413), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT104), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n644), .A2(new_n414), .A3(new_n665), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n580), .A2(new_n537), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n552), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n711), .A2(KEYINPUT103), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n293), .B1(new_n711), .B2(KEYINPUT103), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n562), .A2(new_n573), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n707), .A2(new_n709), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n494), .A2(new_n499), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT38), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n699), .B1(new_n706), .B2(KEYINPUT40), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n269), .ZN(G45));
  NAND3_X1  g535(.A1(new_n644), .A2(new_n655), .A3(new_n690), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n500), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n586), .A2(new_n700), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  AND2_X1   g539(.A1(new_n586), .A2(new_n631), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n398), .A2(new_n399), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n407), .A2(KEYINPUT82), .A3(new_n394), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n407), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n412), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n727), .A2(new_n728), .B1(G469), .B2(new_n730), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n412), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n726), .A2(new_n657), .A3(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT41), .B(G113), .Z(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT106), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n739), .B(new_n741), .ZN(G15));
  INV_X1    g556(.A(new_n266), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n644), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n586), .A2(new_n631), .A3(new_n744), .A4(new_n665), .ZN(new_n745));
  INV_X1    g559(.A(new_n414), .ZN(new_n746));
  INV_X1    g560(.A(new_n496), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n492), .B1(new_n747), .B2(new_n488), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n416), .B1(new_n748), .B2(new_n481), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n497), .A2(new_n415), .A3(new_n498), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n751), .A2(new_n733), .A3(new_n736), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n745), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n282), .ZN(G18));
  INV_X1    g569(.A(new_n312), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n752), .A2(new_n586), .A3(new_n756), .A4(new_n676), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G119), .ZN(G21));
  NOR3_X1   g572(.A1(new_n708), .A2(new_n717), .A3(new_n743), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n582), .A2(new_n537), .ZN(new_n760));
  AOI211_X1 g574(.A(G472), .B(G902), .C1(new_n760), .C2(new_n557), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n680), .B2(G472), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n759), .A2(new_n631), .A3(new_n738), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G122), .ZN(G24));
  INV_X1    g578(.A(new_n722), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n752), .A2(new_n676), .A3(new_n765), .A4(new_n762), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  NAND3_X1  g581(.A1(new_n749), .A2(new_n750), .A3(new_n414), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n413), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n586), .A2(new_n631), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n774));
  INV_X1    g588(.A(new_n691), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n726), .A2(new_n774), .A3(new_n775), .A4(new_n769), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n586), .A2(new_n631), .A3(new_n775), .A4(new_n769), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT107), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  AOI22_X1  g594(.A1(new_n680), .A2(G472), .B1(new_n572), .B2(new_n502), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n655), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT43), .B1(new_n644), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n260), .A2(new_n785), .A3(new_n311), .A4(new_n655), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n782), .A2(new_n676), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT44), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n494), .A2(new_n499), .A3(new_n746), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n387), .A2(new_n392), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n387), .A2(KEYINPUT45), .A3(new_n392), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(G469), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(G469), .A2(G902), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n795), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n729), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n704), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n412), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n788), .A2(new_n789), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  XOR2_X1   g619(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n799), .A2(new_n729), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT46), .B1(new_n794), .B2(new_n795), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n412), .B(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n800), .B2(new_n412), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n811), .A2(new_n813), .A3(new_n722), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n586), .A2(new_n631), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n789), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  NOR2_X1   g631(.A1(G952), .A2(G953), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n657), .A2(new_n781), .A3(new_n409), .A4(new_n638), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n632), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n819), .B1(new_n632), .B2(new_n820), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n641), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n644), .A2(new_n303), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n637), .A2(new_n824), .A3(new_n638), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n683), .A2(new_n826), .A3(new_n763), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n754), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n823), .A2(new_n828), .A3(new_n739), .A4(new_n757), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n762), .A2(new_n676), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n765), .A3(new_n769), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n586), .A2(new_n664), .A3(new_n700), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n303), .A3(new_n690), .A4(new_n789), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n772), .A2(new_n779), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n586), .B(new_n700), .C1(new_n692), .C2(new_n723), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT111), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n409), .A2(new_n628), .A3(new_n412), .A4(new_n675), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n837), .B1(new_n838), .B2(new_n689), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n708), .A2(new_n717), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT81), .B1(new_n395), .B2(new_n404), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n380), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n842), .A2(new_n316), .B1(new_n391), .B2(new_n389), .ZN(new_n843));
  OAI21_X1  g657(.A(G469), .B1(new_n843), .B2(G902), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n411), .B1(new_n844), .B2(new_n729), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n699), .A2(new_n845), .A3(KEYINPUT111), .A4(new_n690), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n715), .A2(new_n839), .A3(new_n840), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n836), .A2(new_n847), .A3(new_n766), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n836), .A2(new_n847), .A3(new_n766), .A4(KEYINPUT52), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n850), .A2(KEYINPUT113), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT113), .B1(new_n850), .B2(new_n851), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n835), .B2(new_n854), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n772), .A2(new_n779), .A3(new_n831), .A4(new_n833), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n683), .A2(new_n826), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n745), .A2(new_n753), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n757), .A4(new_n763), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n632), .A2(new_n820), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT110), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n632), .A2(new_n819), .A3(new_n820), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n739), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n836), .A2(new_n766), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(KEYINPUT112), .A3(KEYINPUT52), .A4(new_n847), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n851), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n868), .A3(new_n850), .ZN(new_n869));
  AND4_X1   g683(.A1(KEYINPUT53), .A2(new_n856), .A3(new_n864), .A4(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n855), .A2(new_n870), .A3(KEYINPUT54), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n835), .A2(new_n854), .A3(KEYINPUT53), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n856), .A2(new_n864), .A3(new_n869), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n872), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n784), .A2(new_n686), .A3(new_n786), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT114), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT114), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n784), .A2(new_n786), .A3(new_n881), .A4(new_n686), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n789), .A2(new_n733), .A3(new_n736), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT116), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n887), .B(new_n884), .C1(new_n880), .C2(new_n882), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n830), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n263), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n631), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n715), .A2(new_n891), .A3(new_n884), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n644), .A2(new_n655), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n734), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n811), .A2(new_n813), .B1(new_n412), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n762), .A2(new_n631), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n897), .B(new_n768), .C1(new_n880), .C2(new_n882), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n737), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n883), .A2(new_n746), .A3(new_n718), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT115), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(KEYINPUT50), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n737), .B(new_n897), .C1(new_n880), .C2(new_n882), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n902), .A2(KEYINPUT50), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n746), .A3(new_n718), .A4(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n889), .A2(new_n899), .A3(new_n903), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT51), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n901), .B(new_n905), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT51), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n889), .A4(new_n899), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n726), .B(new_n913), .C1(new_n886), .C2(new_n888), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n726), .B1(new_n886), .B2(new_n888), .ZN(new_n915));
  NOR2_X1   g729(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n883), .A2(new_n631), .A3(new_n752), .A4(new_n762), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT117), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n262), .A2(G952), .ZN(new_n921));
  INV_X1    g735(.A(new_n656), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n892), .B2(new_n922), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n914), .A2(new_n918), .A3(new_n920), .A4(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n912), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n912), .B2(new_n924), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n818), .B1(new_n878), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n638), .A2(new_n414), .A3(new_n664), .A4(new_n655), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT109), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n895), .A2(KEYINPUT49), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT49), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n718), .B1(new_n933), .B2(new_n734), .ZN(new_n934));
  NOR4_X1   g748(.A1(new_n931), .A2(new_n715), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT120), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n873), .A2(new_n876), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT54), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n912), .A2(new_n924), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT119), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n856), .A2(new_n864), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n850), .A2(new_n851), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT113), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n850), .A2(KEYINPUT113), .A3(new_n851), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n875), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n835), .A2(KEYINPUT53), .A3(new_n869), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n948), .A3(new_n872), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n912), .A2(new_n924), .A3(new_n925), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n938), .A2(new_n940), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n818), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n935), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT120), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n936), .A2(new_n955), .ZN(G75));
  NOR2_X1   g770(.A1(new_n855), .A2(new_n870), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n293), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(G210), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT56), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n490), .B(new_n492), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT55), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n959), .B2(new_n960), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n262), .A2(G952), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(G51));
  NOR3_X1   g780(.A1(new_n957), .A2(new_n293), .A3(new_n794), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n795), .B(KEYINPUT57), .Z(new_n968));
  AOI21_X1  g782(.A(new_n872), .B1(new_n947), .B2(new_n948), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n968), .B1(new_n871), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n405), .A2(new_n406), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT121), .B1(new_n972), .B2(new_n965), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT121), .ZN(new_n974));
  INV_X1    g788(.A(new_n965), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT54), .B1(new_n855), .B2(new_n870), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n949), .ZN(new_n977));
  AOI22_X1  g791(.A1(new_n977), .A2(new_n968), .B1(new_n405), .B2(new_n406), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n974), .B(new_n975), .C1(new_n978), .C2(new_n967), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n973), .A2(new_n979), .ZN(G54));
  NAND3_X1  g794(.A1(new_n958), .A2(KEYINPUT58), .A3(G475), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(new_n253), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n253), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n982), .A2(new_n983), .A3(new_n965), .ZN(G60));
  NAND2_X1  g798(.A1(G478), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT59), .Z(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n650), .A2(new_n651), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT122), .Z(new_n989));
  NAND3_X1  g803(.A1(new_n977), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n878), .A2(new_n986), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n975), .B(new_n990), .C1(new_n991), .C2(new_n989), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(G63));
  NAND2_X1  g807(.A1(G217), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT60), .Z(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n855), .B2(new_n870), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(new_n693), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n996), .B1(new_n696), .B2(new_n616), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n975), .A3(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT61), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(G66));
  NOR2_X1   g815(.A1(new_n864), .A2(G953), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT123), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n262), .B1(new_n264), .B2(G224), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT124), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(KEYINPUT125), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT125), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1003), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n747), .B(new_n488), .C1(G898), .C2(new_n262), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1010), .B(new_n1012), .ZN(G69));
  OAI21_X1  g827(.A(new_n726), .B1(new_n922), .B2(new_n825), .ZN(new_n1014));
  OR3_X1    g828(.A1(new_n1014), .A2(new_n706), .A3(new_n768), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n804), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n720), .ZN(new_n1018));
  AOI21_X1  g832(.A(KEYINPUT62), .B1(new_n1018), .B2(new_n865), .ZN(new_n1019));
  INV_X1    g833(.A(new_n865), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT62), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n720), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n816), .B(new_n1017), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n262), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n225), .A2(new_n202), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1027), .B(KEYINPUT126), .Z(new_n1028));
  NAND2_X1  g842(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT127), .ZN(new_n1030));
  NAND2_X1  g844(.A1(G900), .A2(G953), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n772), .A2(new_n865), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n1032), .A2(new_n816), .ZN(new_n1033));
  AOI22_X1  g847(.A1(new_n788), .A2(new_n789), .B1(new_n726), .B2(new_n840), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n1033), .B(new_n779), .C1(new_n802), .C2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1031), .B(new_n1027), .C1(new_n1035), .C2(G953), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1029), .A2(new_n1030), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1037), .B(new_n1038), .ZN(G72));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1040), .B(KEYINPUT63), .Z(new_n1041));
  OAI21_X1  g855(.A(new_n1041), .B1(new_n1023), .B2(new_n829), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1042), .A2(new_n536), .A3(new_n574), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1041), .B1(new_n1035), .B2(new_n829), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1044), .A2(new_n548), .A3(new_n537), .A4(new_n547), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n575), .A2(new_n552), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n937), .A2(new_n1041), .A3(new_n1046), .ZN(new_n1047));
  AND4_X1   g861(.A1(new_n975), .A2(new_n1043), .A3(new_n1045), .A4(new_n1047), .ZN(G57));
endmodule


