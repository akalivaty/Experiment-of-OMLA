//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n187), .A2(new_n188), .A3(G953), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT94), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G122), .ZN(new_n193));
  INV_X1    g007(.A(G122), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT94), .A3(G116), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(G122), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT95), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT95), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n200), .A3(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n197), .A2(KEYINPUT14), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n197), .A2(KEYINPUT14), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n196), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT70), .B(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT96), .B1(new_n211), .B2(G143), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT96), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G134), .ZN(new_n218));
  INV_X1    g032(.A(G134), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n219), .A3(new_n216), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n204), .A2(KEYINPUT98), .A3(new_n208), .A4(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT98), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n210), .A2(new_n219), .A3(new_n216), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n219), .B1(new_n210), .B2(new_n216), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n208), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(G107), .B1(new_n199), .B2(new_n201), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT99), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT97), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n220), .B(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT13), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n216), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n210), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n216), .A2(new_n233), .ZN(new_n236));
  OAI21_X1  g050(.A(G134), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n202), .A2(new_n203), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n232), .B(new_n237), .C1(new_n238), .C2(new_n227), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n229), .A2(new_n230), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n230), .B1(new_n229), .B2(new_n239), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n190), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n229), .A2(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT99), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n229), .A2(new_n230), .A3(new_n239), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n189), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G902), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G478), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT15), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n251), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n248), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(G210), .B1(G237), .B2(G902), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n214), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n263), .A2(new_n264), .A3(new_n211), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n209), .B1(new_n259), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n214), .A2(G146), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n258), .B2(G143), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n214), .A2(KEYINPUT65), .A3(G146), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n266), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G125), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n259), .A2(new_n260), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n271), .A2(new_n272), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n259), .ZN(new_n281));
  NOR2_X1   g095(.A1(KEYINPUT0), .A2(G128), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G125), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT90), .ZN(new_n287));
  INV_X1    g101(.A(G224), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(G953), .ZN(new_n289));
  INV_X1    g103(.A(G953), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT90), .A3(G224), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(KEYINPUT91), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n286), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n295));
  XNOR2_X1  g109(.A(G116), .B(G119), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT2), .B(G113), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n298), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(KEYINPUT71), .A3(new_n296), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n192), .A2(G119), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT5), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(G113), .B(new_n305), .C1(new_n297), .C2(new_n304), .ZN(new_n306));
  INV_X1    g120(.A(G104), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G107), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n203), .A2(G104), .ZN(new_n309));
  OAI21_X1  g123(.A(G101), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT3), .B1(new_n307), .B2(G107), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n203), .A3(G104), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n307), .A2(G107), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT84), .B(G101), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n310), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n317), .A2(KEYINPUT85), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT85), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n310), .B(new_n319), .C1(new_n315), .C2(new_n316), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n302), .B(new_n306), .C1(new_n318), .C2(new_n321), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n297), .A2(new_n295), .A3(new_n298), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT71), .B1(new_n300), .B2(new_n296), .ZN(new_n324));
  OAI22_X1  g138(.A1(new_n323), .A2(new_n324), .B1(new_n296), .B2(new_n300), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n315), .A2(new_n316), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n315), .A2(G101), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT4), .B1(new_n315), .B2(G101), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n325), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G110), .B(G122), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n322), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT6), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n322), .A2(new_n331), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n332), .B(KEYINPUT89), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(KEYINPUT6), .A3(new_n336), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n294), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n302), .A2(new_n306), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n317), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n332), .B(KEYINPUT8), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n291), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n286), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n276), .A2(new_n285), .A3(new_n347), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n333), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n248), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n257), .B1(new_n340), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n351), .ZN(new_n354));
  AOI21_X1  g168(.A(G902), .B1(new_n354), .B2(new_n345), .ZN(new_n355));
  INV_X1    g169(.A(new_n294), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n333), .A2(KEYINPUT6), .B1(new_n335), .B2(new_n336), .ZN(new_n357));
  INV_X1    g171(.A(new_n339), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n359), .A3(new_n256), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(G214), .B1(G237), .B2(G902), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT16), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G125), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G125), .B(G140), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n275), .A2(KEYINPUT77), .A3(G140), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n369), .B1(new_n374), .B2(new_n364), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n258), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n373), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n368), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G146), .ZN(new_n379));
  NOR2_X1   g193(.A1(G237), .A2(G953), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G214), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(new_n214), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT17), .A3(G131), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(G131), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n381), .B(G143), .ZN(new_n385));
  INV_X1    g199(.A(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT17), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n376), .A2(new_n379), .A3(new_n383), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n374), .A2(G146), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n370), .A2(new_n258), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT18), .A2(G131), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n391), .A2(new_n392), .B1(new_n385), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n382), .A2(KEYINPUT18), .A3(G131), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT92), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G113), .B(G122), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n307), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n377), .A2(KEYINPUT19), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(KEYINPUT19), .B2(new_n370), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n405), .A2(new_n258), .B1(new_n384), .B2(new_n387), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n379), .A2(KEYINPUT79), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n378), .A2(new_n408), .A3(G146), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n402), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n399), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(G475), .A2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT20), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n403), .A2(new_n412), .A3(new_n417), .A4(new_n414), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n400), .B1(new_n419), .B2(new_n402), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n390), .A2(new_n399), .A3(KEYINPUT93), .A4(new_n411), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n248), .A3(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n416), .A2(new_n418), .B1(G475), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G952), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(G953), .ZN(new_n425));
  NAND2_X1  g239(.A1(G234), .A2(G237), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(G898), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(G902), .A3(G953), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT100), .Z(new_n432));
  NAND2_X1  g246(.A1(new_n423), .A2(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n255), .A2(new_n363), .A3(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT10), .B(new_n274), .C1(new_n318), .C2(new_n321), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n284), .B1(new_n329), .B2(new_n330), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n211), .B1(new_n259), .B2(KEYINPUT1), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n266), .B1(new_n262), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n327), .A3(new_n310), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT10), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n435), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n443), .A2(KEYINPUT11), .B1(new_n219), .B2(G137), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n445));
  INV_X1    g259(.A(G137), .ZN(new_n446));
  AND4_X1   g260(.A1(KEYINPUT67), .A2(new_n445), .A3(new_n446), .A4(G134), .ZN(new_n447));
  AOI22_X1  g261(.A1(KEYINPUT67), .A2(new_n445), .B1(new_n446), .B2(G134), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G131), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n386), .B(new_n444), .C1(new_n447), .C2(new_n448), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n442), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G140), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n290), .A2(G227), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT88), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n442), .A2(new_n452), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n453), .B2(new_n456), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n317), .A2(KEYINPUT85), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n259), .B1(new_n263), .B2(new_n264), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n211), .A2(KEYINPUT70), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT70), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G128), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n281), .A2(new_n469), .B1(new_n262), .B2(new_n265), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n470), .A3(new_n320), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT86), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n463), .A2(new_n470), .A3(new_n473), .A4(new_n320), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n439), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n452), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT87), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n475), .A2(new_n479), .A3(KEYINPUT12), .A4(new_n452), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n477), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n453), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n456), .ZN(new_n485));
  OAI211_X1 g299(.A(G469), .B(new_n462), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n482), .A2(new_n457), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n459), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n456), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G469), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n248), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n248), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n486), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n434), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(G472), .A2(G902), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n498), .A2(KEYINPUT32), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n501));
  INV_X1    g315(.A(G210), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n502), .A2(G237), .A3(G953), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n501), .B(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT26), .B(G101), .Z(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n446), .A2(G134), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n219), .A2(G137), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n386), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI22_X1  g323(.A1(KEYINPUT67), .A2(new_n445), .B1(new_n446), .B2(G134), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n443), .A2(KEYINPUT11), .B1(new_n219), .B2(G137), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT67), .A4(G134), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n509), .B1(new_n513), .B2(new_n386), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n452), .A2(new_n284), .B1(new_n274), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n299), .A2(new_n301), .B1(new_n297), .B2(new_n298), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n506), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n518));
  INV_X1    g332(.A(new_n509), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n451), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT68), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT68), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n451), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n523), .A3(new_n274), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n277), .A2(new_n282), .ZN(new_n525));
  OAI211_X1 g339(.A(KEYINPUT66), .B(new_n278), .C1(new_n273), .C2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n278), .B1(new_n273), .B2(new_n525), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT66), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n452), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n518), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n451), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n511), .A2(new_n512), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n386), .B1(new_n533), .B2(new_n444), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n284), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n259), .A2(new_n280), .B1(new_n464), .B2(new_n468), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n261), .A2(new_n267), .A3(new_n211), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n451), .B(new_n519), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n538), .A3(KEYINPUT30), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n325), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n517), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n517), .B(KEYINPUT73), .C1(new_n531), .C2(new_n540), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(KEYINPUT31), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n516), .B1(new_n524), .B2(new_n530), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n535), .A2(new_n538), .A3(new_n516), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT28), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n470), .A2(new_n520), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n527), .B1(new_n450), .B2(new_n451), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT74), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT74), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n535), .A2(new_n538), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n516), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT28), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n506), .ZN(new_n559));
  INV_X1    g373(.A(new_n506), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n547), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n524), .A2(new_n530), .ZN(new_n562));
  INV_X1    g376(.A(new_n518), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n516), .B1(new_n515), .B2(KEYINPUT30), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT31), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND4_X1   g382(.A1(new_n500), .A2(new_n545), .A3(new_n559), .A4(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n558), .A2(new_n506), .B1(new_n567), .B2(new_n566), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n500), .B1(new_n570), .B2(new_n545), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n499), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n564), .A2(new_n565), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n547), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n506), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT29), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n575), .B(new_n576), .C1(new_n506), .C2(new_n558), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n325), .B1(new_n550), .B2(new_n551), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n547), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT28), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n557), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n506), .A2(new_n576), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G472), .ZN(new_n585));
  INV_X1    g399(.A(new_n498), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n545), .A2(new_n559), .A3(new_n568), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT75), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n570), .A2(new_n500), .A3(new_n545), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n572), .B(new_n585), .C1(new_n590), .C2(KEYINPUT32), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT83), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n376), .A2(new_n379), .ZN(new_n593));
  INV_X1    g407(.A(G119), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G128), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n468), .B2(new_n594), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT24), .B(G110), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n599));
  AND2_X1   g413(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n600));
  NOR2_X1   g414(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n601));
  OAI22_X1  g415(.A1(new_n600), .A2(new_n601), .B1(new_n594), .B2(G128), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n599), .A2(new_n595), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G110), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n593), .A2(new_n598), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n596), .A2(new_n597), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n407), .A2(new_n409), .A3(new_n392), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT22), .B(G137), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n290), .A2(G221), .A3(G234), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT80), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n606), .A2(new_n610), .A3(new_n614), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT82), .ZN(new_n619));
  INV_X1    g433(.A(G234), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n620), .B2(G217), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT81), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT25), .ZN(new_n623));
  AOI21_X1  g437(.A(G902), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n616), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G217), .B1(new_n620), .B2(G902), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n625), .B2(new_n626), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n619), .A2(new_n621), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n591), .A2(new_n592), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n592), .B1(new_n591), .B2(new_n630), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n497), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n316), .ZN(G3));
  AOI21_X1  g448(.A(G902), .B1(new_n588), .B2(new_n589), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n590), .B1(new_n636), .B2(G472), .ZN(new_n637));
  INV_X1    g451(.A(new_n496), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n482), .A2(new_n457), .B1(new_n456), .B2(new_n488), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(G902), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n493), .B1(new_n640), .B2(new_n491), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n638), .B1(new_n641), .B2(new_n486), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n637), .A2(new_n642), .A3(new_n630), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n250), .A2(G902), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT33), .B1(new_n247), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  AOI211_X1 g461(.A(KEYINPUT101), .B(new_n647), .C1(new_n242), .C2(new_n246), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n644), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n249), .A2(new_n250), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n423), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n362), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n353), .B2(new_n360), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n651), .A2(new_n432), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n643), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT34), .B(G104), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  INV_X1    g471(.A(new_n433), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n255), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n659), .A2(KEYINPUT102), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(KEYINPUT102), .ZN(new_n661));
  NOR4_X1   g475(.A1(new_n643), .A2(new_n660), .A3(new_n363), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT103), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT35), .B(G107), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  OAI21_X1  g479(.A(new_n498), .B1(new_n569), .B2(new_n571), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n627), .A2(new_n629), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n615), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n611), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n621), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(G472), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n666), .B(new_n671), .C1(new_n635), .C2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT104), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT104), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n497), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  INV_X1    g492(.A(new_n423), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n430), .A2(G900), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n427), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n683), .A2(new_n255), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n671), .A2(new_n653), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n642), .A2(new_n684), .A3(new_n591), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  NAND2_X1  g502(.A1(new_n495), .A2(new_n496), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n681), .B(KEYINPUT39), .Z(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT105), .Z(new_n692));
  INV_X1    g506(.A(KEYINPUT40), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n255), .A2(new_n679), .A3(new_n362), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n543), .A2(new_n544), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n506), .B2(new_n579), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n698), .B2(G902), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n572), .B(new_n699), .C1(new_n590), .C2(KEYINPUT32), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n361), .B(KEYINPUT38), .Z(new_n702));
  NOR4_X1   g516(.A1(new_n696), .A2(new_n701), .A3(new_n671), .A4(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n694), .A2(new_n695), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  AOI211_X1 g519(.A(new_n423), .B(new_n682), .C1(new_n649), .C2(new_n650), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n591), .A3(new_n642), .A4(new_n686), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  NAND2_X1  g522(.A1(new_n588), .A2(new_n589), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT32), .B1(new_n709), .B2(new_n498), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n572), .A2(new_n585), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n630), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n649), .A2(new_n650), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n679), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n653), .A2(new_n432), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(G469), .B1(new_n639), .B2(G902), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n492), .A2(new_n718), .A3(new_n496), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n713), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  NOR2_X1   g537(.A1(new_n660), .A2(new_n661), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n719), .A2(new_n363), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n713), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NOR2_X1   g541(.A1(new_n685), .A2(new_n719), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n255), .A2(new_n433), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n591), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  NAND3_X1  g545(.A1(new_n255), .A2(new_n679), .A3(new_n653), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n733), .A2(new_n432), .A3(new_n720), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n635), .A2(new_n672), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n581), .A2(KEYINPUT106), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n581), .A2(KEYINPUT106), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n506), .A3(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n545), .A2(new_n568), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n586), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n734), .A2(new_n630), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND3_X1  g557(.A1(new_n706), .A2(new_n741), .A3(new_n728), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  NOR2_X1   g559(.A1(new_n361), .A2(new_n652), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n689), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n713), .A2(new_n748), .A3(new_n706), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  XNOR2_X1  g566(.A(new_n684), .B(KEYINPUT107), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n713), .A3(new_n748), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  XNOR2_X1  g569(.A(new_n423), .B(KEYINPUT109), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n714), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n679), .B1(new_n649), .B2(new_n650), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n757), .B(KEYINPUT43), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n759), .B2(KEYINPUT108), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n671), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n637), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n747), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n462), .B1(new_n484), .B2(new_n485), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT45), .B(new_n462), .C1(new_n484), .C2(new_n485), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(G469), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n494), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT46), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n774), .A2(new_n775), .B1(new_n491), .B2(new_n640), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n494), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n778), .A2(new_n638), .A3(new_n690), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n768), .B(new_n779), .C1(new_n767), .C2(new_n766), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n778), .B2(new_n638), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n776), .A2(new_n777), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n496), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n706), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n787), .A2(new_n591), .A3(new_n630), .A4(new_n747), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g603(.A(KEYINPUT110), .B(G140), .Z(new_n790));
  XNOR2_X1  g604(.A(new_n789), .B(new_n790), .ZN(G42));
  INV_X1    g605(.A(new_n741), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n252), .A2(KEYINPUT113), .A3(new_n254), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n253), .B1(new_n247), .B2(new_n248), .ZN(new_n796));
  AOI211_X1 g610(.A(G902), .B(new_n251), .C1(new_n242), .C2(new_n246), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n591), .A2(new_n683), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n671), .B(new_n748), .C1(new_n793), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n754), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n707), .A2(new_n687), .A3(new_n744), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n732), .A2(new_n682), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n642), .A3(new_n764), .A4(new_n700), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(KEYINPUT52), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n707), .A2(new_n804), .A3(new_n744), .A4(new_n687), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n801), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n749), .B(KEYINPUT42), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n726), .A2(new_n742), .A3(new_n721), .A4(new_n730), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n679), .B(new_n716), .C1(new_n794), .C2(new_n798), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n630), .A3(new_n642), .A4(new_n637), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n676), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n717), .A2(new_n630), .A3(new_n642), .A4(new_n637), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n633), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n633), .A2(new_n816), .A3(KEYINPUT112), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT114), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n642), .A2(new_n434), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n712), .A2(KEYINPUT83), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n591), .A2(new_n592), .A3(new_n630), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n818), .B1(new_n825), .B2(new_n655), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n676), .A2(new_n814), .ZN(new_n827));
  AND4_X1   g641(.A1(KEYINPUT114), .A2(new_n826), .A3(new_n820), .A4(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n809), .B(new_n812), .C1(new_n821), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n744), .A2(new_n687), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(KEYINPUT53), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n811), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n751), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n826), .A2(new_n820), .A3(new_n827), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT114), .A4(new_n820), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n841), .B2(new_n809), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT54), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n829), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n839), .A2(new_n840), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n810), .B2(new_n811), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n835), .A2(new_n751), .A3(KEYINPUT115), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n832), .A2(new_n844), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n846), .A2(new_n850), .A3(new_n809), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n845), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n630), .A2(new_n741), .A3(new_n426), .A4(new_n425), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n763), .A2(new_n725), .A3(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n719), .A2(new_n747), .A3(new_n427), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n701), .A3(new_n630), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n856), .B(new_n425), .C1(new_n715), .C2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n763), .A2(new_n713), .A3(new_n857), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n492), .A2(new_n718), .A3(new_n638), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n783), .A2(new_n785), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n763), .A2(new_n746), .A3(new_n855), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n792), .A2(new_n764), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n763), .A2(new_n857), .A3(new_n868), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n858), .A2(new_n679), .A3(new_n714), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n702), .A2(new_n720), .A3(new_n652), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n855), .A2(new_n762), .A3(new_n760), .A4(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT50), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n873), .A2(new_n874), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n871), .B(KEYINPUT51), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n863), .B1(new_n867), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n865), .A2(new_n866), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT116), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n869), .A2(new_n870), .ZN(new_n884));
  INV_X1    g698(.A(new_n877), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n884), .B1(new_n885), .B2(new_n875), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n879), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n843), .A2(new_n854), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n424), .A2(new_n290), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n702), .A2(new_n630), .A3(new_n496), .A4(new_n362), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n492), .A2(new_n718), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT49), .ZN(new_n895));
  NOR4_X1   g709(.A1(new_n893), .A2(new_n895), .A3(new_n700), .A4(new_n757), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT111), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT117), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n892), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(G75));
  NAND2_X1  g716(.A1(new_n845), .A2(new_n852), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(G210), .A3(G902), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n357), .A2(new_n358), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n294), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n359), .ZN(new_n909));
  XOR2_X1   g723(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n904), .A2(new_n905), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n290), .A2(G952), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT121), .Z(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n904), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n919), .B2(new_n911), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n915), .A2(new_n920), .ZN(G51));
  XNOR2_X1  g735(.A(new_n903), .B(new_n853), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n493), .B(KEYINPUT57), .Z(new_n923));
  OAI21_X1  g737(.A(new_n490), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n773), .B(KEYINPUT122), .Z(new_n925));
  NAND3_X1  g739(.A1(new_n903), .A2(G902), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n916), .B1(new_n924), .B2(new_n926), .ZN(G54));
  NAND2_X1  g741(.A1(KEYINPUT58), .A2(G475), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT123), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n903), .A2(G902), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n413), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n413), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n916), .ZN(G60));
  INV_X1    g747(.A(new_n646), .ZN(new_n934));
  INV_X1    g748(.A(new_n648), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT59), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n917), .B1(new_n922), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n843), .B2(new_n854), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n936), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n941), .A2(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  NAND3_X1  g760(.A1(new_n903), .A2(new_n669), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n903), .A2(new_n946), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n917), .B(new_n947), .C1(new_n948), .C2(new_n619), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G66));
  OAI21_X1  g765(.A(G953), .B1(new_n428), .B2(new_n288), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n846), .A2(new_n835), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n952), .B1(new_n954), .B2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n907), .B1(G898), .B2(new_n290), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  NAND2_X1  g771(.A1(new_n564), .A2(new_n539), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n405), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n704), .A2(new_n960), .A3(new_n802), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n794), .A2(new_n798), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n423), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n747), .B1(new_n963), .B2(new_n715), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n692), .B(new_n964), .C1(new_n632), .C2(new_n631), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n780), .A2(new_n789), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n960), .B1(new_n704), .B2(new_n802), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n961), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n959), .B1(new_n968), .B2(G953), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n959), .B1(G900), .B2(G953), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n779), .A2(new_n713), .A3(new_n733), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n751), .A2(new_n754), .A3(new_n802), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n780), .A2(new_n789), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n970), .B1(new_n973), .B2(G953), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n969), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n290), .B1(G227), .B2(G900), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(KEYINPUT124), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n969), .A2(new_n974), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT125), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(new_n968), .A2(new_n954), .ZN(new_n986));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  AOI22_X1  g802(.A1(new_n986), .A2(new_n988), .B1(new_n573), .B2(new_n547), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n973), .A2(new_n953), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n560), .B1(new_n990), .B2(new_n988), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n575), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n845), .B1(new_n829), .B2(new_n833), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n575), .A2(new_n543), .A3(new_n544), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n988), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n916), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n992), .A2(new_n997), .ZN(G57));
endmodule


