

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738;

  AND2_X1 U368 ( .A1(n735), .A2(n365), .ZN(n374) );
  INV_X1 U369 ( .A(G953), .ZN(n684) );
  XOR2_X1 U370 ( .A(n518), .B(n534), .Z(n349) );
  INV_X1 U371 ( .A(n653), .ZN(n606) );
  NOR2_X2 U372 ( .A1(n738), .A2(n737), .ZN(n546) );
  XNOR2_X2 U373 ( .A(n389), .B(KEYINPUT78), .ZN(n650) );
  XNOR2_X2 U374 ( .A(n589), .B(n354), .ZN(n602) );
  XNOR2_X2 U375 ( .A(n581), .B(n392), .ZN(n685) );
  INV_X2 U376 ( .A(G143), .ZN(n515) );
  NOR2_X1 U377 ( .A1(n608), .A2(n662), .ZN(n609) );
  XNOR2_X1 U378 ( .A(n547), .B(KEYINPUT1), .ZN(n653) );
  INV_X1 U379 ( .A(KEYINPUT30), .ZN(n347) );
  NOR2_X1 U380 ( .A1(n414), .A2(n614), .ZN(n615) );
  XNOR2_X1 U381 ( .A(n439), .B(n612), .ZN(n414) );
  XNOR2_X1 U382 ( .A(n510), .B(n509), .ZN(n547) );
  AND2_X1 U383 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X1 U384 ( .A(n422), .B(n421), .ZN(n556) );
  XNOR2_X1 U385 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U386 ( .A(n446), .B(G104), .ZN(n505) );
  INV_X2 U387 ( .A(G113), .ZN(n444) );
  INV_X2 U388 ( .A(G116), .ZN(n443) );
  XNOR2_X1 U389 ( .A(n387), .B(n347), .ZN(n346) );
  NOR2_X1 U390 ( .A1(n622), .A2(G902), .ZN(n476) );
  XNOR2_X1 U391 ( .A(n507), .B(n475), .ZN(n622) );
  NAND2_X1 U392 ( .A1(n512), .A2(n613), .ZN(n513) );
  XNOR2_X2 U393 ( .A(n513), .B(n350), .ZN(n574) );
  NAND2_X2 U394 ( .A1(n555), .A2(n668), .ZN(n543) );
  NOR2_X2 U395 ( .A1(n728), .A2(n395), .ZN(n647) );
  XNOR2_X1 U396 ( .A(n386), .B(n456), .ZN(n467) );
  XNOR2_X1 U397 ( .A(n465), .B(G137), .ZN(n430) );
  INV_X1 U398 ( .A(KEYINPUT70), .ZN(n465) );
  INV_X1 U399 ( .A(KEYINPUT87), .ZN(n407) );
  INV_X1 U400 ( .A(KEYINPUT44), .ZN(n390) );
  BUF_X1 U401 ( .A(n414), .Z(n395) );
  XNOR2_X1 U402 ( .A(n522), .B(n454), .ZN(n523) );
  XNOR2_X1 U403 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n519) );
  XNOR2_X1 U404 ( .A(n396), .B(n376), .ZN(n668) );
  XNOR2_X1 U405 ( .A(KEYINPUT38), .B(KEYINPUT77), .ZN(n376) );
  NAND2_X1 U406 ( .A1(n405), .A2(G902), .ZN(n402) );
  INV_X1 U407 ( .A(G902), .ZN(n400) );
  XOR2_X1 U408 ( .A(G140), .B(G107), .Z(n504) );
  XNOR2_X1 U409 ( .A(n467), .B(G146), .ZN(n428) );
  INV_X1 U410 ( .A(G110), .ZN(n446) );
  XNOR2_X1 U411 ( .A(n590), .B(n353), .ZN(n373) );
  XNOR2_X1 U412 ( .A(n528), .B(n527), .ZN(n557) );
  INV_X1 U413 ( .A(n556), .ZN(n554) );
  XNOR2_X1 U414 ( .A(n464), .B(n463), .ZN(n620) );
  XOR2_X1 U415 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n520) );
  INV_X1 U416 ( .A(KEYINPUT76), .ZN(n426) );
  INV_X1 U417 ( .A(KEYINPUT72), .ZN(n423) );
  OR2_X1 U418 ( .A1(G237), .A2(G902), .ZN(n514) );
  XNOR2_X1 U419 ( .A(n491), .B(n490), .ZN(n492) );
  NOR2_X1 U420 ( .A1(G953), .A2(G237), .ZN(n521) );
  INV_X1 U421 ( .A(G134), .ZN(n420) );
  XNOR2_X1 U422 ( .A(G902), .B(KEYINPUT15), .ZN(n613) );
  XNOR2_X1 U423 ( .A(KEYINPUT92), .B(KEYINPUT18), .ZN(n459) );
  INV_X1 U424 ( .A(n458), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n467), .B(n457), .ZN(n458) );
  INV_X1 U426 ( .A(KEYINPUT45), .ZN(n612) );
  OR2_X1 U427 ( .A1(n359), .A2(n404), .ZN(n548) );
  NAND2_X1 U428 ( .A1(n348), .A2(n656), .ZN(n404) );
  XOR2_X1 U429 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n469) );
  XNOR2_X1 U430 ( .A(G116), .B(G113), .ZN(n468) );
  INV_X1 U431 ( .A(KEYINPUT88), .ZN(n397) );
  XNOR2_X1 U432 ( .A(G122), .B(KEYINPUT7), .ZN(n530) );
  XNOR2_X1 U433 ( .A(n524), .B(n383), .ZN(n701) );
  XNOR2_X1 U434 ( .A(n526), .B(n525), .ZN(n383) );
  INV_X1 U435 ( .A(KEYINPUT33), .ZN(n392) );
  XNOR2_X1 U436 ( .A(n413), .B(n431), .ZN(n412) );
  INV_X1 U437 ( .A(KEYINPUT28), .ZN(n431) );
  NOR2_X1 U438 ( .A1(n671), .A2(n670), .ZN(n540) );
  XNOR2_X1 U439 ( .A(KEYINPUT105), .B(G478), .ZN(n421) );
  OR2_X1 U440 ( .A1(n704), .A2(G902), .ZN(n422) );
  XNOR2_X1 U441 ( .A(n488), .B(n489), .ZN(n706) );
  XNOR2_X1 U442 ( .A(n508), .B(n506), .ZN(n394) );
  XNOR2_X1 U443 ( .A(n438), .B(n437), .ZN(n737) );
  XNOR2_X1 U444 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n437) );
  INV_X1 U445 ( .A(KEYINPUT35), .ZN(n370) );
  INV_X1 U446 ( .A(n591), .ZN(n372) );
  NAND2_X1 U447 ( .A1(n597), .A2(n417), .ZN(n416) );
  NOR2_X1 U448 ( .A1(n591), .A2(n409), .ZN(n408) );
  NOR2_X1 U449 ( .A1(n557), .A2(n556), .ZN(n639) );
  INV_X1 U450 ( .A(KEYINPUT107), .ZN(n441) );
  XNOR2_X1 U451 ( .A(n703), .B(n704), .ZN(n393) );
  INV_X1 U452 ( .A(KEYINPUT56), .ZN(n449) );
  OR2_X1 U453 ( .A1(n585), .A2(n499), .ZN(n348) );
  AND2_X1 U454 ( .A1(G210), .A2(n514), .ZN(n350) );
  AND2_X1 U455 ( .A1(n595), .A2(n442), .ZN(n351) );
  XNOR2_X1 U456 ( .A(n494), .B(n492), .ZN(n436) );
  OR2_X1 U457 ( .A1(n672), .A2(KEYINPUT86), .ZN(n352) );
  INV_X1 U458 ( .A(KEYINPUT16), .ZN(n448) );
  XOR2_X1 U459 ( .A(KEYINPUT82), .B(KEYINPUT34), .Z(n353) );
  XOR2_X1 U460 ( .A(n588), .B(KEYINPUT0), .Z(n354) );
  XOR2_X1 U461 ( .A(n622), .B(n621), .Z(n355) );
  XOR2_X1 U462 ( .A(n701), .B(n700), .Z(n356) );
  XOR2_X1 U463 ( .A(KEYINPUT48), .B(KEYINPUT71), .Z(n357) );
  NOR2_X1 U464 ( .A1(n729), .A2(G952), .ZN(n708) );
  INV_X1 U465 ( .A(n708), .ZN(n451) );
  XOR2_X1 U466 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n358) );
  NAND2_X1 U467 ( .A1(n401), .A2(n398), .ZN(n359) );
  NAND2_X1 U468 ( .A1(n401), .A2(n398), .ZN(n655) );
  NAND2_X1 U469 ( .A1(n615), .A2(n364), .ZN(n389) );
  BUF_X1 U470 ( .A(n636), .Z(n360) );
  NOR2_X2 U471 ( .A1(n560), .A2(n415), .ZN(n636) );
  NAND2_X1 U472 ( .A1(n412), .A2(n511), .ZN(n560) );
  INV_X2 U473 ( .A(G125), .ZN(n380) );
  NAND2_X1 U474 ( .A1(n655), .A2(n656), .ZN(n435) );
  NAND2_X1 U475 ( .A1(n470), .A2(n448), .ZN(n362) );
  NAND2_X1 U476 ( .A1(n361), .A2(KEYINPUT16), .ZN(n363) );
  NAND2_X1 U477 ( .A1(n362), .A2(n363), .ZN(n447) );
  INV_X1 U478 ( .A(n470), .ZN(n361) );
  XNOR2_X2 U479 ( .A(n447), .B(n505), .ZN(n445) );
  NOR2_X1 U480 ( .A1(n578), .A2(n577), .ZN(n364) );
  NOR2_X1 U481 ( .A1(n578), .A2(n577), .ZN(n616) );
  XNOR2_X1 U482 ( .A(n434), .B(KEYINPUT79), .ZN(n433) );
  AND2_X2 U483 ( .A1(n555), .A2(n408), .ZN(n635) );
  BUF_X1 U484 ( .A(n574), .Z(n396) );
  INV_X1 U485 ( .A(n736), .ZN(n365) );
  XNOR2_X1 U486 ( .A(n366), .B(KEYINPUT32), .ZN(n736) );
  NOR2_X2 U487 ( .A1(n596), .A2(n416), .ZN(n366) );
  XNOR2_X2 U488 ( .A(n367), .B(n441), .ZN(n735) );
  NAND2_X1 U489 ( .A1(n599), .A2(n351), .ZN(n367) );
  NOR2_X2 U490 ( .A1(n596), .A2(n606), .ZN(n599) );
  XNOR2_X2 U491 ( .A(n369), .B(n368), .ZN(n391) );
  XNOR2_X2 U492 ( .A(n445), .B(n349), .ZN(n369) );
  XNOR2_X1 U493 ( .A(n369), .B(G101), .ZN(n715) );
  NAND2_X1 U494 ( .A1(n374), .A2(n734), .ZN(n377) );
  XNOR2_X2 U495 ( .A(n371), .B(n370), .ZN(n734) );
  NAND2_X1 U496 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U497 ( .A(n375), .B(n357), .ZN(n578) );
  NAND2_X1 U498 ( .A1(n418), .A2(n567), .ZN(n375) );
  XNOR2_X1 U499 ( .A(n377), .B(n390), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n427), .B(n426), .ZN(n425) );
  AND2_X2 U501 ( .A1(n433), .A2(n346), .ZN(n555) );
  NAND2_X1 U502 ( .A1(n379), .A2(n378), .ZN(n590) );
  INV_X1 U503 ( .A(n608), .ZN(n378) );
  INV_X1 U504 ( .A(n685), .ZN(n379) );
  XNOR2_X2 U505 ( .A(n380), .B(G146), .ZN(n485) );
  NAND2_X1 U506 ( .A1(n636), .A2(KEYINPUT47), .ZN(n564) );
  XNOR2_X1 U507 ( .A(n381), .B(n358), .ZN(G60) );
  NAND2_X1 U508 ( .A1(n385), .A2(n451), .ZN(n381) );
  XNOR2_X1 U509 ( .A(n382), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U510 ( .A1(n384), .A2(n451), .ZN(n382) );
  INV_X1 U511 ( .A(n721), .ZN(n386) );
  BUF_X2 U512 ( .A(n699), .Z(n693) );
  XNOR2_X1 U513 ( .A(n623), .B(n355), .ZN(n384) );
  XNOR2_X1 U514 ( .A(n702), .B(n356), .ZN(n385) );
  NAND2_X1 U515 ( .A1(n650), .A2(n617), .ZN(n618) );
  NAND2_X1 U516 ( .A1(n542), .A2(n667), .ZN(n387) );
  NAND2_X1 U517 ( .A1(n388), .A2(n411), .ZN(n427) );
  NOR2_X2 U518 ( .A1(n410), .A2(n406), .ZN(n388) );
  XNOR2_X2 U519 ( .A(n485), .B(G140), .ZN(n486) );
  XNOR2_X1 U520 ( .A(n419), .B(n423), .ZN(n418) );
  NOR2_X2 U521 ( .A1(n619), .A2(n618), .ZN(n699) );
  NAND2_X1 U522 ( .A1(n602), .A2(n593), .ZN(n594) );
  INV_X1 U523 ( .A(n436), .ZN(n405) );
  NAND2_X1 U524 ( .A1(n436), .A2(n400), .ZN(n399) );
  NOR2_X2 U525 ( .A1(n415), .A2(n587), .ZN(n589) );
  XNOR2_X2 U526 ( .A(n428), .B(n720), .ZN(n507) );
  NOR2_X2 U527 ( .A1(n652), .A2(n547), .ZN(n603) );
  NAND2_X1 U528 ( .A1(n575), .A2(n545), .ZN(n438) );
  XNOR2_X2 U529 ( .A(n476), .B(n477), .ZN(n659) );
  INV_X1 U530 ( .A(n602), .ZN(n608) );
  XNOR2_X2 U531 ( .A(n391), .B(n462), .ZN(n512) );
  NOR2_X1 U532 ( .A1(n393), .A2(n708), .ZN(G63) );
  XNOR2_X1 U533 ( .A(n507), .B(n394), .ZN(n695) );
  XNOR2_X1 U534 ( .A(n616), .B(n397), .ZN(n728) );
  OR2_X1 U535 ( .A1(n706), .A2(n399), .ZN(n398) );
  NAND2_X1 U536 ( .A1(n706), .A2(n405), .ZN(n403) );
  XNOR2_X2 U537 ( .A(n635), .B(n407), .ZN(n406) );
  INV_X1 U538 ( .A(n396), .ZN(n409) );
  NAND2_X1 U539 ( .A1(n566), .A2(n352), .ZN(n410) );
  NAND2_X1 U540 ( .A1(n563), .A2(KEYINPUT86), .ZN(n411) );
  NAND2_X1 U541 ( .A1(n432), .A2(n542), .ZN(n413) );
  NOR2_X1 U542 ( .A1(n395), .A2(G953), .ZN(n709) );
  XNOR2_X2 U543 ( .A(n558), .B(n559), .ZN(n415) );
  NOR2_X1 U544 ( .A1(n653), .A2(n359), .ZN(n417) );
  XNOR2_X2 U545 ( .A(n594), .B(KEYINPUT22), .ZN(n596) );
  NAND2_X1 U546 ( .A1(n425), .A2(n424), .ZN(n419) );
  XNOR2_X2 U547 ( .A(n466), .B(n420), .ZN(n533) );
  XNOR2_X2 U548 ( .A(n515), .B(G128), .ZN(n466) );
  INV_X1 U549 ( .A(n643), .ZN(n424) );
  XNOR2_X2 U550 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n721) );
  XNOR2_X2 U551 ( .A(n533), .B(n429), .ZN(n720) );
  XNOR2_X2 U552 ( .A(n516), .B(n430), .ZN(n429) );
  INV_X1 U553 ( .A(n542), .ZN(n595) );
  INV_X1 U554 ( .A(n548), .ZN(n432) );
  NAND2_X1 U555 ( .A1(n603), .A2(n348), .ZN(n434) );
  XNOR2_X2 U556 ( .A(n435), .B(KEYINPUT68), .ZN(n652) );
  XNOR2_X2 U557 ( .A(n543), .B(KEYINPUT39), .ZN(n575) );
  NAND2_X1 U558 ( .A1(n440), .A2(n611), .ZN(n439) );
  NAND2_X1 U559 ( .A1(n574), .A2(n667), .ZN(n558) );
  INV_X1 U560 ( .A(n359), .ZN(n442) );
  XNOR2_X2 U561 ( .A(n443), .B(G107), .ZN(n534) );
  XNOR2_X2 U562 ( .A(n444), .B(G122), .ZN(n518) );
  XNOR2_X1 U563 ( .A(n450), .B(n449), .ZN(G51) );
  NAND2_X1 U564 ( .A1(n452), .A2(n451), .ZN(n450) );
  XNOR2_X1 U565 ( .A(n453), .B(n620), .ZN(n452) );
  NAND2_X1 U566 ( .A1(n699), .A2(G210), .ZN(n453) );
  AND2_X1 U567 ( .A1(G214), .A2(n521), .ZN(n454) );
  OR2_X1 U568 ( .A1(n672), .A2(n610), .ZN(n455) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n485), .B(n461), .ZN(n462) );
  INV_X1 U571 ( .A(KEYINPUT97), .ZN(n490) );
  XNOR2_X1 U572 ( .A(KEYINPUT13), .B(G475), .ZN(n527) );
  XNOR2_X1 U573 ( .A(n697), .B(n696), .ZN(n698) );
  XOR2_X1 U574 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n464) );
  XNOR2_X2 U575 ( .A(G119), .B(KEYINPUT3), .ZN(n470) );
  XNOR2_X1 U576 ( .A(KEYINPUT67), .B(G101), .ZN(n456) );
  XNOR2_X2 U577 ( .A(KEYINPUT64), .B(n684), .ZN(n729) );
  NAND2_X1 U578 ( .A1(G224), .A2(n729), .ZN(n457) );
  XNOR2_X1 U579 ( .A(n466), .B(KEYINPUT17), .ZN(n460) );
  XNOR2_X1 U580 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U581 ( .A(n512), .B(KEYINPUT84), .ZN(n463) );
  XNOR2_X1 U582 ( .A(G472), .B(KEYINPUT75), .ZN(n477) );
  XOR2_X2 U583 ( .A(KEYINPUT69), .B(G131), .Z(n516) );
  XNOR2_X1 U584 ( .A(n469), .B(n468), .ZN(n474) );
  XNOR2_X1 U585 ( .A(n470), .B(KEYINPUT98), .ZN(n472) );
  NAND2_X1 U586 ( .A1(n521), .A2(G210), .ZN(n471) );
  XNOR2_X1 U587 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U588 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U589 ( .A(n659), .B(KEYINPUT106), .ZN(n542) );
  NAND2_X1 U590 ( .A1(n729), .A2(G234), .ZN(n478) );
  XOR2_X1 U591 ( .A(KEYINPUT8), .B(n478), .Z(n529) );
  NAND2_X1 U592 ( .A1(G221), .A2(n529), .ZN(n489) );
  XOR2_X1 U593 ( .A(G110), .B(G119), .Z(n480) );
  XNOR2_X1 U594 ( .A(G137), .B(G128), .ZN(n479) );
  XNOR2_X1 U595 ( .A(n480), .B(n479), .ZN(n484) );
  XOR2_X1 U596 ( .A(KEYINPUT74), .B(KEYINPUT24), .Z(n482) );
  XNOR2_X1 U597 ( .A(KEYINPUT96), .B(KEYINPUT23), .ZN(n481) );
  XNOR2_X1 U598 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U599 ( .A(n484), .B(n483), .Z(n487) );
  XNOR2_X2 U600 ( .A(n486), .B(KEYINPUT10), .ZN(n719) );
  XNOR2_X1 U601 ( .A(n487), .B(n719), .ZN(n488) );
  XNOR2_X1 U602 ( .A(KEYINPUT25), .B(KEYINPUT80), .ZN(n491) );
  NAND2_X1 U603 ( .A1(G234), .A2(n613), .ZN(n493) );
  XNOR2_X1 U604 ( .A(KEYINPUT20), .B(n493), .ZN(n500) );
  NAND2_X1 U605 ( .A1(n500), .A2(G217), .ZN(n494) );
  NAND2_X1 U606 ( .A1(G234), .A2(G237), .ZN(n495) );
  XNOR2_X1 U607 ( .A(n495), .B(KEYINPUT14), .ZN(n496) );
  NAND2_X1 U608 ( .A1(G952), .A2(n496), .ZN(n681) );
  NOR2_X1 U609 ( .A1(G953), .A2(n681), .ZN(n585) );
  NAND2_X1 U610 ( .A1(G902), .A2(n496), .ZN(n583) );
  NOR2_X1 U611 ( .A1(n729), .A2(n583), .ZN(n497) );
  XOR2_X1 U612 ( .A(KEYINPUT108), .B(n497), .Z(n498) );
  NOR2_X1 U613 ( .A1(G900), .A2(n498), .ZN(n499) );
  NAND2_X1 U614 ( .A1(n500), .A2(G221), .ZN(n501) );
  XOR2_X1 U615 ( .A(n501), .B(KEYINPUT21), .Z(n656) );
  XOR2_X1 U616 ( .A(KEYINPUT95), .B(KEYINPUT81), .Z(n503) );
  NAND2_X1 U617 ( .A1(G227), .A2(n729), .ZN(n502) );
  XNOR2_X1 U618 ( .A(n503), .B(n502), .ZN(n508) );
  NOR2_X1 U619 ( .A1(G902), .A2(n695), .ZN(n510) );
  XOR2_X1 U620 ( .A(KEYINPUT73), .B(G469), .Z(n509) );
  INV_X1 U621 ( .A(n547), .ZN(n511) );
  NAND2_X1 U622 ( .A1(G214), .A2(n514), .ZN(n667) );
  NAND2_X1 U623 ( .A1(n668), .A2(n667), .ZN(n671) );
  XNOR2_X1 U624 ( .A(n516), .B(G143), .ZN(n517) );
  XNOR2_X1 U625 ( .A(n517), .B(G104), .ZN(n526) );
  XNOR2_X1 U626 ( .A(n518), .B(KEYINPUT11), .ZN(n525) );
  XNOR2_X1 U627 ( .A(n520), .B(n519), .ZN(n522) );
  XNOR2_X1 U628 ( .A(n719), .B(n523), .ZN(n524) );
  NOR2_X1 U629 ( .A1(G902), .A2(n701), .ZN(n528) );
  INV_X1 U630 ( .A(n557), .ZN(n544) );
  NAND2_X1 U631 ( .A1(n529), .A2(G217), .ZN(n538) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n531) );
  XNOR2_X1 U633 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U634 ( .A(n532), .B(KEYINPUT104), .Z(n536) );
  XNOR2_X1 U635 ( .A(n533), .B(n534), .ZN(n535) );
  XNOR2_X1 U636 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U637 ( .A(n538), .B(n537), .ZN(n704) );
  NAND2_X1 U638 ( .A1(n544), .A2(n556), .ZN(n670) );
  XNOR2_X1 U639 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n539) );
  XNOR2_X1 U640 ( .A(n540), .B(n539), .ZN(n686) );
  NOR2_X1 U641 ( .A1(n560), .A2(n686), .ZN(n541) );
  XNOR2_X1 U642 ( .A(n541), .B(KEYINPUT42), .ZN(n738) );
  NOR2_X1 U643 ( .A1(n554), .A2(n544), .ZN(n545) );
  XNOR2_X1 U644 ( .A(n546), .B(KEYINPUT46), .ZN(n567) );
  XNOR2_X1 U645 ( .A(n659), .B(KEYINPUT6), .ZN(n598) );
  NOR2_X1 U646 ( .A1(n548), .A2(n598), .ZN(n549) );
  XOR2_X1 U647 ( .A(n549), .B(KEYINPUT109), .Z(n550) );
  NAND2_X1 U648 ( .A1(n545), .A2(n550), .ZN(n568) );
  NOR2_X1 U649 ( .A1(n558), .A2(n568), .ZN(n552) );
  XNOR2_X1 U650 ( .A(KEYINPUT113), .B(KEYINPUT36), .ZN(n551) );
  XNOR2_X1 U651 ( .A(n552), .B(n551), .ZN(n553) );
  NOR2_X1 U652 ( .A1(n653), .A2(n553), .ZN(n643) );
  NAND2_X1 U653 ( .A1(n557), .A2(n554), .ZN(n591) );
  NOR2_X1 U654 ( .A1(n545), .A2(n639), .ZN(n672) );
  INV_X1 U655 ( .A(n672), .ZN(n561) );
  INV_X1 U656 ( .A(KEYINPUT19), .ZN(n559) );
  NAND2_X1 U657 ( .A1(n561), .A2(n636), .ZN(n562) );
  XNOR2_X1 U658 ( .A(n562), .B(KEYINPUT47), .ZN(n563) );
  INV_X1 U659 ( .A(KEYINPUT86), .ZN(n565) );
  NAND2_X1 U660 ( .A1(n565), .A2(n564), .ZN(n566) );
  INV_X1 U661 ( .A(n568), .ZN(n569) );
  NAND2_X1 U662 ( .A1(n569), .A2(n667), .ZN(n570) );
  NOR2_X1 U663 ( .A1(n606), .A2(n570), .ZN(n572) );
  XNOR2_X1 U664 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n571) );
  XNOR2_X1 U665 ( .A(n572), .B(n571), .ZN(n573) );
  NOR2_X1 U666 ( .A1(n396), .A2(n573), .ZN(n646) );
  NAND2_X1 U667 ( .A1(n639), .A2(n575), .ZN(n645) );
  INV_X1 U668 ( .A(n645), .ZN(n576) );
  OR2_X1 U669 ( .A1(n646), .A2(n576), .ZN(n577) );
  INV_X1 U670 ( .A(n598), .ZN(n579) );
  INV_X1 U671 ( .A(n652), .ZN(n605) );
  AND2_X1 U672 ( .A1(n579), .A2(n605), .ZN(n580) );
  NAND2_X1 U673 ( .A1(n606), .A2(n580), .ZN(n581) );
  NOR2_X1 U674 ( .A1(n684), .A2(G898), .ZN(n582) );
  XNOR2_X1 U675 ( .A(n582), .B(KEYINPUT93), .ZN(n716) );
  NOR2_X1 U676 ( .A1(n583), .A2(n716), .ZN(n584) );
  NOR2_X1 U677 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U678 ( .A(n586), .B(KEYINPUT94), .ZN(n587) );
  INV_X1 U679 ( .A(KEYINPUT90), .ZN(n588) );
  INV_X1 U680 ( .A(n656), .ZN(n592) );
  NOR2_X1 U681 ( .A1(n670), .A2(n592), .ZN(n593) );
  XOR2_X1 U682 ( .A(n598), .B(KEYINPUT83), .Z(n597) );
  NAND2_X1 U683 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U684 ( .A(KEYINPUT89), .B(n600), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n601), .A2(n359), .ZN(n624) );
  NAND2_X1 U686 ( .A1(n603), .A2(n378), .ZN(n604) );
  NOR2_X1 U687 ( .A1(n659), .A2(n604), .ZN(n627) );
  AND2_X1 U688 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n659), .A2(n607), .ZN(n662) );
  XOR2_X1 U690 ( .A(KEYINPUT31), .B(n609), .Z(n640) );
  NOR2_X1 U691 ( .A1(n627), .A2(n640), .ZN(n610) );
  AND2_X1 U692 ( .A1(n624), .A2(n455), .ZN(n611) );
  NOR2_X1 U693 ( .A1(n647), .A2(KEYINPUT2), .ZN(n619) );
  INV_X1 U694 ( .A(n613), .ZN(n617) );
  INV_X1 U695 ( .A(KEYINPUT2), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n699), .A2(G472), .ZN(n623) );
  XOR2_X1 U697 ( .A(KEYINPUT62), .B(KEYINPUT91), .Z(n621) );
  XNOR2_X1 U698 ( .A(G101), .B(KEYINPUT114), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n625), .B(n624), .ZN(G3) );
  NAND2_X1 U700 ( .A1(n627), .A2(n545), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n626), .B(G104), .ZN(G6) );
  XOR2_X1 U702 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n629) );
  NAND2_X1 U703 ( .A1(n627), .A2(n639), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n629), .B(n628), .ZN(n631) );
  XOR2_X1 U705 ( .A(G107), .B(KEYINPUT27), .Z(n630) );
  XNOR2_X1 U706 ( .A(n631), .B(n630), .ZN(G9) );
  XOR2_X1 U707 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n633) );
  NAND2_X1 U708 ( .A1(n639), .A2(n360), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U710 ( .A(G128), .B(n634), .ZN(G30) );
  XOR2_X1 U711 ( .A(n635), .B(G143), .Z(G45) );
  NAND2_X1 U712 ( .A1(n360), .A2(n545), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(G146), .ZN(G48) );
  NAND2_X1 U714 ( .A1(n640), .A2(n545), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n638), .B(G113), .ZN(G15) );
  XOR2_X1 U716 ( .A(G116), .B(KEYINPUT117), .Z(n642) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n642), .B(n641), .ZN(G18) );
  XNOR2_X1 U719 ( .A(G125), .B(n643), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n644), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U721 ( .A(G134), .B(n645), .ZN(G36) );
  XOR2_X1 U722 ( .A(G140), .B(n646), .Z(G42) );
  XNOR2_X1 U723 ( .A(KEYINPUT2), .B(KEYINPUT85), .ZN(n649) );
  INV_X1 U724 ( .A(n647), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n690) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT50), .ZN(n661) );
  NOR2_X1 U729 ( .A1(n656), .A2(n359), .ZN(n657) );
  XOR2_X1 U730 ( .A(KEYINPUT49), .B(n657), .Z(n658) );
  NOR2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U733 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT118), .ZN(n665) );
  XNOR2_X1 U735 ( .A(KEYINPUT51), .B(n665), .ZN(n666) );
  NOR2_X1 U736 ( .A1(n686), .A2(n666), .ZN(n678) );
  NOR2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n675) );
  NOR2_X1 U739 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U740 ( .A(KEYINPUT119), .B(n673), .Z(n674) );
  NOR2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n676), .A2(n685), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U744 ( .A(KEYINPUT52), .B(n679), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U746 ( .A(KEYINPUT120), .B(n682), .Z(n683) );
  NAND2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n688) );
  NOR2_X1 U748 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U751 ( .A(n691), .B(KEYINPUT53), .ZN(n692) );
  XNOR2_X1 U752 ( .A(KEYINPUT121), .B(n692), .ZN(G75) );
  NAND2_X1 U753 ( .A1(n693), .A2(G469), .ZN(n697) );
  XOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  NOR2_X1 U755 ( .A1(n708), .A2(n698), .ZN(G54) );
  NAND2_X1 U756 ( .A1(n699), .A2(G475), .ZN(n702) );
  XOR2_X1 U757 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n700) );
  NAND2_X1 U758 ( .A1(G478), .A2(n693), .ZN(n703) );
  NAND2_X1 U759 ( .A1(G217), .A2(n693), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n705), .B(n706), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n708), .A2(n707), .ZN(G66) );
  XNOR2_X1 U762 ( .A(KEYINPUT123), .B(n709), .ZN(n713) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n710) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n710), .ZN(n711) );
  NAND2_X1 U765 ( .A1(n711), .A2(G898), .ZN(n712) );
  NAND2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n714), .B(KEYINPUT124), .ZN(n718) );
  NAND2_X1 U768 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U769 ( .A(n718), .B(n717), .Z(G69) );
  XNOR2_X1 U770 ( .A(n719), .B(n720), .ZN(n722) );
  XOR2_X1 U771 ( .A(n722), .B(n721), .Z(n726) );
  XOR2_X1 U772 ( .A(G227), .B(n726), .Z(n723) );
  NAND2_X1 U773 ( .A1(n723), .A2(G900), .ZN(n724) );
  NAND2_X1 U774 ( .A1(G953), .A2(n724), .ZN(n725) );
  XNOR2_X1 U775 ( .A(n725), .B(KEYINPUT126), .ZN(n732) );
  XNOR2_X1 U776 ( .A(KEYINPUT125), .B(n726), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U780 ( .A(KEYINPUT127), .B(n733), .Z(G72) );
  XNOR2_X1 U781 ( .A(n734), .B(G122), .ZN(G24) );
  XNOR2_X1 U782 ( .A(n735), .B(G110), .ZN(G12) );
  XOR2_X1 U783 ( .A(G119), .B(n736), .Z(G21) );
  XOR2_X1 U784 ( .A(G131), .B(n737), .Z(G33) );
  XOR2_X1 U785 ( .A(n738), .B(G137), .Z(G39) );
endmodule

