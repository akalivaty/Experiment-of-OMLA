//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT97), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  MUX2_X1   g007(.A(new_n207), .B(KEYINPUT14), .S(new_n208), .Z(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  INV_X1    g012(.A(G50gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(KEYINPUT91), .B(G43gat), .Z(new_n216));
  AOI211_X1 g015(.A(KEYINPUT15), .B(new_n215), .C1(new_n216), .C2(new_n214), .ZN(new_n217));
  INV_X1    g016(.A(new_n211), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n212), .B1(new_n219), .B2(new_n209), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT17), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT95), .ZN(new_n222));
  INV_X1    g021(.A(G85gat), .ZN(new_n223));
  INV_X1    g022(.A(G92gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(KEYINPUT8), .A2(new_n228), .B1(new_n223), .B2(new_n224), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n222), .B(new_n230), .C1(new_n223), .C2(new_n224), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G99gat), .ZN(new_n233));
  INV_X1    g032(.A(G106gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n228), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n227), .A2(new_n237), .A3(new_n229), .A4(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT96), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n220), .A2(KEYINPUT17), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n221), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT41), .ZN(new_n243));
  INV_X1    g042(.A(G232gat), .ZN(new_n244));
  INV_X1    g043(.A(G233gat), .ZN(new_n245));
  NOR3_X1   g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n220), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n232), .B(new_n237), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n204), .B1(new_n242), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT97), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(new_n202), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n242), .A2(KEYINPUT97), .A3(new_n249), .A4(new_n203), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT98), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT98), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(new_n256), .A3(new_n253), .ZN(new_n257));
  XNOR2_X1  g056(.A(G134gat), .B(G162gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n255), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n257), .A2(new_n260), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G15gat), .B(G22gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT16), .ZN(new_n266));
  AOI21_X1  g065(.A(G1gat), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G8gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n265), .A2(KEYINPUT92), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G57gat), .B(G64gat), .Z(new_n272));
  INV_X1    g071(.A(KEYINPUT9), .ZN(new_n273));
  INV_X1    g072(.A(G71gat), .ZN(new_n274));
  INV_X1    g073(.A(G78gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G78gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n272), .A2(new_n278), .A3(new_n276), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT93), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n271), .B1(KEYINPUT21), .B2(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT94), .B(G155gat), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT21), .B1(new_n280), .B2(new_n281), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G127gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n286), .B(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n292));
  XNOR2_X1  g091(.A(G183gat), .B(G211gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n291), .B(new_n294), .Z(new_n295));
  NAND2_X1  g094(.A1(new_n264), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n302), .B1(new_n306), .B2(new_n301), .ZN(new_n307));
  AND2_X1   g106(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT27), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G183gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(new_n312), .A3(G183gat), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n310), .A2(new_n311), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G183gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT27), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n313), .A2(new_n321), .A3(KEYINPUT28), .A4(new_n311), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT71), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT27), .B(G183gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT28), .A4(new_n311), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n307), .B1(new_n319), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT25), .B(new_n299), .C1(new_n300), .C2(KEYINPUT23), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(new_n306), .B2(KEYINPUT23), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n333));
  OR2_X1    g132(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n335));
  AOI21_X1  g134(.A(G190gat), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT24), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n333), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n311), .B1(new_n308), .B2(new_n309), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n342), .A2(KEYINPUT68), .A3(new_n338), .A4(new_n339), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n332), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G169gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT65), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(G176gat), .ZN(new_n347));
  INV_X1    g146(.A(G176gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(KEYINPUT65), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT23), .B(new_n345), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n338), .B(new_n339), .C1(G183gat), .C2(G190gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n299), .ZN(new_n352));
  INV_X1    g151(.A(new_n300), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n351), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT25), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n344), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n344), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n330), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G120gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G113gat), .ZN(new_n364));
  INV_X1    g163(.A(G113gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G120gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368));
  XNOR2_X1  g167(.A(G127gat), .B(G134gat), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n368), .C1(new_n369), .C2(KEYINPUT72), .ZN(new_n370));
  INV_X1    g169(.A(G127gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G134gat), .ZN(new_n372));
  INV_X1    g171(.A(G134gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G127gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n368), .A2(KEYINPUT72), .ZN(new_n376));
  XNOR2_X1  g175(.A(G113gat), .B(G120gat), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n375), .B(new_n376), .C1(new_n377), .C2(KEYINPUT1), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n370), .A2(new_n378), .A3(KEYINPUT73), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n383), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n330), .C1(new_n360), .C2(new_n361), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(KEYINPUT64), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n298), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT34), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n390), .A2(KEYINPUT34), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n384), .A2(new_n386), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n396), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n391), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT33), .B1(new_n387), .B2(new_n390), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT74), .B(G71gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(new_n233), .ZN(new_n402));
  XNOR2_X1  g201(.A(G15gat), .B(G43gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n397), .A2(new_n399), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n397), .B2(new_n399), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n297), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT36), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n400), .A2(new_n404), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n398), .A2(new_n391), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n398), .A2(new_n391), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n406), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT36), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n297), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G141gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G148gat), .ZN(new_n419));
  INV_X1    g218(.A(G148gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G141gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT2), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G155gat), .A2(G162gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n425), .A2(KEYINPUT2), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n420), .A2(KEYINPUT79), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G148gat), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n418), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n419), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n430), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n427), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n425), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT80), .B1(new_n426), .B2(new_n427), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n429), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT81), .B(new_n429), .C1(new_n436), .C2(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT3), .ZN(new_n447));
  NAND2_X1  g246(.A1(G211gat), .A2(G218gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT22), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT76), .ZN(new_n451));
  XNOR2_X1  g250(.A(G197gat), .B(G204gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT76), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n453), .A3(new_n449), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G211gat), .B(G218gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n451), .A2(new_n456), .A3(new_n452), .A4(new_n454), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT29), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n447), .B1(new_n460), .B2(KEYINPUT84), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n459), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n462), .A2(KEYINPUT84), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n446), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G228gat), .A2(G233gat), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n447), .B(new_n429), .C1(new_n436), .C2(new_n441), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n463), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT77), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n458), .A2(KEYINPUT77), .A3(new_n459), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n465), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n442), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n466), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G22gat), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n479), .A2(KEYINPUT85), .ZN(new_n480));
  XOR2_X1   g279(.A(G78gat), .B(G106gat), .Z(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT31), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(new_n214), .ZN(new_n483));
  INV_X1    g282(.A(G22gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n474), .A2(new_n477), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n485), .A2(KEYINPUT85), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n483), .B1(new_n486), .B2(new_n479), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n479), .A2(new_n485), .A3(new_n483), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT86), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n479), .A2(new_n490), .A3(new_n485), .A4(new_n483), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n480), .A2(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n493));
  INV_X1    g292(.A(new_n445), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT79), .B(G148gat), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n419), .B1(new_n495), .B2(new_n418), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n496), .A2(new_n430), .A3(new_n440), .A4(new_n439), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT81), .B1(new_n497), .B2(new_n429), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT3), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n379), .A3(new_n468), .ZN(new_n500));
  XOR2_X1   g299(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(G225gat), .B2(G233gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n442), .A2(new_n503), .A3(new_n379), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n437), .A2(new_n425), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(new_n422), .B2(new_n423), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n432), .A2(G148gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n420), .A2(KEYINPUT79), .ZN(new_n508));
  OAI21_X1  g307(.A(G141gat), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n509), .A2(new_n419), .B1(KEYINPUT2), .B2(new_n425), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n439), .A2(new_n440), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n506), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(new_n381), .A3(new_n382), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n504), .B1(new_n503), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n500), .A2(new_n502), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n442), .A2(new_n379), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n446), .B2(new_n379), .ZN(new_n517));
  NAND2_X1  g316(.A1(G225gat), .A2(G233gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n501), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n512), .A2(new_n381), .A3(KEYINPUT4), .A4(new_n382), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n503), .B1(new_n442), .B2(new_n379), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n379), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n446), .B2(KEYINPUT3), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n522), .B1(new_n524), .B2(new_n468), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n515), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G1gat), .B(G29gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT0), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G57gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n223), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n493), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n531), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n515), .B(new_n530), .C1(new_n519), .C2(new_n525), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n532), .B1(new_n535), .B2(new_n493), .ZN(new_n536));
  NAND2_X1  g335(.A1(G226gat), .A2(G233gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n538), .B(new_n330), .C1(new_n360), .C2(new_n361), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n471), .A2(new_n472), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(KEYINPUT29), .ZN(new_n541));
  INV_X1    g340(.A(new_n329), .ZN(new_n542));
  AOI211_X1 g341(.A(new_n542), .B(new_n307), .C1(new_n319), .C2(new_n327), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n344), .A2(new_n358), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n543), .A2(new_n544), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n362), .A2(new_n541), .B1(new_n547), .B2(new_n538), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n546), .B1(new_n548), .B2(new_n540), .ZN(new_n549));
  XNOR2_X1  g348(.A(G8gat), .B(G36gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT78), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G64gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(new_n224), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n546), .B(new_n553), .C1(new_n548), .C2(new_n540), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(KEYINPUT30), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n549), .A2(new_n558), .A3(new_n554), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n536), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n410), .A2(new_n417), .B1(new_n492), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT88), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n362), .A2(new_n541), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n538), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(new_n540), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n539), .A2(new_n545), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n568), .B(KEYINPUT37), .C1(new_n540), .C2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT38), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n565), .A2(new_n570), .A3(new_n571), .A4(new_n553), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n555), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n563), .B1(new_n536), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n554), .B1(new_n549), .B2(new_n564), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n575), .B1(new_n564), .B2(new_n549), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT38), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n549), .A2(new_n554), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n540), .B1(new_n539), .B2(new_n545), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n540), .B2(new_n548), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT38), .B1(new_n580), .B2(KEYINPUT37), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n578), .B1(new_n581), .B2(new_n575), .ZN(new_n582));
  INV_X1    g381(.A(new_n493), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n583), .B1(new_n533), .B2(new_n534), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n582), .B(KEYINPUT88), .C1(new_n584), .C2(new_n532), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n574), .A2(new_n577), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT87), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT40), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n518), .B1(new_n500), .B2(new_n514), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n530), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n517), .A2(new_n518), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n589), .A2(new_n593), .A3(new_n590), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n587), .B(new_n588), .C1(new_n592), .C2(new_n594), .ZN(new_n595));
  AND4_X1   g394(.A1(new_n533), .A2(new_n595), .A3(new_n559), .A4(new_n557), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n587), .B1(new_n592), .B2(new_n594), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT40), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n492), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n586), .A2(new_n599), .A3(KEYINPUT89), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT89), .B1(new_n586), .B2(new_n599), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n562), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n415), .A2(new_n492), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT90), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT35), .ZN(new_n605));
  INV_X1    g404(.A(new_n561), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n487), .A2(new_n480), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n489), .A2(new_n491), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n610), .A2(new_n604), .A3(new_n406), .A4(new_n414), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT35), .B1(new_n611), .B2(new_n561), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n296), .B1(new_n602), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n283), .A2(KEYINPUT10), .A3(new_n248), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n248), .A2(new_n282), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n239), .A2(new_n280), .A3(new_n281), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n282), .A2(new_n236), .A3(new_n238), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n282), .B1(new_n238), .B2(new_n236), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n616), .B(new_n620), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n615), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n617), .A2(new_n618), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n348), .ZN(new_n636));
  INV_X1    g435(.A(G204gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n628), .A2(new_n640), .A3(new_n632), .A4(new_n633), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(KEYINPUT101), .A3(new_n641), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n271), .A2(new_n247), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n221), .A2(new_n241), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n271), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT18), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n271), .B(new_n247), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n648), .B(KEYINPUT13), .Z(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G113gat), .B(G141gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G197gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT11), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n345), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT12), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n652), .A2(new_n662), .A3(new_n656), .A4(new_n655), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n646), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n614), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n536), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g472(.A1(new_n669), .A2(new_n560), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n266), .B2(new_n268), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n266), .B2(new_n268), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n268), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT42), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(KEYINPUT42), .B2(new_n676), .ZN(G1325gat));
  INV_X1    g478(.A(G15gat), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n416), .B1(new_n415), .B2(new_n297), .ZN(new_n681));
  AOI211_X1 g480(.A(KEYINPUT75), .B(KEYINPUT36), .C1(new_n414), .C2(new_n406), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(KEYINPUT102), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n669), .A2(new_n680), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n415), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n670), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n680), .B2(new_n691), .ZN(G1326gat));
  NOR2_X1   g491(.A1(new_n669), .A2(new_n610), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  AOI21_X1  g494(.A(new_n264), .B1(new_n602), .B2(new_n613), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n295), .A2(new_n646), .A3(new_n667), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(G29gat), .A3(new_n536), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n561), .A2(new_n492), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n681), .B2(new_n682), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n586), .A2(new_n599), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT89), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n586), .A2(new_n599), .A3(KEYINPUT89), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n613), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n263), .B(new_n702), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n711), .B(new_n697), .C1(new_n696), .C2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n671), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT105), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n701), .B1(new_n718), .B2(new_n205), .ZN(G1328gat));
  INV_X1    g518(.A(new_n698), .ZN(new_n720));
  INV_X1    g519(.A(new_n560), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n206), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(KEYINPUT106), .B2(KEYINPUT46), .ZN(new_n723));
  NAND2_X1  g522(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n723), .B(new_n724), .Z(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n715), .B2(new_n560), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1329gat));
  INV_X1    g526(.A(new_n216), .ZN(new_n728));
  INV_X1    g527(.A(new_n683), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n715), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n698), .A2(new_n728), .A3(new_n415), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(new_n732), .A3(KEYINPUT47), .ZN(new_n733));
  INV_X1    g532(.A(new_n688), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n716), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n731), .B1(new_n735), .B2(new_n728), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n733), .B1(new_n736), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g536(.A(new_n263), .B1(new_n709), .B2(new_n710), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n713), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n739), .A2(new_n492), .A3(new_n697), .A4(new_n711), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G50gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT107), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n720), .A2(new_n214), .A3(new_n492), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n740), .A2(new_n745), .A3(G50gat), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n602), .A2(new_n613), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n714), .B1(new_n749), .B2(new_n263), .ZN(new_n750));
  INV_X1    g549(.A(new_n702), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n264), .B(new_n751), .C1(new_n602), .C2(new_n613), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n753), .A2(KEYINPUT108), .A3(new_n492), .A4(new_n697), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n715), .B2(new_n610), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n756), .A3(G50gat), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n743), .B1(new_n757), .B2(new_n744), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n748), .A2(new_n758), .A3(KEYINPUT109), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760));
  INV_X1    g559(.A(new_n756), .ZN(new_n761));
  OAI21_X1  g560(.A(G50gat), .B1(new_n740), .B2(new_n755), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n744), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT48), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n760), .B1(new_n764), .B2(new_n747), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n759), .A2(new_n765), .ZN(G1331gat));
  INV_X1    g565(.A(new_n646), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n602), .B2(new_n613), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n296), .A2(new_n666), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n671), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g572(.A1(new_n770), .A2(new_n560), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  AND2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(G1333gat));
  NAND3_X1  g577(.A1(new_n771), .A2(new_n274), .A3(new_n690), .ZN(new_n779));
  OAI21_X1  g578(.A(G71gat), .B1(new_n770), .B2(new_n688), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g581(.A1(new_n770), .A2(new_n610), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(new_n275), .ZN(G1335gat));
  NOR2_X1   g583(.A1(new_n295), .A2(new_n666), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n696), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(new_n646), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n223), .A3(new_n671), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n753), .A2(new_n646), .A3(new_n785), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n536), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1336gat));
  OR3_X1    g592(.A1(new_n791), .A2(KEYINPUT110), .A3(new_n560), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT110), .B1(new_n791), .B2(new_n560), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(G92gat), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n789), .A2(new_n224), .A3(new_n721), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G92gat), .B1(new_n791), .B2(new_n560), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n801), .B2(new_n797), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n791), .B2(new_n688), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n646), .A2(new_n233), .A3(new_n690), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT111), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n788), .A2(new_n234), .A3(new_n646), .A4(new_n492), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(KEYINPUT112), .ZN(new_n810));
  OAI21_X1  g609(.A(G106gat), .B1(new_n791), .B2(new_n610), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n810), .B(new_n812), .ZN(G1339gat));
  XNOR2_X1  g612(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n626), .A2(new_n627), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n626), .B2(new_n627), .ZN(new_n816));
  INV_X1    g615(.A(new_n615), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT99), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n817), .B1(new_n819), .B2(new_n624), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n629), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n638), .B(new_n815), .C1(new_n816), .C2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT114), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n640), .B1(new_n821), .B2(new_n814), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n820), .A2(new_n629), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n628), .A3(KEYINPUT54), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n825), .A2(new_n827), .A3(new_n828), .A4(KEYINPUT55), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n634), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n823), .A2(new_n822), .B1(new_n831), .B2(new_n640), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n666), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n649), .A2(new_n271), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n648), .B1(new_n834), .B2(new_n647), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n653), .A2(new_n654), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n661), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n665), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n644), .A2(new_n645), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n264), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n830), .A2(new_n832), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n263), .A3(new_n838), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n295), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n769), .A2(new_n767), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n721), .A2(new_n536), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n603), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n667), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(new_n365), .ZN(G1340gat));
  NOR2_X1   g652(.A1(new_n851), .A2(new_n767), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(new_n363), .ZN(G1341gat));
  NOR2_X1   g654(.A1(new_n851), .A2(new_n845), .ZN(new_n856));
  XNOR2_X1  g655(.A(KEYINPUT115), .B(G127gat), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n856), .B(new_n857), .ZN(G1342gat));
  NOR2_X1   g657(.A1(new_n264), .A2(new_n721), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n848), .B1(KEYINPUT116), .B2(new_n859), .ZN(new_n860));
  AOI211_X1 g659(.A(new_n536), .B(new_n860), .C1(KEYINPUT116), .C2(new_n859), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n373), .A3(new_n603), .ZN(new_n862));
  XOR2_X1   g661(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n863));
  XNOR2_X1  g662(.A(new_n862), .B(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n851), .B2(new_n264), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT118), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(G1343gat));
  NAND2_X1  g666(.A1(new_n729), .A2(new_n849), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT119), .B1(new_n840), .B2(new_n264), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871));
  AOI211_X1 g670(.A(new_n871), .B(new_n263), .C1(new_n833), .C2(new_n839), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n842), .A2(new_n263), .A3(new_n838), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n869), .B1(new_n874), .B2(new_n295), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n841), .A2(new_n871), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n840), .A2(KEYINPUT119), .A3(new_n264), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n843), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(KEYINPUT120), .A3(new_n845), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n875), .A2(new_n847), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n492), .A2(KEYINPUT57), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT57), .B1(new_n848), .B2(new_n492), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n868), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n418), .B1(new_n886), .B2(new_n666), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n734), .A2(new_n610), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(new_n850), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n666), .A2(new_n418), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT121), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n890), .A2(KEYINPUT121), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT58), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n886), .B2(new_n666), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n884), .B1(new_n880), .B2(new_n882), .ZN(new_n897));
  NOR4_X1   g696(.A1(new_n897), .A2(KEYINPUT122), .A3(new_n667), .A4(new_n868), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n896), .A2(new_n898), .A3(new_n418), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n893), .A2(KEYINPUT58), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n894), .B1(new_n899), .B2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(new_n495), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n889), .A2(new_n902), .A3(new_n646), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n848), .A2(new_n882), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n868), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n646), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n420), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n767), .B1(new_n885), .B2(new_n905), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(KEYINPUT123), .A3(new_n907), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n904), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT59), .B(new_n902), .C1(new_n886), .C2(new_n646), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n903), .B1(new_n913), .B2(new_n914), .ZN(G1345gat));
  AOI21_X1  g714(.A(G155gat), .B1(new_n889), .B2(new_n295), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n295), .A2(G155gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n886), .B2(new_n917), .ZN(G1346gat));
  INV_X1    g717(.A(G162gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n861), .A2(new_n919), .A3(new_n888), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n897), .A2(new_n264), .A3(new_n868), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n919), .ZN(G1347gat));
  AND2_X1   g721(.A1(new_n848), .A2(new_n603), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n671), .A2(new_n560), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(new_n667), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(new_n345), .ZN(G1348gat));
  OAI21_X1  g726(.A(new_n348), .B1(new_n925), .B2(new_n767), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT124), .Z(new_n929));
  NOR4_X1   g728(.A1(new_n925), .A2(new_n767), .A3(new_n347), .A4(new_n349), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(G1349gat));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n933));
  OAI22_X1  g732(.A1(new_n925), .A2(new_n845), .B1(new_n309), .B2(new_n308), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n923), .A2(new_n295), .A3(new_n924), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n933), .B(new_n934), .C1(new_n935), .C2(new_n324), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n936), .B(new_n937), .Z(G1350gat));
  XNOR2_X1  g737(.A(KEYINPUT61), .B(G190gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n264), .ZN(new_n941));
  MUX2_X1   g740(.A(new_n939), .B(new_n940), .S(new_n941), .Z(G1351gat));
  NAND3_X1  g741(.A1(new_n688), .A2(new_n492), .A3(new_n721), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n848), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n943), .A2(new_n944), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n946), .A2(new_n671), .A3(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(new_n666), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n688), .A2(new_n924), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT127), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(new_n906), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(new_n666), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n950), .B1(new_n954), .B2(new_n949), .ZN(G1352gat));
  NAND3_X1  g754(.A1(new_n948), .A2(new_n637), .A3(new_n646), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n911), .A2(new_n952), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G204gat), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(G1353gat));
  INV_X1    g760(.A(G211gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n948), .A2(new_n962), .A3(new_n295), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n953), .A2(new_n295), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n948), .B2(new_n263), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n263), .A2(G218gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n953), .B2(new_n969), .ZN(G1355gat));
endmodule


