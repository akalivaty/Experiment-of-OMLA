//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n548, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(G2104), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR3_X1   g038(.A1(new_n463), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n469), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n466), .A2(new_n473), .A3(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n468), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT70), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n467), .A2(new_n469), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n461), .A2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  OAI22_X1  g062(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n467), .A2(new_n469), .A3(new_n481), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n481), .B1(new_n467), .B2(new_n469), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n461), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n483), .A2(new_n493), .A3(new_n461), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n488), .B1(G136), .B2(new_n495), .ZN(G162));
  NOR2_X1   g071(.A1(new_n478), .A2(new_n479), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(G126), .A3(G2105), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT72), .B(G114), .ZN(new_n501));
  OAI211_X1 g076(.A(G2104), .B(new_n500), .C1(new_n501), .C2(new_n461), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n461), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n498), .A2(new_n499), .A3(new_n502), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT73), .A3(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n510), .A2(new_n512), .B1(KEYINPUT5), .B2(new_n509), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n518), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT74), .Z(new_n528));
  AND2_X1   g103(.A1(new_n517), .A2(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(G51), .B1(new_n513), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n515), .B1(new_n534), .B2(KEYINPUT75), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n535), .B1(KEYINPUT75), .B2(new_n534), .ZN(new_n536));
  INV_X1    g111(.A(new_n518), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n537), .A2(G90), .B1(G52), .B2(new_n529), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  AOI22_X1  g115(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n515), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n518), .A2(new_n543), .B1(new_n520), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  AOI22_X1  g127(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n553), .A2(new_n554), .A3(new_n515), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n553), .B2(new_n515), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n537), .A2(G91), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n559));
  NAND3_X1  g134(.A1(new_n529), .A2(G53), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n520), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n558), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n557), .A2(new_n565), .ZN(G299));
  NAND2_X1  g141(.A1(new_n528), .A2(new_n531), .ZN(G286));
  OR2_X1    g142(.A1(new_n516), .A2(new_n522), .ZN(G303));
  NAND2_X1  g143(.A1(new_n537), .A2(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n529), .A2(G49), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  AOI22_X1  g147(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n515), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  INV_X1    g150(.A(G48), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n518), .A2(new_n575), .B1(new_n520), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n515), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n518), .A2(new_n582), .B1(new_n520), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n513), .A2(G66), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT78), .Z(new_n590));
  AOI21_X1  g165(.A(new_n515), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n529), .A2(G54), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n594));
  OR3_X1    g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n591), .B2(new_n593), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n518), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n595), .A2(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n587), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n587), .B1(new_n601), .B2(G868), .ZN(G321));
  AOI21_X1  g178(.A(new_n564), .B1(new_n556), .B2(new_n555), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT80), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  MUX2_X1   g181(.A(G286), .B(new_n605), .S(new_n606), .Z(G297));
  MUX2_X1   g182(.A(G286), .B(new_n605), .S(new_n606), .Z(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G860), .ZN(G148));
  OAI21_X1  g185(.A(KEYINPUT81), .B1(new_n546), .B2(G868), .ZN(new_n611));
  INV_X1    g186(.A(new_n601), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G559), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(new_n606), .ZN(new_n614));
  MUX2_X1   g189(.A(new_n611), .B(KEYINPUT81), .S(new_n614), .Z(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n465), .A2(new_n497), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT13), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n495), .A2(G135), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n461), .B1(new_n480), .B2(new_n482), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n623), .A2(new_n624), .B1(new_n626), .B2(G2105), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n622), .A2(G123), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n620), .A2(new_n632), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2451), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n637), .B(new_n638), .Z(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n639), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2454), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n650), .A3(G14), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  AOI21_X1  g232(.A(KEYINPUT18), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT20), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  OR3_X1    g248(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1991), .B(G1996), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1981), .B(G1986), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n677), .B(new_n681), .ZN(G229));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G4), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n601), .B2(new_n683), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G1348), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G26), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G140), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n492), .B2(new_n494), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n461), .A2(G116), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n622), .B2(G128), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(KEYINPUT89), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n493), .B1(new_n483), .B2(new_n461), .ZN(new_n699));
  AOI211_X1 g274(.A(KEYINPUT71), .B(G2105), .C1(new_n480), .C2(new_n482), .ZN(new_n700));
  OAI21_X1  g275(.A(G140), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n701), .A2(new_n702), .A3(new_n696), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n690), .B1(new_n704), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G2067), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n686), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G29), .A2(G35), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G162), .B2(G29), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G2090), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n683), .A2(G20), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT23), .Z(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G299), .B2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G1956), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n683), .A2(G19), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n546), .B2(new_n683), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1341), .ZN(new_n720));
  NOR4_X1   g295(.A1(new_n707), .A2(new_n712), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n683), .A2(G23), .ZN(new_n722));
  INV_X1    g297(.A(G288), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n683), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT33), .B(G1976), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G22), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G166), .B2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT88), .B(G1971), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  NOR2_X1   g305(.A1(G6), .A2(G16), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n578), .B2(G16), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT32), .B(G1981), .Z(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  NOR3_X1   g309(.A1(new_n726), .A2(new_n730), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT34), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n688), .A2(G25), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n495), .A2(G131), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n741));
  INV_X1    g316(.A(G107), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G2105), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n622), .B2(G119), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n739), .B1(new_n746), .B2(new_n688), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT35), .B(G1991), .Z(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n747), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G24), .ZN(new_n751));
  OR3_X1    g326(.A1(new_n751), .A2(KEYINPUT87), .A3(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(KEYINPUT87), .B1(new_n751), .B2(G16), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n752), .B(new_n753), .C1(new_n585), .C2(new_n683), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1986), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n737), .A2(new_n738), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT36), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n683), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n683), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT92), .ZN(new_n761));
  INV_X1    g336(.A(G1966), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n688), .A2(G33), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT91), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT25), .Z(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  INV_X1    g343(.A(G127), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n474), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n767), .B1(G2105), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n495), .A2(G139), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n764), .B1(new_n774), .B2(new_n688), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G2072), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n688), .A2(G32), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n495), .A2(G141), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n465), .A2(G105), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT26), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G129), .B2(new_n622), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n777), .B1(new_n785), .B2(new_n688), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT27), .B(G1996), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n786), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n775), .A2(G2072), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n776), .A2(new_n789), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n683), .A2(G5), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G171), .B2(new_n683), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(G1961), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(G1961), .ZN(new_n796));
  NOR2_X1   g371(.A1(G27), .A2(G29), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G164), .B2(G29), .ZN(new_n798));
  INV_X1    g373(.A(G2078), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n688), .B1(KEYINPUT24), .B2(G34), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(KEYINPUT24), .B2(G34), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n466), .A2(new_n473), .A3(new_n476), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G29), .ZN(new_n804));
  INV_X1    g379(.A(G2084), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT30), .B(G28), .ZN(new_n808));
  OR2_X1    g383(.A1(KEYINPUT31), .A2(G11), .ZN(new_n809));
  NAND2_X1  g384(.A1(KEYINPUT31), .A2(G11), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n808), .A2(new_n688), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n806), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G29), .B2(new_n630), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n795), .A2(new_n796), .A3(new_n800), .A4(new_n813), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n763), .A2(new_n792), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT93), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n763), .A2(KEYINPUT93), .A3(new_n792), .A4(new_n814), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n721), .B(new_n758), .C1(new_n817), .C2(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  NAND2_X1  g395(.A1(new_n601), .A2(G559), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT38), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n529), .A2(G55), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n513), .A2(G93), .A3(new_n517), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n823), .A2(KEYINPUT95), .A3(new_n824), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(new_n515), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n546), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n546), .A3(new_n831), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n822), .B(new_n836), .Z(new_n837));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n838));
  AOI21_X1  g413(.A(G860), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n832), .A2(G860), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  INV_X1    g418(.A(G142), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n492), .B2(new_n494), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n461), .A2(G118), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n622), .B2(G130), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n846), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n618), .ZN(new_n853));
  INV_X1    g428(.A(new_n851), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT97), .B1(new_n845), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n853), .B1(new_n852), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n745), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n852), .A2(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n618), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(new_n746), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n698), .A2(new_n703), .A3(G164), .ZN(new_n864));
  AOI21_X1  g439(.A(G164), .B1(new_n698), .B2(new_n703), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n785), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n692), .A2(new_n697), .A3(KEYINPUT89), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n702), .B1(new_n701), .B2(new_n696), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n506), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n698), .A2(new_n703), .A3(G164), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n784), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n866), .A2(new_n774), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n774), .B1(new_n866), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n863), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n864), .A2(new_n865), .A3(new_n785), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n784), .B1(new_n869), .B2(new_n870), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n773), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n858), .A2(new_n862), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n866), .A2(new_n871), .A3(new_n774), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G162), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n630), .A2(KEYINPUT96), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n621), .B2(new_n629), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n803), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n803), .B1(new_n883), .B2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n882), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(G162), .A3(new_n886), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(G37), .B1(new_n881), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n880), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT98), .A4(new_n879), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n889), .A2(new_n891), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n874), .A4(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n893), .A2(KEYINPUT99), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT99), .B1(new_n893), .B2(new_n898), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  INV_X1    g478(.A(new_n880), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n892), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n898), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n893), .A2(KEYINPUT99), .A3(new_n898), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT40), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n902), .A2(new_n911), .ZN(G395));
  NAND3_X1  g487(.A1(new_n829), .A2(new_n606), .A3(new_n831), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n613), .B(new_n836), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n601), .A2(new_n604), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n557), .A2(new_n565), .A3(new_n916), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n601), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n604), .A2(new_n916), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR3_X1    g496(.A1(new_n915), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(G299), .A2(KEYINPUT100), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n601), .A3(new_n918), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT41), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(new_n921), .B2(new_n917), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n915), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n578), .B(new_n585), .Z(new_n931));
  XNOR2_X1  g506(.A(G166), .B(G288), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(KEYINPUT101), .B2(KEYINPUT42), .ZN(new_n934));
  NAND2_X1  g509(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n934), .B(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n937));
  OR3_X1    g512(.A1(new_n930), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n930), .A2(new_n937), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n922), .A2(KEYINPUT102), .A3(new_n929), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n914), .B1(new_n942), .B2(G868), .ZN(G295));
  AOI21_X1  g518(.A(new_n914), .B1(new_n942), .B2(G868), .ZN(G331));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n921), .A2(new_n917), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n834), .A2(new_n835), .A3(G301), .ZN(new_n947));
  AOI21_X1  g522(.A(G301), .B1(new_n834), .B2(new_n835), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(G286), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n836), .A2(G171), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n834), .A2(new_n835), .A3(G301), .ZN(new_n951));
  AOI21_X1  g526(.A(G168), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n946), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(G286), .B1(new_n947), .B2(new_n948), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(G168), .A3(new_n951), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n928), .A2(new_n926), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n933), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(new_n956), .A3(new_n933), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n945), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n945), .A3(new_n960), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(KEYINPUT44), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n959), .A2(new_n945), .A3(new_n960), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n966), .B2(new_n961), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(G397));
  INV_X1    g543(.A(KEYINPUT61), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n604), .B(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G40), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT104), .B1(new_n803), .B2(new_n973), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n465), .A2(G101), .B1(new_n475), .B2(G137), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n975), .A2(new_n976), .A3(G40), .A4(new_n473), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n506), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n978), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT116), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n506), .A2(new_n980), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n974), .A2(new_n977), .B1(KEYINPUT50), .B2(new_n984), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n716), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n991));
  AOI22_X1  g566(.A1(new_n974), .A2(new_n977), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n981), .A2(KEYINPUT45), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT56), .B(G2072), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n972), .B1(new_n990), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G1956), .B1(new_n983), .B2(new_n988), .ZN(new_n997));
  INV_X1    g572(.A(new_n995), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n997), .A2(new_n971), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n969), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1996), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n984), .A2(new_n991), .ZN(new_n1002));
  AND4_X1   g577(.A1(new_n1001), .A2(new_n978), .A3(new_n993), .A4(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n984), .B1(new_n974), .B2(new_n977), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT58), .B(G1341), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT120), .B(new_n546), .C1(new_n1003), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT59), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n546), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(new_n1010), .A3(KEYINPUT59), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n978), .A2(new_n981), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(G2067), .ZN(new_n1016));
  INV_X1    g591(.A(new_n985), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1348), .B1(new_n986), .B2(new_n1017), .ZN(new_n1018));
  NOR4_X1   g593(.A1(new_n1016), .A2(new_n1018), .A3(new_n612), .A4(KEYINPUT60), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n612), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n1020), .B2(new_n601), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1019), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n990), .A2(new_n972), .A3(new_n995), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n971), .B1(new_n997), .B2(new_n998), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(KEYINPUT61), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1000), .A2(new_n1014), .A3(new_n1025), .A4(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1021), .A2(KEYINPUT119), .A3(new_n601), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1020), .B2(new_n612), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1027), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1026), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n978), .A2(new_n993), .A3(new_n799), .A4(new_n1002), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(KEYINPUT123), .A3(new_n1037), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n986), .A2(new_n1017), .ZN(new_n1042));
  INV_X1    g617(.A(G1961), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1040), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(G301), .B(KEYINPUT54), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n975), .A2(KEYINPUT124), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(G40), .A3(new_n473), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1002), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(KEYINPUT125), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n993), .A2(KEYINPUT53), .A3(new_n799), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT125), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1046), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n991), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n981), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT45), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n984), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n978), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1040), .A2(new_n1041), .A3(new_n1044), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1045), .A2(new_n1055), .B1(new_n1063), .B2(new_n1046), .ZN(new_n1064));
  INV_X1    g639(.A(G1981), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT113), .B1(new_n578), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(G1981), .C1(new_n574), .C2(new_n577), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT112), .B(G1981), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n578), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT49), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT109), .B(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1004), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n1080));
  INV_X1    g655(.A(G1976), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G288), .A2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1004), .A2(new_n1082), .A3(new_n1077), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1077), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1082), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1015), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G303), .A2(G8), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT108), .B(G2090), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1042), .A2(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT107), .B(G1971), .Z(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n992), .B2(new_n993), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1093), .B(G8), .C1(new_n1096), .C2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT52), .B1(G288), .B2(new_n1081), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1015), .A2(new_n1087), .A3(new_n1086), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT111), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1083), .A2(new_n1103), .A3(new_n1100), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  AND4_X1   g680(.A1(new_n1079), .A2(new_n1090), .A3(new_n1099), .A4(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n983), .A2(new_n988), .A3(new_n1094), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n978), .A2(new_n993), .A3(new_n1002), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1097), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1077), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1111), .A2(new_n1093), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1064), .A2(new_n1106), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(G286), .A2(new_n1086), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1060), .A2(new_n762), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n986), .A2(new_n805), .A3(new_n1017), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1077), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1114), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G8), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(new_n1114), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT121), .B(KEYINPUT51), .Z(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1117), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1113), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1035), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1110), .B1(new_n1042), .B2(new_n1095), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G8), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1093), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1136), .B2(new_n1135), .ZN(new_n1138));
  AOI211_X1 g713(.A(G286), .B(new_n1077), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1139));
  AND4_X1   g714(.A1(new_n1079), .A2(new_n1090), .A3(new_n1139), .A4(new_n1105), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1133), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1079), .A2(new_n1090), .A3(new_n1105), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1133), .B(new_n1139), .C1(new_n1111), .C2(new_n1093), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1099), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1078), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1079), .A2(new_n1081), .A3(new_n723), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1070), .B(KEYINPUT115), .Z(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1141), .A2(new_n1144), .A3(new_n1148), .ZN(new_n1149));
  AND4_X1   g724(.A1(G171), .A2(new_n1106), .A3(new_n1112), .A4(new_n1063), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1130), .A2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1120), .A2(new_n1123), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT62), .B1(new_n1153), .B2(new_n1117), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1132), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n784), .B(G1996), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT105), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n704), .A2(G2067), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n704), .A2(G2067), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1161), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1163), .A2(KEYINPUT105), .A3(new_n1159), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1157), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1002), .B1(new_n977), .B2(new_n974), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  OR3_X1    g742(.A1(new_n1165), .A2(KEYINPUT106), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT106), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n746), .A2(new_n748), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n745), .A2(new_n749), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1166), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(new_n1169), .A3(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n585), .B(G1986), .Z(new_n1174));
  AOI21_X1  g749(.A(new_n1173), .B1(new_n1166), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1156), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1166), .A2(new_n1001), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT46), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(KEYINPUT126), .B2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(KEYINPUT126), .B(KEYINPUT46), .Z(new_n1180));
  AOI21_X1  g755(.A(new_n1179), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n784), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1181), .B1(new_n1182), .B2(new_n1167), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT47), .ZN(new_n1184));
  OR3_X1    g759(.A1(new_n1167), .A2(G1986), .A3(G290), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT48), .Z(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1173), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1167), .B1(new_n1188), .B2(new_n1163), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1176), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g766(.A1(G401), .A2(new_n458), .A3(G227), .A4(G229), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1193), .B1(new_n966), .B2(new_n961), .ZN(new_n1194));
  AOI21_X1  g768(.A(new_n1194), .B1(new_n909), .B2(new_n910), .ZN(G308));
  OAI221_X1 g769(.A(new_n1193), .B1(new_n966), .B2(new_n961), .C1(new_n899), .C2(new_n900), .ZN(G225));
endmodule


