//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT22), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT77), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT24), .B(G110), .Z(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n194), .A2(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT71), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT71), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n192), .B1(new_n200), .B2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n195), .A2(new_n197), .A3(new_n193), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT72), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT72), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n211), .A2(new_n193), .A3(KEYINPUT23), .A4(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G110), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n208), .A2(new_n213), .A3(new_n202), .A4(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT75), .B1(new_n205), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT75), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT71), .B1(new_n201), .B2(G128), .ZN(new_n219));
  INV_X1    g033(.A(new_n199), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT67), .B(G119), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(new_n193), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n219), .B1(KEYINPUT71), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n218), .B(new_n215), .C1(new_n223), .C2(new_n192), .ZN(new_n224));
  INV_X1    g038(.A(G140), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G125), .ZN(new_n226));
  INV_X1    g040(.A(G125), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G140), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT16), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT73), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n226), .A2(KEYINPUT16), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT73), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n228), .A3(new_n232), .A4(KEYINPUT16), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n230), .A2(G146), .A3(new_n231), .A4(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT65), .A2(G146), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT65), .A2(G146), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n226), .A2(new_n228), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n217), .A2(new_n224), .A3(new_n234), .A4(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n242));
  INV_X1    g056(.A(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT74), .A3(new_n234), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n223), .A2(new_n192), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT74), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n247), .A3(new_n243), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n208), .A2(new_n213), .A3(new_n202), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G110), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n245), .A2(new_n246), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n241), .A2(KEYINPUT76), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT76), .B1(new_n241), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n191), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G902), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n241), .A2(new_n251), .A3(new_n190), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n254), .A2(KEYINPUT25), .A3(new_n255), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(G217), .ZN(new_n262));
  INV_X1    g076(.A(G234), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G902), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n254), .A2(new_n256), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n265), .A2(G902), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G472), .A2(G902), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT0), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(new_n193), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT65), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n243), .ZN(new_n278));
  INV_X1    g092(.A(G143), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT65), .A2(G146), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n243), .A2(G143), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n275), .B(new_n276), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(G143), .B1(new_n235), .B2(new_n236), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(G146), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n275), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT66), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT11), .ZN(new_n289));
  INV_X1    g103(.A(G134), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n289), .B1(new_n290), .B2(G137), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(G137), .ZN(new_n292));
  INV_X1    g106(.A(G137), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT11), .A3(G134), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G131), .ZN(new_n296));
  INV_X1    g110(.A(G131), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n291), .A2(new_n294), .A3(new_n297), .A4(new_n292), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n281), .A2(new_n282), .ZN(new_n300));
  INV_X1    g114(.A(new_n275), .ZN(new_n301));
  INV_X1    g115(.A(new_n276), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n286), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n288), .A2(new_n299), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n284), .A2(new_n307), .A3(G128), .A4(new_n285), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n193), .B1(new_n284), .B2(KEYINPUT1), .ZN(new_n309));
  INV_X1    g123(.A(new_n282), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(new_n237), .B2(new_n279), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n308), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n292), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n290), .A2(G137), .ZN(new_n314));
  OAI21_X1  g128(.A(G131), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n298), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n306), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n299), .A2(new_n303), .A3(new_n286), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n316), .A2(KEYINPUT30), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n201), .A2(G116), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT2), .B(G113), .Z(new_n324));
  OAI211_X1 g138(.A(new_n323), .B(new_n324), .C1(G116), .C2(new_n194), .ZN(new_n325));
  INV_X1    g139(.A(new_n324), .ZN(new_n326));
  INV_X1    g140(.A(G116), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n221), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n194), .A2(G116), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n319), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G101), .ZN(new_n333));
  INV_X1    g147(.A(G237), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT68), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G237), .ZN(new_n337));
  AOI21_X1  g151(.A(G953), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G210), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT27), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n341), .A3(G210), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT26), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n343), .A2(KEYINPUT26), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n333), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n346), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(G101), .A3(new_n344), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT31), .ZN(new_n351));
  INV_X1    g165(.A(new_n331), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n316), .A2(new_n352), .A3(new_n320), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n332), .A2(new_n350), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(KEYINPUT28), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n316), .A2(new_n352), .A3(new_n356), .A4(new_n320), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n317), .A2(new_n331), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n347), .A2(new_n349), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n353), .ZN(new_n364));
  INV_X1    g178(.A(new_n318), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n306), .B2(new_n316), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(new_n321), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n367), .B2(new_n331), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n351), .B1(new_n368), .B2(new_n350), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT32), .B(new_n273), .C1(new_n363), .C2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n332), .A2(new_n353), .A3(new_n350), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT31), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n354), .A3(new_n362), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT32), .B1(new_n374), .B2(new_n273), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n366), .A2(new_n352), .A3(new_n321), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n361), .B1(new_n377), .B2(new_n364), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n350), .A2(new_n359), .A3(new_n358), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n361), .A2(new_n379), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n316), .A2(new_n320), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n331), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n355), .B2(new_n357), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G472), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT69), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT69), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n391), .A3(G472), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n272), .B1(new_n376), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT78), .A3(G104), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT3), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(G104), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n400), .A2(new_n395), .A3(KEYINPUT78), .A4(G104), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G101), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n397), .A2(new_n399), .A3(new_n333), .A4(new_n401), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(KEYINPUT4), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT79), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n403), .A2(KEYINPUT4), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n403), .A2(new_n408), .A3(KEYINPUT4), .A4(new_n404), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n406), .A2(new_n331), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n323), .B(KEYINPUT5), .C1(G116), .C2(new_n194), .ZN(new_n411));
  OR3_X1    g225(.A1(new_n221), .A2(KEYINPUT5), .A3(new_n327), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(G113), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G104), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G107), .ZN(new_n415));
  OAI21_X1  g229(.A(G101), .B1(new_n398), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n404), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n413), .A2(new_n325), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(G110), .B(G122), .Z(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n420), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n410), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n283), .A2(new_n287), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G125), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n312), .A2(new_n227), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n187), .A2(G224), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n419), .A2(new_n431), .A3(new_n420), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n424), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(KEYINPUT7), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n426), .B2(new_n427), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT83), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n426), .A2(new_n427), .A3(new_n434), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n413), .A2(new_n325), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n404), .A2(new_n416), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n418), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n420), .B(KEYINPUT8), .Z(new_n445));
  AOI22_X1  g259(.A1(new_n444), .A2(new_n445), .B1(new_n439), .B2(new_n438), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n437), .A2(new_n440), .A3(new_n446), .A4(new_n423), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n433), .A2(new_n255), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n433), .A2(new_n447), .A3(new_n255), .A4(new_n449), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n453), .A2(new_n452), .ZN(new_n455));
  INV_X1    g269(.A(G469), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n406), .A2(new_n425), .A3(new_n407), .A4(new_n409), .ZN(new_n457));
  INV_X1    g271(.A(new_n299), .ZN(new_n458));
  INV_X1    g272(.A(new_n308), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT1), .B1(new_n279), .B2(G146), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n193), .B1(new_n460), .B2(KEYINPUT80), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n282), .A2(new_n462), .A3(KEYINPUT1), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n461), .A2(new_n463), .B1(new_n284), .B2(new_n285), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n417), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT10), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n312), .A2(new_n417), .A3(KEYINPUT10), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n457), .A2(new_n458), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G140), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n187), .A2(G227), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n442), .B(new_n308), .C1(new_n311), .C2(new_n309), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n458), .B1(new_n465), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n457), .A2(new_n467), .A3(new_n468), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n299), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n472), .B1(new_n480), .B2(new_n469), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n456), .B(new_n255), .C1(new_n478), .C2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n456), .A2(new_n255), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n472), .ZN(new_n485));
  INV_X1    g299(.A(new_n469), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n477), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n480), .A2(new_n469), .A3(new_n472), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(G469), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n482), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n454), .A2(new_n455), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n245), .A2(new_n248), .ZN(new_n492));
  AOI21_X1  g306(.A(G143), .B1(new_n338), .B2(G214), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n338), .A2(G143), .A3(G214), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT17), .A3(G131), .ZN(new_n497));
  INV_X1    g311(.A(new_n495), .ZN(new_n498));
  OAI21_X1  g312(.A(G131), .B1(new_n498), .B2(new_n493), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(new_n297), .A3(new_n495), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n492), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n414), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT18), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n506), .A2(new_n297), .A3(KEYINPUT85), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n496), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n496), .A2(new_n507), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n240), .B1(new_n243), .B2(new_n239), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n503), .A2(new_n505), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n503), .A2(new_n511), .A3(KEYINPUT86), .A4(new_n505), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n499), .A2(new_n500), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n239), .B(KEYINPUT19), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n238), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n234), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n505), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G475), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n255), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n503), .A2(new_n511), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n522), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n516), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n255), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G475), .ZN(new_n533));
  INV_X1    g347(.A(G478), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT13), .B1(new_n193), .B2(G143), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n290), .ZN(new_n538));
  XNOR2_X1  g352(.A(G128), .B(G143), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G122), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G116), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT87), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n327), .A2(G122), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(new_n395), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n543), .A2(new_n395), .A3(new_n544), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n540), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n543), .B1(KEYINPUT14), .B2(new_n544), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n544), .A2(KEYINPUT14), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT88), .ZN(new_n551));
  OAI21_X1  g365(.A(G107), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n547), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n539), .B(new_n290), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT9), .B(G234), .Z(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(new_n187), .A3(new_n262), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n558), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n548), .A2(new_n555), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n536), .B1(new_n562), .B2(new_n255), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G952), .ZN(new_n565));
  AOI211_X1 g379(.A(G953), .B(new_n565), .C1(G234), .C2(G237), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT21), .B(G898), .Z(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT90), .ZN(new_n568));
  OAI211_X1 g382(.A(G902), .B(G953), .C1(new_n263), .C2(new_n334), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT89), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n562), .A2(new_n255), .A3(new_n536), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(G475), .B1(new_n516), .B2(new_n523), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(KEYINPUT20), .A3(new_n255), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n528), .A2(new_n533), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n557), .A2(new_n255), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n579), .A2(G221), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G214), .B1(G237), .B2(G902), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n582), .B(KEYINPUT81), .Z(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n491), .A2(new_n578), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n394), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  NAND3_X1  g402(.A1(new_n528), .A2(new_n533), .A3(new_n577), .ZN(new_n589));
  AOI21_X1  g403(.A(G478), .B1(new_n562), .B2(new_n255), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n590), .A2(KEYINPUT91), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(KEYINPUT91), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n562), .B(KEYINPUT33), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(G478), .A3(new_n255), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n571), .A2(new_n583), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n451), .B2(new_n453), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n589), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT92), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n589), .A2(KEYINPUT92), .A3(new_n596), .A4(new_n599), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n264), .B1(new_n259), .B2(new_n260), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n270), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n490), .A2(new_n581), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n374), .A2(new_n255), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n608), .A2(G472), .B1(new_n273), .B2(new_n374), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  AOI21_X1  g427(.A(KEYINPUT20), .B1(new_n576), .B2(new_n255), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n514), .A2(new_n515), .B1(new_n522), .B2(new_n521), .ZN(new_n615));
  NOR4_X1   g429(.A1(new_n615), .A2(new_n527), .A3(G475), .A4(G902), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n525), .B1(new_n531), .B2(new_n255), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n564), .A2(new_n573), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n618), .A2(new_n619), .A3(new_n599), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n610), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  NOR2_X1   g437(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT93), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n252), .A2(new_n253), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n268), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n266), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n609), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n586), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(KEYINPUT94), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT37), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n214), .ZN(G12));
  OAI21_X1  g450(.A(new_n273), .B1(new_n363), .B2(new_n369), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT32), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n391), .B1(new_n388), .B2(G472), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  AOI211_X1 g455(.A(KEYINPUT69), .B(new_n641), .C1(new_n381), .C2(new_n387), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n639), .B(new_n370), .C1(new_n640), .C2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n583), .B1(new_n451), .B2(new_n453), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n643), .A2(new_n607), .A3(new_n629), .A4(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n619), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n570), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n566), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n589), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  NOR2_X1   g466(.A1(new_n350), .A2(new_n364), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n255), .B1(new_n654), .B2(new_n385), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n368), .A2(new_n361), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n376), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n490), .A2(new_n581), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n649), .B(KEYINPUT39), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT96), .B(KEYINPUT40), .Z(new_n663));
  OAI211_X1 g477(.A(new_n619), .B(new_n589), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n659), .B(new_n664), .C1(new_n662), .C2(new_n663), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n454), .A2(new_n455), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT95), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n454), .A2(new_n455), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT95), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT38), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n668), .A2(KEYINPUT38), .A3(new_n670), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n665), .A2(new_n584), .A3(new_n630), .A4(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT97), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  INV_X1    g493(.A(new_n649), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n589), .A2(new_n607), .A3(new_n596), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n451), .A2(new_n453), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n584), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n393), .B2(new_n376), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n681), .A2(new_n684), .A3(KEYINPUT98), .A4(new_n629), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT98), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n643), .A2(new_n629), .A3(new_n644), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n589), .A2(new_n607), .A3(new_n596), .A4(new_n680), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT99), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n243), .ZN(G48));
  OAI21_X1  g506(.A(new_n255), .B1(new_n478), .B2(new_n481), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G469), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n694), .A2(new_n482), .A3(new_n581), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n640), .A2(new_n642), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n639), .A2(new_n370), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n606), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n604), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT100), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT100), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n604), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT41), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G113), .ZN(G15));
  NAND2_X1  g520(.A1(new_n699), .A2(new_n620), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NOR4_X1   g522(.A1(new_n614), .A2(new_n616), .A3(new_n617), .A4(new_n574), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n684), .A2(new_n709), .A3(new_n629), .A4(new_n695), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  AOI21_X1  g525(.A(KEYINPUT101), .B1(new_n266), .B2(new_n271), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n605), .A2(new_n713), .A3(new_n270), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n589), .A2(new_n619), .A3(new_n599), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n608), .A2(G472), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n354), .B1(new_n350), .B2(new_n386), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n273), .B1(new_n718), .B2(new_n369), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n715), .A2(new_n695), .A3(new_n716), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NAND3_X1  g536(.A1(new_n589), .A2(new_n596), .A3(new_n680), .ZN(new_n723));
  OR2_X1    g537(.A1(new_n625), .A2(new_n626), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n625), .A2(new_n626), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n269), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n717), .B(new_n719), .C1(new_n726), .C2(new_n605), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n695), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n683), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  INV_X1    g546(.A(new_n723), .ZN(new_n733));
  AND4_X1   g547(.A1(KEYINPUT102), .A2(new_n669), .A3(new_n584), .A4(new_n607), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n583), .B1(new_n454), .B2(new_n455), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT102), .B1(new_n735), .B2(new_n607), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n394), .B(new_n733), .C1(new_n734), .C2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n607), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n735), .A2(KEYINPUT102), .A3(new_n607), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n643), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n745), .A2(new_n712), .A3(new_n714), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(KEYINPUT42), .A3(new_n746), .A4(new_n733), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n739), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  OAI211_X1 g563(.A(new_n394), .B(new_n650), .C1(new_n734), .C2(new_n736), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND2_X1  g565(.A1(new_n618), .A2(new_n596), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n631), .A3(new_n629), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT44), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n735), .B(KEYINPUT105), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT106), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n487), .A2(new_n488), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n487), .A2(KEYINPUT45), .A3(new_n488), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(G469), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n484), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n482), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT103), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  INV_X1    g583(.A(new_n765), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n770), .B2(new_n483), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT104), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT104), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n773), .B(new_n769), .C1(new_n770), .C2(new_n483), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT103), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n766), .A2(new_n775), .A3(new_n482), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n768), .A2(new_n772), .A3(new_n774), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n581), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n661), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n759), .A2(KEYINPUT106), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n760), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n777), .A2(new_n783), .A3(new_n581), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n783), .B1(new_n777), .B2(new_n581), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n785), .A3(new_n643), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n272), .A3(new_n733), .A4(new_n735), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT107), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n225), .ZN(G42));
  AND2_X1   g603(.A1(new_n673), .A2(new_n674), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n694), .A2(new_n482), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT49), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n752), .A2(new_n712), .A3(new_n714), .A4(new_n585), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n790), .A2(new_n659), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n645), .A2(new_n650), .B1(new_n728), .B2(new_n730), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n618), .A2(new_n683), .A3(new_n646), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n629), .A2(new_n649), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n607), .A3(new_n797), .A4(new_n658), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n690), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT112), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n690), .A2(new_n795), .A3(new_n801), .A4(new_n798), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT113), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(new_n800), .B2(new_n802), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n690), .A2(new_n795), .A3(KEYINPUT52), .A4(new_n798), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT111), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n728), .B1(new_n734), .B2(new_n736), .ZN(new_n813));
  INV_X1    g627(.A(new_n740), .ZN(new_n814));
  INV_X1    g628(.A(new_n573), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT108), .B1(new_n815), .B2(new_n563), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT108), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n564), .A2(new_n817), .A3(new_n573), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n393), .B2(new_n376), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n589), .A2(new_n649), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n814), .A2(new_n629), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n750), .A2(new_n813), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n823), .A2(new_n824), .B1(new_n739), .B2(new_n747), .ZN(new_n825));
  AOI211_X1 g639(.A(KEYINPUT100), .B(new_n698), .C1(new_n602), .C2(new_n603), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n702), .B1(new_n604), .B2(new_n699), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n633), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n643), .A2(new_n709), .A3(new_n629), .A4(new_n644), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n829), .A2(new_n695), .B1(new_n394), .B2(new_n586), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n528), .A2(new_n819), .A3(new_n533), .A4(new_n577), .ZN(new_n831));
  INV_X1    g645(.A(new_n596), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n831), .B1(new_n618), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n610), .A2(new_n833), .A3(new_n666), .A4(new_n597), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n830), .A2(new_n707), .A3(new_n721), .A4(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n828), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n750), .A2(new_n813), .A3(new_n822), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT109), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n825), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n812), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  XNOR2_X1  g657(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n803), .A2(new_n804), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n807), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(new_n839), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n842), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n754), .A2(new_n566), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n669), .A2(new_n584), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n729), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n746), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT48), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n565), .A2(G953), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n589), .A2(new_n596), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n851), .A2(new_n606), .A3(new_n566), .A4(new_n659), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n853), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n790), .A2(KEYINPUT117), .A3(new_n583), .A4(new_n695), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n715), .A2(new_n720), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n754), .A2(new_n859), .A3(new_n566), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n673), .A2(new_n583), .A3(new_n674), .A4(new_n695), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n858), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n858), .A2(KEYINPUT50), .A3(new_n860), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n791), .A2(new_n580), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n784), .B2(new_n785), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n566), .A2(new_n758), .A3(new_n859), .A4(new_n754), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n870), .A2(KEYINPUT116), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT116), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n849), .A2(new_n851), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n727), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n856), .A2(new_n589), .A3(new_n596), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n868), .A2(new_n874), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n857), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n860), .A2(new_n730), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n876), .B(new_n878), .C1(new_n866), .C2(new_n867), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n870), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g701(.A(KEYINPUT118), .B(new_n869), .C1(new_n784), .C2(new_n785), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n871), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n889), .A2(KEYINPUT51), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n884), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n878), .B1(new_n866), .B2(new_n867), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n884), .A2(new_n892), .A3(new_n890), .A4(new_n877), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n882), .B(new_n883), .C1(new_n891), .C2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n633), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n701), .B2(new_n703), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n721), .A2(new_n834), .A3(new_n710), .A4(new_n587), .ZN(new_n897));
  INV_X1    g711(.A(new_n707), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n838), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n748), .B1(KEYINPUT109), .B2(new_n837), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT110), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT110), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n825), .A2(new_n836), .A3(new_n903), .A4(new_n838), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n808), .B1(new_n803), .B2(new_n804), .ZN(new_n906));
  AOI211_X1 g720(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n800), .C2(new_n802), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n908), .B2(new_n811), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT114), .B1(new_n909), .B2(KEYINPUT53), .ZN(new_n910));
  OR3_X1    g724(.A1(new_n846), .A2(new_n839), .A3(new_n844), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT114), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n806), .A2(new_n809), .A3(new_n811), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n912), .B(new_n840), .C1(new_n913), .C2(new_n905), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n848), .B(new_n894), .C1(KEYINPUT54), .C2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n794), .B1(new_n916), .B2(new_n917), .ZN(G75));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n842), .A2(new_n847), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(G902), .ZN(new_n921));
  INV_X1    g735(.A(G210), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n424), .A2(new_n432), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(new_n430), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT55), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n923), .A2(new_n926), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n187), .A2(G952), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT120), .Z(new_n930));
  NOR3_X1   g744(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(G51));
  XNOR2_X1  g745(.A(new_n483), .B(KEYINPUT57), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n843), .B1(new_n842), .B2(new_n847), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n848), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n478), .A2(new_n481), .ZN(new_n937));
  OAI211_X1 g751(.A(KEYINPUT121), .B(new_n932), .C1(new_n848), .C2(new_n933), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n921), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n770), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n929), .B1(new_n939), .B2(new_n941), .ZN(G54));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT58), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n525), .ZN(new_n945));
  NAND3_X1  g759(.A1(KEYINPUT122), .A2(KEYINPUT58), .A3(G475), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n940), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n947), .A2(new_n615), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n615), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n929), .ZN(G60));
  INV_X1    g764(.A(new_n930), .ZN(new_n951));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT59), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n848), .B2(new_n933), .ZN(new_n954));
  INV_X1    g768(.A(new_n594), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n915), .A2(KEYINPUT54), .ZN(new_n957));
  INV_X1    g771(.A(new_n848), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n953), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n956), .B1(new_n960), .B2(new_n955), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n920), .A2(new_n627), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n966), .A3(new_n951), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n920), .A2(new_n964), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n267), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n951), .A3(new_n965), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n968), .B(new_n971), .ZN(G66));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n836), .B(KEYINPUT124), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n187), .ZN(new_n975));
  INV_X1    g789(.A(G224), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n568), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n973), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n973), .B2(new_n977), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n924), .B1(G898), .B2(new_n187), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n979), .B(new_n980), .Z(G69));
  XOR2_X1   g795(.A(new_n367), .B(new_n518), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(G900), .B1(new_n983), .B2(G227), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n187), .B(new_n984), .C1(G227), .C2(new_n983), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n690), .A2(new_n795), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n987), .A2(new_n748), .A3(new_n750), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n779), .A2(new_n746), .A3(new_n796), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n781), .A2(new_n787), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(G953), .B1(new_n991), .B2(new_n983), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n678), .A2(new_n987), .ZN(new_n993));
  XNOR2_X1  g807(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n678), .A2(new_n987), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n995), .A2(new_n781), .A3(new_n787), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n850), .A2(new_n662), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n999), .A2(new_n394), .A3(new_n833), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n982), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n985), .B1(new_n992), .B2(new_n1001), .ZN(G72));
  NOR3_X1   g816(.A1(new_n998), .A2(new_n974), .A3(new_n1000), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n656), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n990), .B2(new_n974), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n654), .A2(new_n377), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n929), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1009), .A2(new_n656), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n915), .A2(new_n1012), .A3(new_n1005), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n915), .A2(KEYINPUT127), .A3(new_n1012), .A4(new_n1005), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1011), .B1(new_n1015), .B2(new_n1016), .ZN(G57));
endmodule


