//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n193), .A3(new_n197), .A4(new_n191), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT65), .B1(new_n205), .B2(G146), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(G146), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n201), .B(new_n204), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n203), .A2(G143), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n200), .B(new_n209), .C1(new_n207), .C2(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n194), .A2(KEYINPUT66), .A3(G131), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n199), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(G143), .B2(new_n203), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n216), .A2(new_n217), .B1(new_n207), .B2(new_n210), .ZN(new_n218));
  OAI211_X1 g032(.A(G128), .B(new_n204), .C1(new_n206), .C2(new_n207), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(KEYINPUT1), .ZN(new_n220));
  INV_X1    g034(.A(new_n191), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n189), .A2(G137), .ZN(new_n222));
  OAI21_X1  g036(.A(G131), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(new_n198), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT64), .B1(new_n214), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT70), .B1(new_n214), .B2(new_n224), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT30), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n187), .A2(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n214), .A2(new_n224), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT70), .A3(KEYINPUT30), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT68), .A2(G119), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT68), .A2(G119), .ZN(new_n234));
  OAI21_X1  g048(.A(G116), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT2), .A2(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT67), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT2), .A3(G113), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT2), .A2(G113), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n235), .A2(new_n243), .A3(new_n244), .A4(new_n237), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(KEYINPUT69), .A3(new_n247), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n228), .A2(new_n232), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G101), .ZN(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n254), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n250), .A2(new_n214), .A3(new_n251), .A4(new_n224), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n253), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT31), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n252), .A2(new_n229), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(new_n260), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n252), .A2(new_n229), .A3(KEYINPUT73), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(KEYINPUT28), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n229), .A2(KEYINPUT74), .ZN(new_n268));
  INV_X1    g082(.A(new_n251), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT69), .B1(new_n246), .B2(new_n247), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT74), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n214), .A2(new_n272), .A3(new_n224), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n268), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n259), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n280));
  NAND4_X1  g094(.A1(new_n253), .A2(new_n259), .A3(new_n260), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n262), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n282), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n267), .A2(new_n259), .A3(new_n276), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n259), .B1(new_n253), .B2(new_n260), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT29), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n263), .A2(new_n260), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n276), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n259), .A2(KEYINPUT29), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT75), .B(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G472), .B1(new_n290), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n286), .A2(new_n287), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G128), .B1(new_n233), .B2(new_n234), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT23), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n304));
  INV_X1    g118(.A(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT68), .A2(G119), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n217), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT76), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n306), .A2(new_n310), .A3(new_n217), .A4(new_n307), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n303), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n305), .A2(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(KEYINPUT77), .A3(new_n314), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(G110), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(G125), .ZN(new_n323));
  INV_X1    g137(.A(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n326), .B2(new_n320), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n203), .ZN(new_n328));
  OAI211_X1 g142(.A(G146), .B(new_n322), .C1(new_n326), .C2(new_n320), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n306), .A2(new_n307), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n313), .B1(new_n332), .B2(G128), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n319), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n315), .A2(G110), .B1(new_n333), .B2(new_n334), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G125), .B(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT16), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n341), .A2(KEYINPUT78), .A3(G146), .A4(new_n322), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n337), .B(new_n343), .C1(G146), .C2(new_n326), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT79), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n336), .A2(new_n347), .A3(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(G953), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(G221), .A3(G234), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT22), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(new_n192), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n352), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n345), .A2(KEYINPUT79), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n298), .B2(G234), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G902), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(KEYINPUT81), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n348), .A2(new_n352), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n347), .B1(new_n336), .B2(new_n344), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n355), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n298), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT25), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n297), .B1(new_n353), .B2(new_n355), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(KEYINPUT80), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n371), .A3(new_n358), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n301), .A2(new_n361), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT9), .B(G234), .Z(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n199), .A2(new_n213), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT12), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(new_n379), .B2(G107), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G104), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(G107), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n380), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n382), .A2(G104), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n379), .A2(G107), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n216), .A2(KEYINPUT82), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G128), .B1(new_n216), .B2(KEYINPUT82), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n206), .A2(new_n207), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(new_n215), .A3(G128), .A4(new_n204), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n390), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n390), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(new_n220), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n377), .B(new_n378), .C1(new_n398), .C2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n380), .A2(new_n383), .A3(new_n385), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G101), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT4), .A3(new_n386), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n405), .A3(G101), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n212), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n220), .A3(KEYINPUT10), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n407), .B(new_n408), .C1(new_n398), .C2(KEYINPUT10), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n401), .B1(new_n409), .B2(new_n377), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n377), .B1(new_n398), .B2(new_n400), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(KEYINPUT12), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT83), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  INV_X1    g228(.A(G227), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G953), .ZN(new_n416));
  XOR2_X1   g230(.A(new_n414), .B(new_n416), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n407), .A2(new_n408), .ZN(new_n419));
  INV_X1    g233(.A(new_n377), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n419), .B(new_n420), .C1(KEYINPUT10), .C2(new_n398), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n411), .A2(KEYINPUT12), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .A4(new_n401), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n413), .A2(new_n418), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n409), .A2(new_n377), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n426), .A3(new_n417), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n427), .A3(G469), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n410), .A2(new_n412), .A3(new_n418), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n417), .B1(new_n421), .B2(new_n426), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n430), .B(new_n298), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G902), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n376), .B1(new_n429), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT96), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT15), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n439), .A2(KEYINPUT15), .ZN(new_n442));
  OAI21_X1  g256(.A(G478), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n205), .A2(G128), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n217), .A2(G143), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n446), .A2(new_n189), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n447), .A2(KEYINPUT92), .ZN(new_n448));
  INV_X1    g262(.A(new_n444), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n449), .A2(KEYINPUT13), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(KEYINPUT13), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(new_n445), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G134), .ZN(new_n453));
  XNOR2_X1  g267(.A(G116), .B(G122), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(new_n382), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n447), .A2(KEYINPUT92), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n448), .A2(new_n453), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n382), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT94), .B1(new_n236), .B2(G122), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n236), .A2(G122), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n460), .B1(KEYINPUT14), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G122), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n463), .B2(G116), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT93), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT93), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT14), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(new_n236), .A3(KEYINPUT94), .A4(G122), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n462), .A2(new_n465), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n459), .B1(new_n470), .B2(G107), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n446), .B(new_n189), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n471), .A2(KEYINPUT95), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT95), .B1(new_n471), .B2(new_n472), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n457), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n375), .A2(new_n357), .A3(G953), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n457), .B(new_n476), .C1(new_n473), .C2(new_n474), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n443), .B1(new_n480), .B2(new_n298), .ZN(new_n481));
  INV_X1    g295(.A(new_n443), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n297), .B(new_n482), .C1(new_n478), .C2(new_n479), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n326), .A2(KEYINPUT19), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT19), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n340), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n485), .B1(new_n489), .B2(G146), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(G143), .B1(new_n255), .B2(G214), .ZN(new_n493));
  OAI21_X1  g307(.A(G131), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G237), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n349), .A3(G214), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n205), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n197), .A3(new_n491), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT90), .A4(new_n203), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n343), .A2(new_n490), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n340), .B(new_n203), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n497), .B(new_n491), .C1(new_n503), .C2(new_n197), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n502), .B(new_n504), .C1(new_n503), .C2(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(new_n379), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n494), .A2(new_n511), .A3(new_n498), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n494), .A2(new_n511), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n494), .A2(KEYINPUT91), .A3(new_n511), .A4(new_n498), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n514), .A2(new_n330), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n508), .A3(new_n505), .ZN(new_n518));
  AOI21_X1  g332(.A(G475), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n519), .A2(KEYINPUT20), .A3(new_n434), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT20), .B1(new_n519), .B2(new_n434), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(G234), .A2(G237), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(G952), .A3(new_n349), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n297), .A2(G953), .A3(new_n523), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT21), .B(G898), .Z(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n518), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n508), .B1(new_n517), .B2(new_n505), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n434), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G475), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n484), .A2(new_n522), .A3(new_n531), .A4(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G214), .B1(G237), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n438), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT84), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n212), .B2(new_n324), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n208), .A2(new_n211), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(KEYINPUT84), .A3(G125), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(KEYINPUT85), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT85), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT84), .B1(new_n542), .B2(G125), .ZN(new_n546));
  AOI211_X1 g360(.A(new_n540), .B(new_n324), .C1(new_n208), .C2(new_n211), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT86), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n220), .B2(G125), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n397), .A2(KEYINPUT86), .A3(new_n324), .A4(new_n218), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n544), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G224), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(G953), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n553), .A2(KEYINPUT88), .A3(KEYINPUT7), .A4(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT88), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n544), .A2(new_n548), .A3(new_n556), .A4(new_n552), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n404), .A2(new_n406), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n269), .B2(new_n270), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n235), .A2(KEYINPUT5), .A3(new_n237), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n565), .B(G113), .C1(KEYINPUT5), .C2(new_n235), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n247), .A3(new_n399), .ZN(new_n567));
  XOR2_X1   g381(.A(G110), .B(G122), .Z(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n564), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n552), .A2(new_n541), .A3(new_n543), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n560), .A2(KEYINPUT87), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n560), .A2(KEYINPUT87), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n556), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n566), .A2(new_n247), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n390), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n567), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n568), .B(KEYINPUT8), .Z(new_n578));
  AOI22_X1  g392(.A1(new_n571), .A2(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n557), .A2(new_n561), .A3(new_n570), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n544), .A2(new_n548), .A3(new_n552), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n555), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n559), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n562), .B1(new_n250), .B2(new_n251), .ZN(new_n584));
  INV_X1    g398(.A(new_n567), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n568), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n570), .A3(KEYINPUT6), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT6), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n588), .B(new_n568), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n583), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(new_n590), .A3(new_n434), .ZN(new_n591));
  OAI21_X1  g405(.A(G210), .B1(G237), .B2(G902), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT89), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n580), .A2(new_n590), .A3(new_n434), .A4(new_n592), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(new_n595), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n539), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n373), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT97), .B(G101), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G3));
  NAND2_X1  g417(.A1(new_n594), .A2(new_n596), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT98), .B1(new_n604), .B2(new_n537), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n606));
  AOI211_X1 g420(.A(new_n606), .B(new_n538), .C1(new_n594), .C2(new_n596), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n480), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n478), .A2(KEYINPUT33), .A3(new_n479), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n298), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G478), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n519), .A2(new_n434), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT20), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n519), .A2(KEYINPUT20), .A3(new_n434), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n535), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n480), .A2(new_n298), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(G478), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n612), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NOR4_X1   g435(.A1(new_n605), .A2(new_n607), .A3(new_n530), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n282), .A2(new_n298), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n623), .A2(G472), .B1(new_n283), .B2(new_n282), .ZN(new_n624));
  INV_X1    g438(.A(new_n438), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n624), .A2(new_n372), .A3(new_n625), .A4(new_n361), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NOR3_X1   g444(.A1(new_n605), .A2(new_n607), .A3(new_n530), .ZN(new_n631));
  INV_X1    g445(.A(new_n484), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n615), .A2(new_n535), .A3(new_n616), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n627), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NOR2_X1   g452(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n345), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n360), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n372), .A2(new_n643), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n599), .A2(new_n644), .A3(new_n539), .A4(new_n624), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT100), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n525), .B1(new_n527), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n632), .A2(new_n633), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n644), .A2(new_n625), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n604), .A2(new_n537), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n606), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n604), .A2(KEYINPUT98), .A3(new_n537), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n301), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n649), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n438), .B(new_n653), .C1(new_n372), .C2(new_n643), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n605), .A2(new_n607), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n661), .A2(KEYINPUT101), .A3(new_n301), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT102), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n217), .ZN(G30));
  NAND2_X1  g480(.A1(new_n597), .A2(new_n598), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT38), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n651), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n625), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n674));
  INV_X1    g488(.A(new_n644), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n253), .A2(new_n260), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n259), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n434), .B1(new_n291), .B2(new_n259), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n286), .A2(new_n287), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n633), .A2(new_n484), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n683), .B1(new_n673), .B2(KEYINPUT40), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n671), .A2(new_n537), .A3(new_n674), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  NAND2_X1  g501(.A1(new_n644), .A2(new_n625), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n659), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n621), .A2(new_n651), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  INV_X1    g506(.A(new_n432), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n421), .A2(new_n417), .A3(new_n423), .A4(new_n401), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI211_X1 g509(.A(KEYINPUT104), .B(new_n430), .C1(new_n695), .C2(new_n298), .ZN(new_n696));
  INV_X1    g510(.A(new_n376), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n430), .A2(KEYINPUT104), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n297), .B(new_n698), .C1(new_n693), .C2(new_n694), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  AND4_X1   g514(.A1(new_n361), .A2(new_n301), .A3(new_n372), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n622), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT105), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT41), .B(G113), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND3_X1  g519(.A1(new_n701), .A2(new_n631), .A3(new_n635), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  INV_X1    g521(.A(new_n700), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n708), .A2(new_n605), .A3(new_n607), .ZN(new_n709));
  INV_X1    g523(.A(new_n536), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n301), .A3(new_n710), .A4(new_n644), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT106), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  AND3_X1   g527(.A1(new_n662), .A2(new_n531), .A3(new_n683), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n293), .A2(new_n278), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n262), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n262), .A2(new_n715), .A3(KEYINPUT108), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n281), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n283), .B(KEYINPUT107), .Z(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n623), .A2(G472), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n372), .A2(new_n361), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n724), .A2(new_n725), .A3(new_n708), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n714), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n463), .ZN(G24));
  AOI22_X1  g542(.A1(new_n720), .A2(new_n721), .B1(G472), .B2(new_n623), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n729), .A2(new_n644), .A3(new_n690), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n709), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  NAND2_X1  g546(.A1(new_n286), .A2(KEYINPUT110), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n284), .A2(new_n734), .A3(new_n285), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n287), .A3(new_n300), .A4(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n437), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n425), .A2(KEYINPUT109), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n413), .A2(new_n424), .A3(new_n739), .A4(new_n418), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n738), .A2(G469), .A3(new_n427), .A4(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n697), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n667), .A2(new_n742), .A3(new_n537), .ZN(new_n743));
  INV_X1    g557(.A(new_n725), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n736), .A2(new_n743), .A3(new_n744), .A4(new_n690), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT42), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n667), .A2(new_n742), .A3(new_n537), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n373), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n690), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n654), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT111), .B(G134), .Z(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G36));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n619), .B1(G478), .B2(new_n611), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n633), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT113), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n762), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n757), .A2(KEYINPUT43), .A3(new_n633), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n624), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n644), .B1(new_n768), .B2(new_n769), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n756), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n772), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT44), .A3(new_n770), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n667), .A2(new_n537), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n738), .A2(KEYINPUT45), .A3(new_n427), .A4(new_n740), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n425), .A2(new_n427), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(G469), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n778), .B1(new_n784), .B2(new_n435), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n436), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n433), .A3(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n787), .A2(new_n376), .A3(new_n672), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n773), .A2(new_n775), .A3(new_n777), .A4(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT116), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n192), .ZN(G39));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n787), .A2(new_n792), .A3(new_n376), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n792), .B1(new_n787), .B2(new_n376), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n793), .A2(new_n794), .A3(new_n776), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n744), .A2(new_n301), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n690), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  INV_X1    g612(.A(new_n671), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n725), .A2(new_n681), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n696), .A2(new_n699), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n758), .B1(new_n802), .B2(KEYINPUT49), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(KEYINPUT49), .B2(new_n802), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n804), .A2(new_n538), .A3(new_n697), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n799), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n776), .A2(new_n708), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n800), .A3(new_n525), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n621), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n524), .B1(new_n764), .B2(new_n767), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n538), .A3(new_n726), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n671), .A2(new_n811), .A3(KEYINPUT50), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n808), .A2(new_n617), .A3(new_n757), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI22_X1  g628(.A1(new_n793), .A2(new_n794), .B1(new_n376), .B2(new_n802), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n724), .A2(new_n725), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(new_n816), .A3(new_n777), .A4(new_n810), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n810), .A2(new_n807), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n644), .A3(new_n729), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT50), .B1(new_n671), .B2(new_n811), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n814), .A2(new_n817), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT120), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT51), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(KEYINPUT120), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n736), .A2(new_n744), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n818), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT48), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n810), .A2(new_n709), .A3(new_n816), .ZN(new_n829));
  AND4_X1   g643(.A1(G952), .A2(new_n828), .A3(new_n349), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(new_n825), .A3(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n689), .A2(new_n690), .B1(new_n730), .B2(new_n709), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n662), .A2(new_n683), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n742), .A2(new_n652), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n675), .A3(new_n681), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n664), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n832), .A2(new_n664), .A3(KEYINPUT52), .A4(new_n835), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n714), .A2(new_n726), .B1(new_n701), .B2(new_n622), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n634), .A2(new_n621), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n530), .A2(new_n538), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n598), .A3(new_n597), .A4(new_n843), .ZN(new_n844));
  OAI22_X1  g658(.A1(new_n373), .A2(new_n600), .B1(new_n626), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n645), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n841), .A2(new_n846), .A3(new_n706), .A4(new_n711), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n730), .B2(new_n743), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n729), .A2(new_n644), .A3(new_n690), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n850), .A2(KEYINPUT117), .A3(new_n747), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n632), .A2(new_n617), .A3(new_n651), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n777), .A2(new_n301), .A3(new_n852), .ZN(new_n853));
  OAI22_X1  g667(.A1(new_n849), .A2(new_n851), .B1(new_n853), .B2(new_n688), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n746), .A2(new_n750), .A3(new_n753), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n847), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n840), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n840), .A2(new_n856), .A3(KEYINPUT53), .ZN(new_n860));
  XOR2_X1   g674(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n863), .A2(KEYINPUT119), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n840), .A2(new_n856), .A3(KEYINPUT53), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n840), .B2(new_n856), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n863), .B(KEYINPUT119), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n809), .B(new_n831), .C1(new_n864), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(G952), .A2(G953), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n806), .B1(new_n870), .B2(new_n871), .ZN(G75));
  OAI211_X1 g686(.A(new_n297), .B(new_n593), .C1(new_n865), .C2(new_n866), .ZN(new_n873));
  NOR2_X1   g687(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT55), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n587), .A2(new_n589), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n559), .A3(new_n582), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n878), .A2(new_n590), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT55), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n873), .A2(new_n880), .A3(new_n874), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n876), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n876), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n349), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n297), .B(new_n784), .C1(new_n865), .C2(new_n866), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n435), .B(KEYINPUT57), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n865), .A2(new_n866), .A3(new_n861), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n862), .B1(new_n859), .B2(new_n860), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n888), .B1(new_n892), .B2(new_n695), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n886), .B1(new_n893), .B2(new_n884), .ZN(new_n894));
  INV_X1    g708(.A(new_n884), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n863), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n897), .A2(new_n889), .B1(new_n693), .B2(new_n694), .ZN(new_n898));
  OAI211_X1 g712(.A(KEYINPUT122), .B(new_n895), .C1(new_n898), .C2(new_n888), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(G54));
  NOR2_X1   g714(.A1(new_n867), .A2(new_n298), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(new_n518), .A3(new_n510), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n510), .A2(new_n518), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .A4(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n903), .A2(new_n895), .A3(new_n905), .ZN(G60));
  NAND2_X1  g720(.A1(G478), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT59), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n864), .A2(new_n869), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n609), .A2(new_n610), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n897), .A2(new_n609), .A3(new_n610), .A4(new_n908), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n911), .A2(new_n895), .A3(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(new_n859), .A2(new_n860), .ZN(new_n914));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT123), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT60), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n356), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n884), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT61), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n914), .A2(new_n640), .A3(new_n917), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n919), .B(new_n922), .C1(new_n920), .C2(KEYINPUT61), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(G66));
  OAI21_X1  g740(.A(G953), .B1(new_n529), .B2(new_n554), .ZN(new_n927));
  INV_X1    g741(.A(new_n847), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(G953), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n877), .B1(G898), .B2(new_n349), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  AND2_X1   g745(.A1(new_n832), .A2(new_n664), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n686), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n789), .A2(new_n797), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n776), .A2(new_n673), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n937), .A2(new_n744), .A3(new_n301), .A4(new_n842), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n228), .A2(new_n232), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n489), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n349), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n826), .A2(new_n833), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n855), .B1(new_n788), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n789), .A2(new_n797), .A3(new_n945), .A4(new_n932), .ZN(new_n946));
  MUX2_X1   g760(.A(new_n650), .B(new_n946), .S(new_n349), .Z(new_n947));
  OAI21_X1  g761(.A(new_n943), .B1(new_n947), .B2(new_n942), .ZN(new_n948));
  OAI21_X1  g762(.A(G953), .B1(new_n415), .B2(new_n650), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G72));
  NAND2_X1  g764(.A1(G472), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT63), .Z(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT125), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n939), .B2(new_n847), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n678), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n946), .B2(new_n847), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n676), .A2(new_n259), .ZN(new_n959));
  OAI211_X1 g773(.A(KEYINPUT126), .B(new_n953), .C1(new_n946), .C2(new_n847), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n959), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n914), .A2(new_n677), .A3(new_n962), .A4(new_n952), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n955), .A2(new_n961), .A3(new_n895), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT127), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n884), .B1(new_n954), .B2(new_n678), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n966), .A2(new_n967), .A3(new_n961), .A4(new_n963), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n965), .A2(new_n968), .ZN(G57));
endmodule


