//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT26), .ZN(new_n205));
  AND3_X1   g004(.A1(new_n204), .A2(KEYINPUT68), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT68), .B1(new_n204), .B2(new_n205), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n202), .B(new_n203), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT27), .B(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT28), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT27), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G183gat), .ZN(new_n216));
  AND4_X1   g015(.A1(KEYINPUT28), .A2(new_n214), .A3(new_n216), .A4(new_n211), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n208), .B(new_n209), .C1(new_n212), .C2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT23), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n222), .A2(new_n224), .A3(new_n202), .ZN(new_n225));
  NOR2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n209), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT25), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT25), .A4(new_n202), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n209), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n227), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n226), .B1(KEYINPUT65), .B2(new_n229), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n238), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n232), .B1(new_n240), .B2(KEYINPUT66), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n236), .A2(new_n237), .A3(new_n242), .A4(new_n239), .ZN(new_n243));
  AOI211_X1 g042(.A(new_n219), .B(new_n231), .C1(new_n241), .C2(new_n243), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n234), .A2(new_n227), .A3(new_n235), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n229), .A2(KEYINPUT65), .ZN(new_n246));
  INV_X1    g045(.A(new_n226), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n239), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT66), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n232), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n243), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n231), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT67), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n218), .B1(new_n244), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G127gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G134gat), .ZN(new_n256));
  INV_X1    g055(.A(G134gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G127gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  INV_X1    g060(.A(G113gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(G120gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(G120gat), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n260), .A2(new_n267), .A3(KEYINPUT71), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n265), .A2(G113gat), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT1), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n256), .A2(KEYINPUT69), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n270), .A2(new_n271), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n254), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G227gat), .A2(G233gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n272), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n260), .A2(KEYINPUT71), .A3(new_n267), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT71), .B1(new_n260), .B2(new_n267), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n284), .B(new_n218), .C1(new_n244), .C2(new_n253), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT32), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT33), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G15gat), .B(G43gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT72), .ZN(new_n291));
  XNOR2_X1  g090(.A(G71gat), .B(G99gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n287), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n251), .A2(new_n252), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n219), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n231), .B1(new_n241), .B2(new_n243), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n284), .B1(new_n299), .B2(new_n218), .ZN(new_n300));
  INV_X1    g099(.A(new_n285), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n279), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT34), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n280), .B1(new_n278), .B2(new_n285), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT34), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n288), .B1(new_n293), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n307), .B2(new_n293), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n303), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT74), .B1(new_n294), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n304), .B(KEYINPUT34), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n287), .A2(new_n289), .A3(new_n293), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .A4(new_n310), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n310), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n306), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT75), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT79), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n284), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n281), .B(KEYINPUT79), .C1(new_n282), .C2(new_n283), .ZN(new_n328));
  XOR2_X1   g127(.A(G141gat), .B(G148gat), .Z(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(KEYINPUT2), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G141gat), .B(G148gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n333), .B(new_n332), .C1(new_n337), .C2(KEYINPUT2), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT3), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n336), .A2(new_n338), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n327), .A2(new_n328), .A3(new_n340), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(new_n284), .B2(new_n339), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n277), .A2(KEYINPUT4), .A3(new_n341), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n344), .A2(new_n345), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n327), .A2(new_n328), .A3(new_n339), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n277), .A2(new_n341), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n349), .B(KEYINPUT5), .C1(new_n352), .C2(new_n345), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT4), .B1(new_n277), .B2(new_n341), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n284), .A2(new_n346), .A3(new_n339), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n348), .A2(new_n347), .A3(KEYINPUT80), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT5), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n344), .A2(new_n360), .A3(new_n345), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT0), .ZN(new_n365));
  XNOR2_X1  g164(.A(G57gat), .B(G85gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n363), .A2(new_n368), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n362), .A3(new_n367), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G8gat), .B(G36gat), .Z(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT78), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n254), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n218), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n297), .A2(new_n382), .A3(KEYINPUT77), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n295), .B2(new_n218), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n379), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G197gat), .B(G204gat), .ZN(new_n387));
  INV_X1    g186(.A(G211gat), .ZN(new_n388));
  INV_X1    g187(.A(G218gat), .ZN(new_n389));
  OAI22_X1  g188(.A1(new_n388), .A2(new_n389), .B1(KEYINPUT76), .B2(KEYINPUT22), .ZN(new_n390));
  AND2_X1   g189(.A1(KEYINPUT76), .A2(KEYINPUT22), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n387), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G211gat), .B(G218gat), .Z(new_n393));
  AND2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(new_n393), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n381), .A2(new_n386), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT77), .B1(new_n297), .B2(new_n382), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n295), .A2(new_n384), .A3(new_n218), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n380), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n379), .B(new_n218), .C1(new_n244), .C2(new_n253), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n377), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  INV_X1    g203(.A(new_n396), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n381), .A2(new_n386), .A3(new_n396), .ZN(new_n407));
  INV_X1    g206(.A(new_n377), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n403), .A2(KEYINPUT30), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n406), .A2(new_n407), .A3(new_n411), .A4(new_n408), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n369), .A2(new_n373), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(G50gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n418), .B(KEYINPUT82), .Z(new_n419));
  OAI21_X1  g218(.A(new_n342), .B1(new_n396), .B2(KEYINPUT29), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n339), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n339), .A2(KEYINPUT3), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n396), .B1(new_n422), .B2(KEYINPUT29), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G22gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n423), .A3(G22gat), .ZN(new_n427));
  INV_X1    g226(.A(G228gat), .ZN(new_n428));
  INV_X1    g227(.A(G233gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n426), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n426), .B2(new_n427), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n419), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n427), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n430), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n418), .A2(KEYINPUT82), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n431), .A3(new_n427), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n440), .A2(KEYINPUT35), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n414), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n325), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n440), .B1(new_n319), .B2(new_n318), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n317), .A2(new_n413), .A3(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n445), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT84), .B1(new_n445), .B2(KEYINPUT35), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT38), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n406), .A2(new_n407), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT83), .B1(new_n450), .B2(KEYINPUT37), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n406), .A2(new_n407), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n408), .B1(new_n450), .B2(KEYINPUT37), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n449), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n373), .A2(new_n369), .A3(new_n409), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n404), .A2(new_n396), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n381), .A2(new_n386), .A3(new_n405), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT37), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n449), .A3(new_n377), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n451), .B2(new_n454), .ZN(new_n463));
  OR3_X1    g262(.A1(new_n457), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n344), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n357), .B2(new_n358), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(new_n345), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n352), .B2(new_n345), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n466), .B2(new_n345), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT40), .A4(new_n367), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n370), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n368), .B1(new_n467), .B2(new_n468), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT40), .B1(new_n474), .B2(new_n471), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n410), .A2(new_n412), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n440), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n464), .A2(new_n479), .B1(new_n414), .B2(new_n440), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n324), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n318), .B2(new_n319), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n317), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n448), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G85gat), .A2(G92gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT7), .ZN(new_n489));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490));
  INV_X1    g289(.A(G85gat), .ZN(new_n491));
  INV_X1    g290(.A(G92gat), .ZN(new_n492));
  AOI22_X1  g291(.A1(KEYINPUT8), .A2(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G99gat), .B(G106gat), .Z(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n495), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n489), .A3(new_n493), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(KEYINPUT98), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT98), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n494), .A2(new_n500), .A3(new_n495), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G50gat), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n504), .A2(G43gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(G43gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT15), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  OR2_X1    g307(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n510));
  AOI21_X1  g309(.A(G36gat), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT14), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n512), .A2(new_n513), .A3(G29gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n508), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n507), .B(KEYINPUT86), .C1(new_n511), .C2(new_n514), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g318(.A1(KEYINPUT87), .A2(KEYINPUT15), .ZN(new_n520));
  NAND2_X1  g319(.A1(KEYINPUT87), .A2(KEYINPUT15), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n520), .B(new_n521), .C1(new_n506), .C2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n505), .A2(new_n506), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(new_n522), .ZN(new_n525));
  INV_X1    g324(.A(new_n515), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT41), .ZN(new_n529));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT97), .Z(new_n531));
  OAI22_X1  g330(.A1(new_n503), .A2(new_n528), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT91), .B1(new_n528), .B2(KEYINPUT17), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n517), .A2(new_n518), .B1(new_n526), .B2(new_n525), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n502), .B1(new_n536), .B2(new_n534), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G190gat), .B(G218gat), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n540), .A2(new_n542), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n531), .A2(new_n529), .ZN(new_n546));
  XOR2_X1   g345(.A(G134gat), .B(G162gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  OAI22_X1  g347(.A1(new_n544), .A2(new_n545), .B1(KEYINPUT99), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n545), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n548), .B(KEYINPUT99), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n543), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT93), .ZN(new_n556));
  INV_X1    g355(.A(G57gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(G64gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(G64gat), .ZN(new_n559));
  INV_X1    g358(.A(G64gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT93), .A3(G57gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  OR2_X1    g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n562), .A2(new_n566), .A3(KEYINPUT94), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT94), .B1(new_n562), .B2(new_n566), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n560), .A2(G57gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n559), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n571), .A2(new_n572), .B1(new_n565), .B2(new_n563), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n572), .B2(new_n571), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n564), .A2(new_n563), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT21), .ZN(new_n579));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(KEYINPUT21), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT90), .ZN(new_n583));
  XNOR2_X1  g382(.A(G15gat), .B(G22gat), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n585));
  INV_X1    g384(.A(G1gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(KEYINPUT89), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n585), .A2(KEYINPUT16), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n586), .B1(new_n585), .B2(new_n587), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n583), .B(G8gat), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  INV_X1    g391(.A(G8gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(KEYINPUT90), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(KEYINPUT90), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n592), .A2(new_n595), .A3(new_n588), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n582), .A2(KEYINPUT96), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT96), .B1(new_n582), .B2(new_n598), .ZN(new_n600));
  OR3_X1    g399(.A1(new_n581), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n581), .B1(new_n599), .B2(new_n600), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT95), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n601), .A2(new_n602), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n601), .B2(new_n602), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n555), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n534), .A2(new_n536), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n598), .B(new_n613), .C1(new_n533), .C2(new_n537), .ZN(new_n614));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n591), .A2(new_n597), .A3(new_n534), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT18), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n614), .A2(KEYINPUT18), .A3(new_n615), .A4(new_n616), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n615), .B(KEYINPUT13), .Z(new_n621));
  INV_X1    g420(.A(new_n616), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n534), .B1(new_n591), .B2(new_n597), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G113gat), .B(G141gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G169gat), .B(G197gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n619), .A2(new_n620), .A3(new_n624), .A4(new_n631), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT101), .Z(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT100), .B(KEYINPUT10), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n496), .A2(new_n498), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n569), .A2(new_n644), .A3(new_n576), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI22_X1  g445(.A1(new_n569), .A2(new_n576), .B1(new_n499), .B2(new_n501), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n502), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n641), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n577), .A2(new_n502), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n641), .A3(new_n645), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n639), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n641), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n642), .B1(new_n651), .B2(new_n645), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n503), .A2(new_n577), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n655), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(new_n652), .A3(new_n638), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n612), .A2(new_n635), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n487), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n373), .A2(new_n369), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n478), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT102), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT16), .B(G8gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT103), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n668), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(G8gat), .ZN(new_n674));
  OR3_X1    g473(.A1(new_n669), .A2(new_n668), .A3(new_n672), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(G1325gat));
  INV_X1    g475(.A(new_n663), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n312), .A2(new_n316), .B1(new_n320), .B2(KEYINPUT75), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT36), .B1(new_n678), .B2(new_n323), .ZN(new_n679));
  INV_X1    g478(.A(new_n484), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT104), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n482), .A2(new_n682), .A3(new_n484), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G15gat), .B1(new_n677), .B2(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n324), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n677), .B2(new_n687), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n663), .A2(new_n440), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT105), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  AOI21_X1  g491(.A(new_n555), .B1(new_n448), .B2(new_n486), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n611), .A2(new_n635), .A3(new_n661), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(G29gat), .A3(new_n664), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT45), .Z(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT106), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n324), .A2(new_n414), .A3(new_n441), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n445), .A2(KEYINPUT35), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT84), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n445), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n440), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n474), .A2(new_n471), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT40), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n370), .A3(new_n472), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n706), .B1(new_n710), .B2(new_n477), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n457), .A2(new_n458), .A3(new_n463), .ZN(new_n712));
  OAI22_X1  g511(.A1(new_n711), .A2(new_n712), .B1(new_n413), .B2(new_n706), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n324), .A2(new_n481), .B1(new_n317), .B2(new_n483), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n554), .B1(new_n705), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT44), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n681), .A2(new_n480), .A3(new_n683), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n448), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n698), .A3(new_n554), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n699), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n694), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n664), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n697), .A2(new_n724), .ZN(G1328gat));
  NAND2_X1  g524(.A1(new_n478), .A2(new_n513), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  AOI211_X1 g526(.A(new_n726), .B(new_n695), .C1(new_n727), .C2(KEYINPUT46), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n695), .A2(new_n726), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G36gat), .B1(new_n723), .B2(new_n477), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT108), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(new_n735), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1329gat));
  NOR3_X1   g536(.A1(new_n695), .A2(G43gat), .A3(new_n324), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT109), .Z(new_n739));
  OAI21_X1  g538(.A(G43gat), .B1(new_n723), .B2(new_n685), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n739), .A2(KEYINPUT47), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(G1330gat));
  OAI21_X1  g544(.A(new_n504), .B1(new_n695), .B2(new_n706), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n440), .A2(G50gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n723), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n633), .A2(new_n634), .ZN(new_n750));
  INV_X1    g549(.A(new_n661), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n612), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n720), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n664), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT110), .B(G57gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1332gat));
  XNOR2_X1  g555(.A(new_n477), .B(KEYINPUT111), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  AND2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(G1333gat));
  NOR3_X1   g562(.A1(new_n753), .A2(G71gat), .A3(new_n324), .ZN(new_n764));
  INV_X1    g563(.A(new_n753), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n684), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n764), .B1(G71gat), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n440), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g569(.A1(new_n611), .A2(new_n750), .A3(new_n751), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n722), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n664), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n555), .B1(new_n719), .B2(new_n448), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n611), .A2(new_n750), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n780));
  NAND3_X1  g579(.A1(new_n774), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n751), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n491), .A3(new_n665), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n773), .A2(new_n783), .ZN(G1336gat));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n781), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n758), .A2(G92gat), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n785), .A2(new_n661), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(KEYINPUT52), .ZN(new_n788));
  OAI21_X1  g587(.A(G92gat), .B1(new_n772), .B2(new_n758), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n722), .A2(new_n478), .A3(new_n771), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n791), .A2(KEYINPUT113), .A3(G92gat), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT113), .B1(new_n791), .B2(G92gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(new_n787), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n790), .B1(new_n794), .B2(new_n795), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n772), .B2(new_n685), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n324), .A2(G99gat), .A3(new_n751), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n785), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1338gat));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  INV_X1    g600(.A(G106gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n802), .A3(new_n440), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT114), .B1(new_n772), .B2(new_n706), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G106gat), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n772), .A2(KEYINPUT114), .A3(new_n706), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n801), .B(new_n803), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G106gat), .B1(new_n772), .B2(new_n706), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n803), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT53), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(G1339gat));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n648), .A2(new_n641), .A3(new_n649), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n659), .A2(new_n813), .A3(KEYINPUT54), .ZN(new_n814));
  XNOR2_X1  g613(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n639), .B1(new_n659), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n812), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n638), .B1(new_n650), .B2(new_n815), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n659), .A2(new_n813), .A3(KEYINPUT54), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n818), .A2(new_n660), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n750), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n622), .A2(new_n623), .A3(new_n621), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n630), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n634), .A2(new_n661), .A3(new_n826), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT117), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(KEYINPUT117), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n823), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n555), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n634), .A2(new_n826), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(KEYINPUT116), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n833), .A2(new_n554), .A3(new_n834), .A4(new_n822), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n611), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n612), .A2(new_n750), .A3(new_n661), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n440), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n839), .A2(new_n665), .A3(new_n325), .A4(new_n758), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(KEYINPUT118), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(G113gat), .A3(new_n750), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n838), .A2(new_n664), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n317), .A2(new_n444), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n847), .A3(new_n758), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n262), .B1(new_n848), .B2(new_n635), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n844), .A2(new_n849), .ZN(G1340gat));
  NAND3_X1  g649(.A1(new_n843), .A2(G120gat), .A3(new_n661), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n265), .B1(new_n848), .B2(new_n751), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(G1341gat));
  AOI21_X1  g652(.A(new_n255), .B1(new_n843), .B2(new_n611), .ZN(new_n854));
  INV_X1    g653(.A(new_n611), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n848), .A2(G127gat), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n854), .A2(new_n856), .ZN(G1342gat));
  NOR2_X1   g656(.A1(new_n555), .A2(new_n478), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n845), .A2(new_n257), .A3(new_n847), .A4(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n861), .A2(new_n862), .B1(new_n863), .B2(KEYINPUT56), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(KEYINPUT121), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n863), .B(KEYINPUT56), .C1(new_n861), .C2(new_n862), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n841), .A2(new_n842), .A3(new_n554), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n868), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT120), .B1(new_n868), .B2(G134gat), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n866), .B(new_n867), .C1(new_n869), .C2(new_n870), .ZN(G1343gat));
  NOR2_X1   g670(.A1(new_n684), .A2(new_n706), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n845), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n757), .ZN(new_n874));
  INV_X1    g673(.A(G141gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n750), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n684), .A2(new_n664), .A3(new_n757), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n440), .B1(new_n836), .B2(new_n837), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(KEYINPUT122), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n706), .A2(new_n879), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n634), .A2(new_n883), .A3(new_n661), .A4(new_n826), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n827), .A2(KEYINPUT123), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n818), .A2(new_n660), .A3(new_n821), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n884), .B(new_n885), .C1(new_n635), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n555), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n835), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n837), .B1(new_n889), .B2(new_n855), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n880), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT122), .B1(new_n878), .B2(new_n879), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n877), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n635), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n876), .B1(new_n894), .B2(new_n875), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT58), .ZN(G1344gat));
  OAI21_X1  g695(.A(new_n881), .B1(new_n836), .B2(new_n837), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n822), .A2(new_n750), .B1(KEYINPUT123), .B2(new_n827), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n554), .B1(new_n898), .B2(new_n884), .ZN(new_n899));
  INV_X1    g698(.A(new_n835), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n855), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n837), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n706), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n897), .B1(new_n903), .B2(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n661), .ZN(new_n905));
  INV_X1    g704(.A(new_n877), .ZN(new_n906));
  OAI21_X1  g705(.A(G148gat), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT59), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n661), .B(new_n877), .C1(new_n891), .C2(new_n892), .ZN(new_n909));
  INV_X1    g708(.A(G148gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(KEYINPUT59), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n909), .A2(KEYINPUT124), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT124), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n874), .A2(new_n910), .A3(new_n661), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(G155gat), .B1(new_n893), .B2(new_n855), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n874), .A2(new_n330), .A3(new_n611), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n893), .B2(new_n555), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n858), .A2(new_n331), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n873), .B2(new_n921), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n665), .A2(new_n477), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n839), .A2(new_n325), .A3(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n220), .A3(new_n635), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n838), .A2(new_n665), .A3(new_n758), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(new_n847), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n750), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n928), .B2(new_n220), .ZN(G1348gat));
  NOR3_X1   g728(.A1(new_n924), .A2(new_n221), .A3(new_n751), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n661), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n221), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n927), .A2(new_n210), .A3(new_n611), .ZN(new_n933));
  OAI21_X1  g732(.A(G183gat), .B1(new_n924), .B2(new_n855), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n924), .B2(new_n555), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT61), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n211), .A3(new_n554), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1351gat));
  NAND2_X1  g739(.A1(new_n926), .A2(new_n872), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n750), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n681), .A2(new_n683), .A3(new_n923), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n879), .B1(new_n890), .B2(new_n706), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n897), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(G197gat), .A3(new_n750), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n943), .A2(new_n947), .ZN(G1352gat));
  INV_X1    g747(.A(G204gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n661), .A2(new_n949), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n941), .A2(new_n950), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g750(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n952));
  INV_X1    g751(.A(new_n944), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n904), .A2(new_n661), .A3(new_n953), .ZN(new_n954));
  AOI22_X1  g753(.A1(new_n951), .A2(new_n952), .B1(G204gat), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n955), .B1(new_n951), .B2(new_n952), .ZN(G1353gat));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n904), .A2(new_n958), .A3(new_n611), .A4(new_n953), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n946), .B2(new_n611), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n904), .A2(new_n611), .A3(new_n953), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n959), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n942), .A2(new_n388), .A3(new_n611), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT127), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n970), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1354gat));
  NOR3_X1   g771(.A1(new_n941), .A2(G218gat), .A3(new_n555), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n389), .B1(new_n946), .B2(new_n554), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n973), .A2(new_n974), .ZN(G1355gat));
endmodule


