

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  NOR2_X1 U323 ( .A1(n426), .A2(n425), .ZN(n427) );
  XOR2_X1 U324 ( .A(n357), .B(n356), .Z(n517) );
  XNOR2_X1 U325 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n456) );
  XNOR2_X1 U326 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U327 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n462) );
  XNOR2_X1 U328 ( .A(n348), .B(G92GAT), .ZN(n349) );
  XNOR2_X1 U329 ( .A(n463), .B(n462), .ZN(n522) );
  XNOR2_X1 U330 ( .A(n350), .B(n349), .ZN(n353) );
  NOR2_X1 U331 ( .A1(n514), .A2(n466), .ZN(n564) );
  NOR2_X1 U332 ( .A1(n525), .A2(n470), .ZN(n561) );
  XOR2_X1 U333 ( .A(KEYINPUT79), .B(n548), .Z(n536) );
  XOR2_X1 U334 ( .A(KEYINPUT110), .B(n447), .Z(n520) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n471) );
  XNOR2_X1 U336 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U337 ( .A(n472), .B(n471), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n292) );
  XNOR2_X1 U339 ( .A(G113GAT), .B(G197GAT), .ZN(n291) );
  XNOR2_X1 U340 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U341 ( .A(G50GAT), .B(G36GAT), .Z(n294) );
  XOR2_X1 U342 ( .A(G141GAT), .B(G22GAT), .Z(n391) );
  XOR2_X1 U343 ( .A(G169GAT), .B(G8GAT), .Z(n351) );
  XNOR2_X1 U344 ( .A(n391), .B(n351), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U346 ( .A(n296), .B(n295), .Z(n298) );
  NAND2_X1 U347 ( .A1(G229GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U349 ( .A(n299), .B(KEYINPUT30), .Z(n302) );
  XNOR2_X1 U350 ( .A(G15GAT), .B(G1GAT), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n300), .B(KEYINPUT71), .ZN(n327) );
  XNOR2_X1 U352 ( .A(n327), .B(KEYINPUT29), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U354 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n304) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G29GAT), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U357 ( .A(KEYINPUT70), .B(n305), .Z(n440) );
  XNOR2_X1 U358 ( .A(n306), .B(n440), .ZN(n565) );
  XOR2_X1 U359 ( .A(G92GAT), .B(G85GAT), .Z(n308) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G106GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n432) );
  XOR2_X1 U362 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n310) );
  XNOR2_X1 U363 ( .A(G204GAT), .B(KEYINPUT72), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U365 ( .A(n432), .B(n311), .Z(n313) );
  XOR2_X1 U366 ( .A(G120GAT), .B(G71GAT), .Z(n403) );
  XOR2_X1 U367 ( .A(G148GAT), .B(G78GAT), .Z(n390) );
  XNOR2_X1 U368 ( .A(n403), .B(n390), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n320) );
  XOR2_X1 U370 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n315) );
  NAND2_X1 U371 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U373 ( .A(n316), .B(KEYINPUT74), .Z(n318) );
  XOR2_X1 U374 ( .A(G57GAT), .B(KEYINPUT13), .Z(n323) );
  XOR2_X1 U375 ( .A(G176GAT), .B(G64GAT), .Z(n344) );
  XNOR2_X1 U376 ( .A(n323), .B(n344), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U378 ( .A(n320), .B(n319), .Z(n571) );
  XNOR2_X1 U379 ( .A(n571), .B(KEYINPUT41), .ZN(n557) );
  NAND2_X1 U380 ( .A1(n565), .A2(n557), .ZN(n504) );
  INV_X1 U381 ( .A(n504), .ZN(n446) );
  XNOR2_X1 U382 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n445) );
  XOR2_X1 U383 ( .A(G78GAT), .B(G71GAT), .Z(n322) );
  XNOR2_X1 U384 ( .A(G183GAT), .B(G127GAT), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U386 ( .A(n324), .B(n323), .Z(n326) );
  XNOR2_X1 U387 ( .A(G22GAT), .B(G155GAT), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n326), .B(n325), .ZN(n331) );
  XOR2_X1 U389 ( .A(n327), .B(KEYINPUT12), .Z(n329) );
  NAND2_X1 U390 ( .A1(G231GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U392 ( .A(n331), .B(n330), .Z(n339) );
  XOR2_X1 U393 ( .A(KEYINPUT82), .B(G64GAT), .Z(n333) );
  XNOR2_X1 U394 ( .A(G8GAT), .B(G211GAT), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U396 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n335) );
  XNOR2_X1 U397 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n560) );
  XOR2_X1 U401 ( .A(G183GAT), .B(KEYINPUT17), .Z(n341) );
  XNOR2_X1 U402 ( .A(KEYINPUT18), .B(KEYINPUT86), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n343) );
  XOR2_X1 U404 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n342) );
  XNOR2_X1 U405 ( .A(n343), .B(n342), .ZN(n413) );
  INV_X1 U406 ( .A(n413), .ZN(n357) );
  XOR2_X1 U407 ( .A(G36GAT), .B(G190GAT), .Z(n428) );
  XNOR2_X1 U408 ( .A(n344), .B(n428), .ZN(n355) );
  XOR2_X1 U409 ( .A(G204GAT), .B(G211GAT), .Z(n346) );
  XNOR2_X1 U410 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n345) );
  XNOR2_X1 U411 ( .A(n346), .B(n345), .ZN(n388) );
  INV_X1 U412 ( .A(KEYINPUT93), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n388), .B(n347), .ZN(n350) );
  NAND2_X1 U414 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XOR2_X1 U415 ( .A(n351), .B(G218GAT), .Z(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n356) );
  INV_X1 U418 ( .A(n517), .ZN(n464) );
  XOR2_X1 U419 ( .A(KEYINPUT27), .B(n464), .Z(n420) );
  XOR2_X1 U420 ( .A(G127GAT), .B(KEYINPUT0), .Z(n359) );
  XNOR2_X1 U421 ( .A(G113GAT), .B(G134GAT), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n407) );
  XOR2_X1 U423 ( .A(KEYINPUT92), .B(n407), .Z(n361) );
  NAND2_X1 U424 ( .A1(G225GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n376) );
  XOR2_X1 U426 ( .A(G85GAT), .B(G162GAT), .Z(n363) );
  XNOR2_X1 U427 ( .A(G29GAT), .B(G120GAT), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U429 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n365) );
  XNOR2_X1 U430 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U432 ( .A(n367), .B(n366), .Z(n374) );
  XOR2_X1 U433 ( .A(G155GAT), .B(KEYINPUT2), .Z(n369) );
  XNOR2_X1 U434 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n369), .B(n368), .ZN(n385) );
  XOR2_X1 U436 ( .A(G57GAT), .B(G148GAT), .Z(n371) );
  XNOR2_X1 U437 ( .A(G1GAT), .B(G141GAT), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n385), .B(n372), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n514) );
  NAND2_X1 U442 ( .A1(n420), .A2(n514), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n377), .B(KEYINPUT94), .ZN(n523) );
  XNOR2_X1 U444 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n396) );
  XOR2_X1 U445 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n379) );
  XNOR2_X1 U446 ( .A(G106GAT), .B(KEYINPUT24), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n379), .B(n378), .ZN(n395) );
  XOR2_X1 U448 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n381) );
  NAND2_X1 U449 ( .A1(G228GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U450 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U451 ( .A(n382), .B(KEYINPUT91), .Z(n387) );
  XOR2_X1 U452 ( .A(G162GAT), .B(KEYINPUT76), .Z(n384) );
  XNOR2_X1 U453 ( .A(G50GAT), .B(G218GAT), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n429) );
  XNOR2_X1 U455 ( .A(n429), .B(n385), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n389) );
  XOR2_X1 U457 ( .A(n389), .B(n388), .Z(n393) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n467) );
  XNOR2_X1 U461 ( .A(n396), .B(n467), .ZN(n528) );
  NOR2_X1 U462 ( .A1(n523), .A2(n528), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n397), .B(KEYINPUT95), .ZN(n414) );
  XOR2_X1 U464 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n399) );
  XNOR2_X1 U465 ( .A(G169GAT), .B(G15GAT), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n411) );
  XOR2_X1 U467 ( .A(G176GAT), .B(G99GAT), .Z(n401) );
  XNOR2_X1 U468 ( .A(G43GAT), .B(G190GAT), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U470 ( .A(n403), .B(n402), .Z(n405) );
  NAND2_X1 U471 ( .A1(G227GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U472 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U473 ( .A(n406), .B(KEYINPUT20), .Z(n409) );
  XNOR2_X1 U474 ( .A(n407), .B(KEYINPUT84), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X2 U477 ( .A(n413), .B(n412), .ZN(n519) );
  NOR2_X1 U478 ( .A1(n414), .A2(n519), .ZN(n426) );
  INV_X1 U479 ( .A(n467), .ZN(n416) );
  INV_X1 U480 ( .A(n519), .ZN(n525) );
  NOR2_X1 U481 ( .A1(n525), .A2(n464), .ZN(n415) );
  NOR2_X1 U482 ( .A1(n416), .A2(n415), .ZN(n418) );
  XNOR2_X1 U483 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n422) );
  NOR2_X1 U485 ( .A1(n467), .A2(n519), .ZN(n419) );
  XNOR2_X1 U486 ( .A(n419), .B(KEYINPUT26), .ZN(n563) );
  NAND2_X1 U487 ( .A1(n420), .A2(n563), .ZN(n421) );
  NAND2_X1 U488 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U489 ( .A(KEYINPUT97), .B(n423), .ZN(n424) );
  NOR2_X1 U490 ( .A1(n514), .A2(n424), .ZN(n425) );
  XOR2_X1 U491 ( .A(KEYINPUT98), .B(n427), .Z(n475) );
  XOR2_X1 U492 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n431) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n432), .B(G134GAT), .ZN(n434) );
  NAND2_X1 U496 ( .A1(G232GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U497 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n442) );
  XOR2_X1 U499 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n438) );
  XNOR2_X1 U500 ( .A(KEYINPUT78), .B(KEYINPUT9), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n548) );
  XNOR2_X1 U504 ( .A(KEYINPUT36), .B(n536), .ZN(n580) );
  NAND2_X1 U505 ( .A1(n475), .A2(n580), .ZN(n443) );
  NOR2_X1 U506 ( .A1(n560), .A2(n443), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n445), .B(n444), .ZN(n486) );
  NAND2_X1 U508 ( .A1(n446), .A2(n486), .ZN(n447) );
  NAND2_X1 U509 ( .A1(n520), .A2(n528), .ZN(n451) );
  XOR2_X1 U510 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n449) );
  INV_X1 U511 ( .A(G106GAT), .ZN(n448) );
  XNOR2_X1 U512 ( .A(n451), .B(n450), .ZN(G1339GAT) );
  XOR2_X1 U513 ( .A(KEYINPUT118), .B(KEYINPUT55), .Z(n469) );
  INV_X1 U514 ( .A(n565), .ZN(n551) );
  NAND2_X1 U515 ( .A1(n551), .A2(n557), .ZN(n452) );
  XNOR2_X1 U516 ( .A(KEYINPUT46), .B(n452), .ZN(n454) );
  NOR2_X1 U517 ( .A1(n548), .A2(n560), .ZN(n453) );
  NAND2_X1 U518 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U519 ( .A(n455), .B(KEYINPUT47), .ZN(n461) );
  NAND2_X1 U520 ( .A1(n580), .A2(n560), .ZN(n457) );
  NAND2_X1 U521 ( .A1(n458), .A2(n571), .ZN(n459) );
  NOR2_X1 U522 ( .A1(n459), .A2(n551), .ZN(n460) );
  NOR2_X1 U523 ( .A1(n461), .A2(n460), .ZN(n463) );
  NOR2_X1 U524 ( .A1(n522), .A2(n464), .ZN(n465) );
  XOR2_X1 U525 ( .A(KEYINPUT54), .B(n465), .Z(n466) );
  NAND2_X1 U526 ( .A1(n564), .A2(n467), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n561), .A2(n536), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n571), .A2(n551), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT75), .ZN(n487) );
  INV_X1 U531 ( .A(n487), .ZN(n477) );
  INV_X1 U532 ( .A(n560), .ZN(n576) );
  NOR2_X1 U533 ( .A1(n536), .A2(n576), .ZN(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT16), .B(n474), .ZN(n476) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n503) );
  NOR2_X1 U536 ( .A1(n477), .A2(n503), .ZN(n484) );
  NAND2_X1 U537 ( .A1(n514), .A2(n484), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(KEYINPUT34), .ZN(n479) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  XOR2_X1 U540 ( .A(G8GAT), .B(KEYINPUT99), .Z(n481) );
  NAND2_X1 U541 ( .A1(n484), .A2(n517), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT35), .Z(n483) );
  NAND2_X1 U544 ( .A1(n484), .A2(n519), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NAND2_X1 U546 ( .A1(n528), .A2(n484), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n485), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n492) );
  NAND2_X1 U549 ( .A1(n487), .A2(n486), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n488), .B(KEYINPUT38), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n499) );
  NAND2_X1 U553 ( .A1(n499), .A2(n514), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(n493), .ZN(G1328GAT) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n495) );
  NAND2_X1 U557 ( .A1(n517), .A2(n499), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(G1329GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n497) );
  NAND2_X1 U560 ( .A1(n499), .A2(n519), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n501) );
  NAND2_X1 U564 ( .A1(n499), .A2(n528), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n502), .ZN(G1331GAT) );
  NOR2_X1 U567 ( .A1(n504), .A2(n503), .ZN(n511) );
  NAND2_X1 U568 ( .A1(n514), .A2(n511), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(KEYINPUT42), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n511), .A2(n517), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT109), .Z(n510) );
  NAND2_X1 U575 ( .A1(n511), .A2(n519), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U578 ( .A1(n511), .A2(n528), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  XOR2_X1 U580 ( .A(G85GAT), .B(KEYINPUT111), .Z(n516) );
  NAND2_X1 U581 ( .A1(n520), .A2(n514), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n517), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(G113GAT), .B(KEYINPUT115), .Z(n530) );
  NOR2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(KEYINPUT113), .ZN(n540) );
  NOR2_X1 U590 ( .A1(n525), .A2(n540), .ZN(n526) );
  XOR2_X1 U591 ( .A(KEYINPUT114), .B(n526), .Z(n527) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n537), .A2(n551), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U596 ( .A1(n537), .A2(n557), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n534) );
  NAND2_X1 U599 ( .A1(n537), .A2(n560), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n535), .Z(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  INV_X1 U605 ( .A(n563), .ZN(n541) );
  NOR2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n551), .A2(n549), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n544) );
  NAND2_X1 U610 ( .A1(n549), .A2(n557), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .Z(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n549), .A2(n560), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U618 ( .A(G169GAT), .B(KEYINPUT119), .Z(n553) );
  NAND2_X1 U619 ( .A1(n561), .A2(n551), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(n556), .Z(n559) );
  NAND2_X1 U625 ( .A1(n561), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n579) );
  NOR2_X1 U630 ( .A1(n565), .A2(n579), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT59), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n579), .A2(n571), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n579), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(n577), .Z(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n583) );
  INV_X1 U645 ( .A(n579), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

