//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948;
  XOR2_X1   g000(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G43gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n209), .A2(G43gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT14), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n214), .A2(new_n215), .ZN(new_n220));
  OR3_X1    g019(.A1(new_n213), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n212), .B1(new_n222), .B2(new_n210), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n209), .A2(KEYINPUT91), .A3(G43gat), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT15), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT89), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n219), .A2(new_n227), .B1(new_n214), .B2(new_n215), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT89), .B1(new_n216), .B2(new_n218), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n213), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT90), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(KEYINPUT90), .B(new_n213), .C1(new_n228), .C2(new_n229), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n226), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT17), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT94), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT94), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n237), .A3(KEYINPUT17), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G15gat), .B(G22gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT93), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT16), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n242), .A2(G1gat), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n241), .A2(G1gat), .ZN(new_n245));
  OR3_X1    g044(.A1(new_n244), .A2(new_n245), .A3(G8gat), .ZN(new_n246));
  OAI21_X1  g045(.A(G8gat), .B1(new_n244), .B2(new_n245), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n250));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n239), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G229gat), .A2(G233gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n234), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT18), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n253), .A2(KEYINPUT18), .A3(new_n254), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n249), .A2(new_n234), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n256), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n254), .B(KEYINPUT13), .Z(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND4_X1   g063(.A1(new_n208), .A2(new_n259), .A3(new_n260), .A4(new_n264), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n257), .A2(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n208), .B1(new_n266), .B2(new_n260), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT66), .B(G190gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT27), .B(G183gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT28), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(KEYINPUT68), .A3(G183gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT27), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n270), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n272), .B1(new_n278), .B2(KEYINPUT28), .ZN(new_n279));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  INV_X1    g079(.A(G169gat), .ZN(new_n281));
  INV_X1    g080(.A(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n283), .B2(KEYINPUT26), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n279), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT23), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n293), .A2(KEYINPUT25), .A3(new_n280), .A4(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT66), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G190gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT67), .B1(new_n300), .B2(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n270), .A2(new_n302), .A3(new_n276), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT65), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(new_n288), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n295), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n280), .A3(new_n294), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT64), .B1(new_n289), .B2(KEYINPUT24), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT64), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n276), .A2(new_n296), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n311), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT25), .B1(new_n310), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n291), .B1(new_n308), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G113gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT69), .B(G113gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(new_n320), .ZN(new_n323));
  INV_X1    g122(.A(G134gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G127gat), .ZN(new_n325));
  OR2_X1    g124(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n326));
  INV_X1    g125(.A(G127gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G134gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n329));
  AND4_X1   g128(.A1(new_n325), .A2(new_n326), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n320), .A2(G113gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n320), .A2(G113gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n325), .A2(new_n328), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n323), .A2(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n269), .B1(new_n319), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n302), .B1(new_n270), .B2(new_n276), .ZN(new_n339));
  AND4_X1   g138(.A1(new_n302), .A2(new_n297), .A3(new_n299), .A4(new_n276), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n307), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n295), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n315), .B(new_n316), .C1(new_n312), .C2(new_n313), .ZN(new_n345));
  INV_X1    g144(.A(new_n314), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n344), .B1(new_n347), .B2(new_n309), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n343), .A2(new_n348), .B1(new_n279), .B2(new_n290), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(KEYINPUT71), .A3(new_n336), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n349), .B2(new_n336), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n319), .A2(KEYINPUT72), .A3(new_n337), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n338), .A2(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G227gat), .A2(G233gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT32), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT33), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n354), .B2(new_n355), .ZN(new_n358));
  XOR2_X1   g157(.A(G15gat), .B(G43gat), .Z(new_n359));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n354), .A2(new_n355), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT34), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT34), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n354), .A2(new_n365), .A3(new_n355), .ZN(new_n366));
  INV_X1    g165(.A(new_n361), .ZN(new_n367));
  OAI221_X1 g166(.A(KEYINPUT32), .B1(new_n357), .B2(new_n367), .C1(new_n354), .C2(new_n355), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n362), .A2(new_n364), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n362), .A2(new_n368), .B1(new_n366), .B2(new_n364), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n349), .B2(KEYINPUT29), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT74), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n349), .B2(new_n373), .ZN(new_n376));
  XNOR2_X1  g175(.A(G197gat), .B(G204gat), .ZN(new_n377));
  INV_X1    g176(.A(G211gat), .ZN(new_n378));
  INV_X1    g177(.A(G218gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n377), .B1(KEYINPUT22), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G211gat), .B(G218gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n373), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n319), .A2(KEYINPUT74), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n374), .A2(new_n376), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n319), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n349), .A2(new_n373), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n383), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(G64gat), .ZN(new_n393));
  INV_X1    g192(.A(G92gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n387), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n387), .B2(new_n391), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n387), .A2(new_n391), .ZN(new_n400));
  INV_X1    g199(.A(new_n395), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n400), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G162gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G155gat), .ZN(new_n406));
  INV_X1    g205(.A(G155gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G162gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G141gat), .B(G148gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT76), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(KEYINPUT76), .B(new_n409), .C1(new_n410), .C2(new_n411), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT77), .B(G141gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G148gat), .ZN(new_n417));
  INV_X1    g216(.A(G141gat), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT78), .B1(new_n418), .B2(G148gat), .ZN(new_n419));
  OR3_X1    g218(.A1(new_n418), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT2), .B1(new_n405), .B2(KEYINPUT79), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n422), .A2(new_n406), .A3(new_n408), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n414), .A2(new_n415), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n384), .B1(new_n426), .B2(new_n388), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n427), .A2(KEYINPUT83), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(KEYINPUT83), .ZN(new_n429));
  INV_X1    g228(.A(G228gat), .ZN(new_n430));
  INV_X1    g229(.A(G233gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n425), .B1(new_n383), .B2(KEYINPUT29), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n416), .A2(G148gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n420), .A2(new_n419), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n423), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n415), .ZN(new_n436));
  OR2_X1    g235(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n437));
  NAND2_X1  g236(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n418), .A2(G148gat), .ZN(new_n439));
  INV_X1    g238(.A(G148gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(G141gat), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT76), .B1(new_n442), .B2(new_n409), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n435), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  AOI211_X1 g243(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n384), .A2(new_n388), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n424), .B1(new_n447), .B2(new_n425), .ZN(new_n448));
  OAI22_X1  g247(.A1(new_n448), .A2(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT31), .B(G50gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n451), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n446), .A2(new_n453), .A3(new_n449), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G78gat), .B(G106gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(G22gat), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n452), .A2(new_n457), .A3(new_n454), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n372), .A2(new_n404), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n337), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n336), .B(new_n435), .C1(new_n443), .C2(new_n436), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT81), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT5), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n463), .ZN(new_n469));
  INV_X1    g268(.A(new_n465), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n414), .A2(new_n415), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n336), .B1(new_n471), .B2(new_n435), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n467), .B(new_n469), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT82), .B1(new_n468), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n469), .B1(new_n470), .B2(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT81), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT5), .A4(new_n473), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n336), .B1(new_n444), .B2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT4), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT4), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n424), .A2(new_n482), .A3(new_n336), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n426), .A2(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT80), .A3(new_n463), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n480), .A2(new_n426), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n483), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n463), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n475), .A2(new_n479), .A3(new_n485), .A4(new_n490), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n488), .A2(KEYINPUT5), .ZN(new_n492));
  XNOR2_X1  g291(.A(G1gat), .B(G29gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT0), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(G57gat), .ZN(new_n495));
  INV_X1    g294(.A(G85gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n491), .B2(new_n492), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI211_X1 g301(.A(new_n499), .B(new_n497), .C1(new_n491), .C2(new_n492), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n462), .A2(KEYINPUT35), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT35), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n372), .A2(new_n404), .A3(new_n461), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(new_n504), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n492), .ZN(new_n511));
  INV_X1    g310(.A(new_n497), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT84), .B1(new_n484), .B2(new_n463), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n486), .A2(new_n487), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT84), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n469), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT39), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n470), .A2(new_n472), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n519), .B1(new_n521), .B2(new_n463), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(new_n517), .A3(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n520), .A2(KEYINPUT40), .A3(new_n497), .A4(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT40), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n497), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT39), .B1(new_n514), .B2(new_n517), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n403), .A2(new_n513), .A3(new_n524), .A4(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT85), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n497), .A3(new_n523), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n525), .A2(new_n532), .B1(new_n511), .B2(new_n512), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(KEYINPUT85), .A3(new_n403), .A4(new_n524), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT38), .ZN(new_n536));
  XOR2_X1   g335(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n537));
  OAI211_X1 g336(.A(new_n536), .B(new_n401), .C1(new_n400), .C2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n374), .A2(new_n376), .A3(new_n386), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n383), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT86), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(KEYINPUT86), .A3(new_n383), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n389), .A2(new_n390), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n542), .B(new_n543), .C1(new_n383), .C2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n538), .B1(new_n545), .B2(KEYINPUT37), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n400), .A2(new_n537), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n395), .B1(new_n400), .B2(KEYINPUT37), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n536), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n546), .A2(new_n396), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n503), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n513), .A2(new_n499), .A3(new_n498), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n461), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n404), .B1(new_n502), .B2(new_n503), .ZN(new_n555));
  INV_X1    g354(.A(new_n461), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(new_n370), .B2(new_n371), .ZN(new_n558));
  INV_X1    g357(.A(new_n371), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(KEYINPUT36), .A3(new_n369), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n555), .A2(new_n556), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n268), .B1(new_n510), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564));
  AND2_X1   g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(KEYINPUT41), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n564), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G99gat), .B(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT7), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(KEYINPUT8), .A2(new_n573), .B1(new_n496), .B2(new_n394), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n568), .B(KEYINPUT97), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n570), .A2(new_n575), .A3(KEYINPUT98), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n255), .A2(new_n583), .B1(KEYINPUT41), .B2(new_n565), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n236), .A2(new_n238), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT99), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n583), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n252), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n584), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n567), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n584), .B(new_n592), .C1(new_n585), .C2(new_n588), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT100), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n584), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n583), .B(KEYINPUT99), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n251), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n598), .B2(new_n239), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT100), .B1(new_n599), .B2(new_n592), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n591), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(KEYINPUT102), .B(new_n591), .C1(new_n595), .C2(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n593), .A2(new_n594), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n599), .A2(KEYINPUT100), .A3(new_n592), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT101), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n590), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT101), .B1(new_n606), .B2(new_n607), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n567), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  XOR2_X1   g418(.A(G57gat), .B(G64gat), .Z(new_n620));
  INV_X1    g419(.A(KEYINPUT9), .ZN(new_n621));
  INV_X1    g420(.A(G71gat), .ZN(new_n622));
  INV_X1    g421(.A(G78gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G71gat), .B(G78gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  OAI21_X1  g426(.A(new_n249), .B1(new_n619), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT96), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n619), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT95), .Z(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n629), .A2(new_n633), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n618), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n634), .A3(new_n617), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n627), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n583), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n627), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n576), .A3(new_n579), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n581), .A2(new_n627), .A3(new_n582), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n641), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n648), .ZN(new_n653));
  INV_X1    g452(.A(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT105), .B(G204gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT104), .B(G176gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n659), .B(new_n660), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n661), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n652), .A2(new_n655), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n605), .A2(new_n612), .A3(new_n640), .A4(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n595), .B2(new_n600), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n608), .A3(new_n609), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n672), .A2(new_n567), .B1(new_n603), .B2(new_n604), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n673), .A2(KEYINPUT106), .A3(new_n640), .A4(new_n666), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n563), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n505), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g477(.A1(new_n676), .A2(new_n404), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  AND2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(KEYINPUT42), .ZN(new_n683));
  INV_X1    g482(.A(G8gat), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n679), .ZN(G1325gat));
  NAND2_X1  g484(.A1(new_n558), .A2(new_n560), .ZN(new_n686));
  OAI21_X1  g485(.A(G15gat), .B1(new_n676), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n372), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n676), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n676), .A2(new_n461), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT107), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n691), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(new_n640), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n605), .A2(new_n612), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n563), .A2(new_n695), .A3(new_n696), .A4(new_n666), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n697), .A2(G29gat), .A3(new_n505), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT45), .Z(new_n699));
  AND3_X1   g498(.A1(new_n554), .A2(KEYINPUT108), .A3(new_n561), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT108), .B1(new_n554), .B2(new_n561), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n510), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n702), .B2(new_n696), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n696), .A2(KEYINPUT44), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n510), .B2(new_n562), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n268), .A2(new_n640), .A3(new_n665), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n505), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n699), .A2(new_n709), .ZN(G1328gat));
  NOR3_X1   g509(.A1(new_n697), .A2(G36gat), .A3(new_n404), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n708), .B2(new_n404), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(new_n686), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n706), .A2(new_n715), .A3(new_n707), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G43gat), .ZN(new_n717));
  OR3_X1    g516(.A1(new_n697), .A2(G43gat), .A3(new_n688), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n717), .A2(new_n718), .B1(KEYINPUT109), .B2(KEYINPUT47), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n708), .B2(new_n461), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT48), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n556), .A2(new_n209), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n722), .B1(new_n697), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n724), .B(new_n726), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n506), .A2(new_n509), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n562), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n554), .A2(KEYINPUT108), .A3(new_n561), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n673), .A2(new_n268), .A3(new_n640), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n732), .A2(new_n666), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n504), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n403), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  NAND2_X1  g539(.A1(new_n734), .A2(new_n715), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G71gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n734), .A2(new_n622), .A3(new_n372), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT111), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n556), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  INV_X1    g550(.A(new_n268), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n640), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n706), .A2(new_n665), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n505), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT112), .B1(new_n732), .B2(new_n673), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n702), .A2(new_n757), .A3(new_n696), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n753), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n753), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n702), .A2(new_n696), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(KEYINPUT112), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT51), .B1(new_n764), .B2(new_n758), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n665), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n504), .A2(new_n496), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n755), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  NOR4_X1   g567(.A1(new_n703), .A2(new_n666), .A3(new_n705), .A4(new_n762), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n394), .B1(new_n769), .B2(new_n403), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(KEYINPUT52), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n761), .A2(new_n765), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n665), .A2(new_n394), .A3(new_n403), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT113), .Z(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT114), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n764), .A2(new_n758), .A3(new_n776), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT52), .B1(new_n780), .B2(new_n770), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n775), .A2(new_n781), .ZN(G1337gat));
  INV_X1    g581(.A(G99gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n769), .A2(new_n715), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(KEYINPUT115), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(KEYINPUT115), .B2(new_n784), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n372), .A2(new_n783), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n766), .B2(new_n787), .ZN(G1338gat));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  OAI21_X1  g588(.A(G106gat), .B1(new_n754), .B2(new_n461), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n461), .A2(G106gat), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n789), .B(new_n790), .C1(new_n766), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n665), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n776), .B1(new_n764), .B2(new_n758), .ZN(new_n796));
  AND4_X1   g595(.A1(new_n753), .A2(new_n756), .A3(new_n758), .A4(new_n776), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n790), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT116), .B1(new_n799), .B2(KEYINPUT53), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n794), .B1(new_n778), .B2(new_n779), .ZN(new_n801));
  INV_X1    g600(.A(G106gat), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n769), .B2(new_n556), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT116), .B(KEYINPUT53), .C1(new_n801), .C2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n793), .B1(new_n800), .B2(new_n805), .ZN(G1339gat));
  NOR2_X1   g605(.A1(new_n505), .A2(new_n403), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809));
  INV_X1    g608(.A(new_n263), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n261), .A2(new_n256), .A3(new_n810), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT117), .Z(new_n812));
  AOI21_X1  g611(.A(new_n254), .B1(new_n253), .B2(new_n256), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n206), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n266), .A2(new_n208), .A3(new_n260), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(new_n665), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n645), .A2(new_n654), .A3(new_n649), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n652), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n650), .A2(new_n820), .A3(new_n651), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n661), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n817), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n652), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n661), .A4(new_n821), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n664), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n816), .B1(new_n268), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n673), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n814), .A2(new_n815), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n696), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n640), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n733), .A2(new_n665), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n809), .B1(new_n834), .B2(new_n556), .ZN(new_n835));
  OAI211_X1 g634(.A(KEYINPUT118), .B(new_n461), .C1(new_n832), .C2(new_n833), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n688), .B(new_n808), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n268), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n834), .A2(new_n505), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n462), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n268), .A2(new_n322), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(G1340gat));
  INV_X1    g642(.A(new_n841), .ZN(new_n844));
  AOI21_X1  g643(.A(G120gat), .B1(new_n844), .B2(new_n665), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n666), .A2(new_n320), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT119), .ZN(G1341gat));
  OAI21_X1  g647(.A(G127gat), .B1(new_n838), .B2(new_n695), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n844), .A2(new_n327), .A3(new_n640), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1342gat));
  NOR3_X1   g650(.A1(new_n841), .A2(G134gat), .A3(new_n673), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT56), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n838), .B2(new_n673), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n807), .A2(new_n686), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT120), .ZN(new_n857));
  INV_X1    g656(.A(new_n834), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT57), .A3(new_n556), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n834), .B2(new_n461), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n857), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n416), .B1(new_n862), .B2(new_n752), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n715), .A2(new_n403), .A3(new_n461), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n840), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n865), .A2(G141gat), .A3(new_n268), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT58), .Z(G1344gat));
  OAI21_X1  g667(.A(KEYINPUT59), .B1(new_n865), .B2(new_n666), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n666), .A2(KEYINPUT59), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n869), .A2(new_n440), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n859), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n752), .B1(new_n669), .B2(new_n674), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n832), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n556), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n874), .A2(new_n832), .A3(new_n873), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n860), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT122), .B(new_n860), .C1(new_n876), .C2(new_n877), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n666), .B(new_n857), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n871), .B1(new_n882), .B2(new_n883), .ZN(G1345gat));
  NOR2_X1   g683(.A1(new_n865), .A2(new_n695), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n886), .A2(KEYINPUT123), .ZN(new_n887));
  AOI21_X1  g686(.A(G155gat), .B1(new_n886), .B2(KEYINPUT123), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n695), .A2(new_n407), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n887), .A2(new_n888), .B1(new_n862), .B2(new_n889), .ZN(G1346gat));
  XNOR2_X1  g689(.A(KEYINPUT79), .B(G162gat), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n862), .B2(new_n696), .ZN(new_n892));
  AND4_X1   g691(.A1(new_n696), .A2(new_n840), .A3(new_n864), .A4(new_n891), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT124), .Z(G1347gat));
  NOR2_X1   g694(.A1(new_n504), .A2(new_n404), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n834), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n461), .A3(new_n372), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n752), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n372), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n835), .B2(new_n836), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n268), .A2(new_n281), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(G1348gat));
  NAND3_X1  g704(.A1(new_n900), .A2(new_n282), .A3(new_n665), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n903), .A2(new_n665), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n282), .ZN(G1349gat));
  AOI21_X1  g707(.A(new_n276), .B1(new_n903), .B2(new_n640), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n640), .A2(new_n271), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g711(.A1(new_n900), .A2(new_n270), .A3(new_n696), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n296), .B1(new_n903), .B2(new_n696), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(KEYINPUT125), .B(new_n913), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n715), .A2(new_n461), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n898), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(G197gat), .B1(new_n925), .B2(new_n752), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n897), .A2(new_n715), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n928), .B1(new_n880), .B2(new_n881), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n752), .A2(G197gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  NOR3_X1   g730(.A1(new_n924), .A2(G204gat), .A3(new_n666), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT62), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n929), .A2(new_n665), .ZN(new_n934));
  INV_X1    g733(.A(G204gat), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(G1353gat));
  AOI211_X1 g735(.A(new_n695), .B(new_n928), .C1(new_n880), .C2(new_n881), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT63), .B1(new_n937), .B2(new_n378), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n880), .A2(new_n881), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n640), .A3(new_n927), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n941), .A3(G211gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n378), .A3(new_n640), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT126), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n938), .A2(new_n942), .A3(new_n944), .ZN(G1354gat));
  AOI21_X1  g744(.A(G218gat), .B1(new_n925), .B2(new_n696), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n673), .A2(new_n379), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT127), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n929), .B2(new_n948), .ZN(G1355gat));
endmodule


