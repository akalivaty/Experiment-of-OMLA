//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n461), .A2(KEYINPUT64), .A3(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT64), .B1(new_n461), .B2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G101), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G137), .A3(new_n461), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n467), .B1(new_n474), .B2(G2105), .ZN(G160));
  AOI21_X1  g050(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT65), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT66), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n465), .A2(new_n461), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n478), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT67), .Z(G162));
  AND2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n461), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(G114), .B2(new_n461), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G62), .ZN(new_n504));
  NAND2_X1  g079(.A1(G75), .A2(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n506), .A2(KEYINPUT68), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(new_n500), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n501), .A2(new_n502), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n512), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(G88), .B1(new_n513), .B2(G50), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n506), .B2(KEYINPUT68), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n507), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND2_X1  g092(.A1(new_n509), .A2(new_n510), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n501), .B2(new_n502), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n520), .A2(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n500), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n513), .A2(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n503), .A2(new_n518), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n511), .A2(G81), .B1(new_n513), .B2(G43), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n500), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  NAND4_X1  g114(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  INV_X1    g118(.A(G78), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT71), .B1(new_n544), .B2(new_n512), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n546), .A2(G78), .A3(G543), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n503), .A2(G65), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n500), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n550), .B1(new_n549), .B2(new_n548), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(KEYINPUT70), .B2(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n513), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n554), .A2(new_n555), .B1(new_n511), .B2(G91), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n513), .B(new_n553), .C1(KEYINPUT70), .C2(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n551), .A2(new_n556), .A3(new_n557), .ZN(G299));
  XOR2_X1   g133(.A(G171), .B(KEYINPUT73), .Z(G301));
  INV_X1    g134(.A(G168), .ZN(G286));
  OAI21_X1  g135(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT74), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n511), .A2(G87), .B1(new_n513), .B2(G49), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(G288));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  INV_X1    g140(.A(G86), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n531), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n511), .A2(KEYINPUT75), .A3(G86), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(G48), .A2(G543), .ZN(new_n570));
  AND2_X1   g145(.A1(KEYINPUT6), .A2(G651), .ZN(new_n571));
  NOR2_X1   g146(.A1(KEYINPUT6), .A2(G651), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT76), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n575), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n501), .B2(new_n502), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n569), .A2(new_n577), .A3(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n511), .A2(G85), .B1(new_n513), .B2(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n500), .B2(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n503), .A2(new_n518), .A3(G92), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(KEYINPUT10), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n590), .A2(new_n591), .B1(G54), .B2(new_n513), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n503), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n500), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n594), .B2(new_n593), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n592), .A2(KEYINPUT78), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT78), .B1(new_n592), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n588), .B1(new_n600), .B2(new_n587), .ZN(G284));
  AOI21_X1  g176(.A(new_n588), .B1(new_n600), .B2(new_n587), .ZN(G321));
  NOR2_X1   g177(.A1(G286), .A2(new_n587), .ZN(new_n603));
  XOR2_X1   g178(.A(G299), .B(KEYINPUT79), .Z(new_n604));
  AOI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n587), .ZN(G297));
  AOI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n587), .ZN(G280));
  NOR2_X1   g181(.A1(new_n599), .A2(G559), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(G860), .B2(new_n600), .ZN(G148));
  INV_X1    g183(.A(new_n538), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(new_n587), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n607), .B2(new_n587), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g187(.A1(new_n462), .A2(new_n463), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n465), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT12), .Z(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT13), .Z(new_n616));
  INV_X1    g191(.A(G2100), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n476), .A2(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n461), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G135), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n620), .B1(new_n621), .B2(new_n622), .C1(new_n623), .C2(new_n483), .ZN(new_n624));
  INV_X1    g199(.A(G2096), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n618), .A2(new_n619), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT80), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2430), .Z(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n641), .A2(new_n642), .A3(G14), .ZN(G401));
  INV_X1    g218(.A(KEYINPUT18), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(new_n617), .ZN(new_n651));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n647), .B2(KEYINPUT18), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n625), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n658), .B2(new_n661), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n657), .A3(new_n661), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n664), .B(new_n667), .C1(new_n657), .C2(new_n666), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  MUX2_X1   g249(.A(G6), .B(G305), .S(G16), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT84), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT32), .B(G1981), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n682), .A2(G23), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G288), .B2(G16), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT33), .ZN(new_n685));
  INV_X1    g260(.A(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(G16), .A2(G22), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G166), .B2(G16), .ZN(new_n689));
  INV_X1    g264(.A(G1971), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n680), .A2(new_n681), .A3(new_n687), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT83), .B(KEYINPUT34), .Z(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(G25), .A2(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n476), .A2(G119), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n461), .A2(G107), .ZN(new_n698));
  OAI21_X1  g273(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n699));
  INV_X1    g274(.A(G131), .ZN(new_n700));
  OAI221_X1 g275(.A(new_n697), .B1(new_n698), .B2(new_n699), .C1(new_n700), .C2(new_n483), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT82), .Z(new_n702));
  AOI21_X1  g277(.A(new_n696), .B1(new_n702), .B2(G29), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n703), .A2(new_n705), .ZN(new_n707));
  MUX2_X1   g282(.A(G24), .B(G290), .S(G16), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1986), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n694), .A2(new_n695), .A3(new_n706), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(KEYINPUT87), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n712), .A2(KEYINPUT86), .A3(KEYINPUT36), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n711), .B2(KEYINPUT87), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(G33), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT25), .Z(new_n719));
  INV_X1    g294(.A(G139), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n483), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(new_n461), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n721), .B1(KEYINPUT89), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(KEYINPUT89), .B2(new_n723), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n717), .B1(new_n725), .B2(G29), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G2072), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT90), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n716), .A2(G32), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n484), .A2(G141), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n613), .A2(G105), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n476), .A2(G129), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT26), .Z(new_n735));
  NAND4_X1  g310(.A1(new_n731), .A2(new_n732), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n730), .B1(new_n737), .B2(new_n716), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT27), .B(G1996), .Z(new_n739));
  OAI21_X1  g314(.A(new_n716), .B1(KEYINPUT24), .B2(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(KEYINPUT24), .B2(G34), .ZN(new_n741));
  INV_X1    g316(.A(G160), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G29), .ZN(new_n743));
  INV_X1    g318(.A(G2084), .ZN(new_n744));
  OAI22_X1  g319(.A1(new_n738), .A2(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n727), .B2(G2072), .ZN(new_n746));
  AOI21_X1  g321(.A(KEYINPUT91), .B1(new_n729), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n682), .A2(G19), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n538), .B2(new_n682), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT88), .Z(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G1341), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(G1341), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n600), .A2(new_n682), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G4), .B2(new_n682), .ZN(new_n754));
  INV_X1    g329(.A(G1348), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n747), .A2(new_n751), .A3(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n738), .A2(new_n739), .B1(new_n743), .B2(new_n744), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n682), .A2(G5), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G171), .B2(new_n682), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT93), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n758), .B1(new_n761), .B2(G1961), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT94), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n716), .A2(G26), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT28), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n476), .A2(G128), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n461), .A2(G116), .ZN(new_n767));
  OAI21_X1  g342(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n768));
  INV_X1    g343(.A(G140), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n766), .B1(new_n767), .B2(new_n768), .C1(new_n769), .C2(new_n483), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n765), .B1(new_n770), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2067), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  NAND2_X1  g348(.A1(G164), .A2(G29), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G27), .B2(G29), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n772), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n773), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n761), .A2(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n682), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1956), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n682), .A2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G168), .B2(new_n682), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n784), .A2(G1966), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(G1966), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT31), .B(G11), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT92), .B(G28), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n788), .B2(KEYINPUT30), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(KEYINPUT30), .B2(new_n788), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n787), .B(new_n790), .C1(new_n624), .C2(new_n716), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n785), .A2(new_n786), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n777), .A2(new_n778), .A3(new_n782), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n716), .A2(G35), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT95), .Z(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G162), .B2(new_n716), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT29), .B(G2090), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AOI211_X1 g373(.A(new_n793), .B(new_n798), .C1(new_n755), .C2(new_n754), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n729), .A2(KEYINPUT91), .A3(new_n746), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n757), .A2(new_n763), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT86), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n711), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n713), .A2(new_n715), .A3(new_n803), .ZN(G311));
  NAND3_X1  g379(.A1(new_n713), .A2(new_n715), .A3(new_n803), .ZN(G150));
  AOI22_X1  g380(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n500), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n807), .A2(KEYINPUT96), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT98), .B(G93), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT97), .B(G55), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n511), .A2(new_n809), .B1(new_n513), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n807), .B2(KEYINPUT96), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G860), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT37), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n600), .A2(G559), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT38), .Z(new_n818));
  INV_X1    g393(.A(new_n813), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n538), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n813), .A2(new_n536), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT99), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n820), .A2(new_n824), .A3(new_n821), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n818), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n814), .B1(new_n828), .B2(KEYINPUT39), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n816), .B1(new_n829), .B2(new_n830), .ZN(G145));
  INV_X1    g406(.A(KEYINPUT104), .ZN(new_n832));
  XNOR2_X1  g407(.A(G160), .B(KEYINPUT100), .ZN(new_n833));
  XNOR2_X1  g408(.A(G162), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n624), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n498), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G114), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n495), .B1(new_n838), .B2(G2105), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G126), .B2(new_n476), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n840), .A2(KEYINPUT101), .A3(new_n493), .A4(new_n492), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n770), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n725), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n737), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n476), .A2(G130), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT102), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n484), .A2(G142), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n461), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n615), .ZN(new_n852));
  INV_X1    g427(.A(new_n702), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n835), .B1(new_n845), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n845), .B2(new_n854), .ZN(new_n856));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n854), .A2(KEYINPUT103), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n859), .A2(new_n845), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n845), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n835), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n832), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n863), .A2(new_n856), .A3(KEYINPUT104), .A4(new_n857), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g443(.A(G305), .B(KEYINPUT107), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G303), .ZN(new_n870));
  XNOR2_X1  g445(.A(G288), .B(G290), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT42), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n826), .A2(KEYINPUT105), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n823), .A2(new_n875), .A3(new_n825), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n607), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n607), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n592), .A2(new_n596), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G299), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n879), .A2(new_n880), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n873), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n891), .A2(KEYINPUT109), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n885), .A2(new_n873), .A3(new_n890), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n893), .A2(KEYINPUT108), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(KEYINPUT108), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(KEYINPUT109), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n892), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G868), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(G868), .B2(new_n813), .ZN(G295));
  OAI21_X1  g474(.A(new_n898), .B1(G868), .B2(new_n813), .ZN(G331));
  NOR2_X1   g475(.A1(G301), .A2(G286), .ZN(new_n901));
  NOR2_X1   g476(.A1(G168), .A2(G171), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n826), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n823), .B(new_n825), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n826), .A2(KEYINPUT110), .A3(new_n903), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n883), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT111), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n904), .A2(new_n906), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n909), .A2(new_n910), .B1(new_n912), .B2(new_n889), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n913), .A3(new_n872), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n914), .A2(new_n857), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(new_n872), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT43), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n912), .A2(new_n883), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n883), .A2(new_n888), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n886), .B2(new_n883), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n907), .A2(new_n908), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(new_n923), .B2(KEYINPUT112), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(KEYINPUT112), .B2(new_n923), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n917), .ZN(new_n926));
  AND4_X1   g501(.A1(KEYINPUT43), .A2(new_n926), .A3(new_n857), .A4(new_n914), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n919), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n915), .B2(new_n918), .ZN(new_n931));
  AND4_X1   g506(.A1(new_n930), .A2(new_n926), .A3(new_n857), .A4(new_n914), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n933), .ZN(G397));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n842), .B2(G1384), .ZN(new_n936));
  OAI21_X1  g511(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n937), .A2(G40), .A3(new_n464), .A4(new_n466), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G1996), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n736), .B(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G2067), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n770), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT113), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n853), .A2(new_n705), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n702), .A2(new_n704), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n939), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(G290), .B(G1986), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n939), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(G299), .B(KEYINPUT57), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n498), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n954), .B1(new_n498), .B2(new_n955), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n957), .A2(new_n958), .A3(new_n938), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(G1956), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n498), .A2(new_n955), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n938), .B1(new_n961), .B2(new_n935), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n935), .A2(G1384), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n837), .A2(new_n841), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(KEYINPUT56), .B(G2072), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n953), .A2(new_n960), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n959), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n961), .A2(new_n938), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n968), .A2(new_n755), .B1(new_n942), .B2(new_n969), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n967), .A2(new_n599), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n960), .A2(new_n966), .ZN(new_n972));
  XOR2_X1   g547(.A(G299), .B(KEYINPUT57), .Z(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n962), .A2(new_n964), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n940), .ZN(new_n977));
  INV_X1    g552(.A(new_n969), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT124), .B(KEYINPUT58), .Z(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(G1341), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n609), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT59), .Z(new_n983));
  INV_X1    g558(.A(KEYINPUT61), .ZN(new_n984));
  OR3_X1    g559(.A1(new_n974), .A2(new_n967), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n974), .B2(new_n967), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n970), .A2(new_n600), .A3(KEYINPUT60), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(KEYINPUT60), .B2(new_n970), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n970), .A2(KEYINPUT60), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n599), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n975), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n498), .A2(new_n963), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n962), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(G1966), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n995), .A2(KEYINPUT120), .B1(new_n744), .B2(new_n959), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT120), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n994), .B2(G1966), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(G168), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G8), .ZN(new_n1000));
  AOI21_X1  g575(.A(G168), .B1(new_n996), .B2(new_n998), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT51), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n1003), .A3(G8), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT53), .B1(new_n976), .B2(new_n773), .ZN(new_n1006));
  INV_X1    g581(.A(G1961), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n968), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n773), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n474), .A2(KEYINPUT125), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n461), .B1(new_n474), .B2(KEYINPUT125), .ZN(new_n1011));
  AOI211_X1 g586(.A(new_n467), .B(new_n1009), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(new_n936), .A3(new_n964), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n528), .B(new_n532), .C1(new_n1008), .C2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n994), .A2(KEYINPUT53), .A3(new_n773), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1008), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G301), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT54), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1008), .A2(G301), .A3(new_n1013), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n992), .A2(new_n1005), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1020), .ZN(new_n1026));
  NOR2_X1   g601(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1028));
  AND2_X1   g603(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1005), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1025), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n978), .B(G8), .C1(new_n686), .C2(G288), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT52), .B1(G288), .B2(new_n686), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(KEYINPUT52), .B2(new_n1033), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n978), .A2(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n511), .A2(G86), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n577), .A2(new_n582), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G1981), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT116), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1044), .A3(G1981), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1981), .B1(new_n574), .B2(new_n576), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT75), .B1(new_n511), .B2(G86), .ZN(new_n1048));
  AND4_X1   g623(.A1(KEYINPUT75), .A2(new_n503), .A3(new_n518), .A4(G86), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1047), .B(new_n582), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT115), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n569), .A2(new_n1052), .A3(new_n582), .A4(new_n1047), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1046), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1039), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1043), .A2(new_n1045), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT117), .B1(new_n1058), .B2(KEYINPUT49), .ZN(new_n1059));
  AND4_X1   g634(.A1(KEYINPUT117), .A2(new_n1046), .A3(new_n1054), .A4(KEYINPUT49), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT118), .B(new_n1057), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1038), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n507), .B2(new_n515), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT55), .B(G8), .C1(new_n507), .C2(new_n515), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1971), .B1(new_n962), .B2(new_n964), .ZN(new_n1071));
  NOR4_X1   g646(.A1(new_n957), .A2(new_n958), .A3(G2090), .A4(new_n938), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1070), .B(G8), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n962), .A2(new_n964), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n690), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n958), .A2(new_n938), .ZN(new_n1078));
  INV_X1    g653(.A(G2090), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n956), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(KEYINPUT114), .A3(G8), .A4(new_n1070), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1077), .A2(KEYINPUT119), .A3(new_n1080), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1085), .A3(G8), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1070), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1075), .A2(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1065), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1032), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1065), .A2(new_n1075), .A3(new_n1082), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G288), .A2(G1976), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1092), .A2(new_n1093), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1091), .B1(new_n1094), .B2(new_n1039), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1096));
  NAND2_X1  g671(.A1(G168), .A2(G8), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n996), .B2(new_n998), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1081), .A2(G8), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(new_n1087), .ZN(new_n1101));
  AND4_X1   g676(.A1(new_n1065), .A2(new_n1096), .A3(new_n1098), .A4(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1092), .A2(new_n1088), .A3(new_n1037), .A4(new_n1098), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1065), .A2(KEYINPUT121), .A3(new_n1088), .A4(new_n1098), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1099), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1102), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1105), .A2(new_n1106), .A3(KEYINPUT122), .A4(new_n1099), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1095), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1090), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g688(.A(KEYINPUT123), .B(new_n1095), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n952), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n939), .ZN(new_n1116));
  OR3_X1    g691(.A1(new_n1116), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT46), .B1(new_n1116), .B2(G1996), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n943), .A2(new_n737), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1117), .A2(new_n1118), .B1(new_n939), .B2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n1120), .B(KEYINPUT47), .Z(new_n1121));
  NOR3_X1   g696(.A1(new_n1116), .A2(G1986), .A3(G290), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT48), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n950), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n946), .A2(new_n947), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(G2067), .B2(new_n770), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(KEYINPUT127), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(new_n1116), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(KEYINPUT127), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1115), .A2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g706(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1133));
  OAI211_X1 g707(.A(new_n867), .B(new_n1133), .C1(new_n931), .C2(new_n932), .ZN(G225));
  INV_X1    g708(.A(G225), .ZN(G308));
endmodule


