//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1379, new_n1380, new_n1381, new_n1382;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OR2_X1    g0012(.A1(KEYINPUT64), .A2(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(KEYINPUT64), .A2(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n203), .A2(G50), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n201), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n218), .B2(new_n219), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT17), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n252), .B1(new_n206), .B2(G20), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n216), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n254), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n253), .A2(new_n257), .B1(new_n258), .B2(new_n252), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G58), .A2(G68), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT76), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(KEYINPUT76), .A2(G58), .A3(G68), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(new_n203), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n264), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n267), .A2(new_n268), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT7), .ZN(new_n270));
  OAI21_X1  g0070(.A(G68), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n215), .A2(new_n272), .A3(KEYINPUT7), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n266), .B(KEYINPUT16), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n255), .A2(new_n216), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT7), .B1(new_n215), .B2(new_n272), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n269), .A2(new_n270), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(G68), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT16), .B1(new_n279), .B2(new_n266), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n259), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(G226), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G1698), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n285), .B1(G223), .B2(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G87), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(new_n283), .A3(G274), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n292), .B1(new_n221), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g0096(.A(KEYINPUT79), .B(G190), .Z(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n296), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n251), .B1(new_n281), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n279), .A2(new_n266), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT16), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(new_n275), .A3(new_n274), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n288), .A2(new_n295), .A3(new_n297), .ZN(new_n307));
  INV_X1    g0107(.A(new_n288), .ZN(new_n308));
  INV_X1    g0108(.A(new_n295), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n307), .B1(G200), .B2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n306), .A2(new_n311), .A3(KEYINPUT17), .A4(new_n259), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n302), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n281), .A2(KEYINPUT77), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT77), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n259), .C1(new_n276), .C2(new_n280), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n296), .A2(G179), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n296), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n314), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT18), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(KEYINPUT78), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n313), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT80), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT78), .B(KEYINPUT18), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n314), .A2(new_n316), .A3(new_n319), .A4(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n320), .A2(new_n322), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n302), .A2(new_n312), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n326), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT80), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G1698), .ZN(new_n333));
  OAI211_X1 g0133(.A(G222), .B(new_n333), .C1(new_n267), .C2(new_n268), .ZN(new_n334));
  OAI211_X1 g0134(.A(G223), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n335));
  INV_X1    g0135(.A(G77), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n334), .B(new_n335), .C1(new_n336), .C2(new_n272), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT68), .ZN(new_n340));
  INV_X1    g0140(.A(new_n294), .ZN(new_n341));
  INV_X1    g0141(.A(G274), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n217), .B2(new_n282), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n341), .A2(G226), .B1(new_n343), .B2(new_n291), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n340), .B1(new_n339), .B2(new_n344), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n318), .ZN(new_n349));
  INV_X1    g0149(.A(new_n347), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n345), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n354));
  INV_X1    g0154(.A(G150), .ZN(new_n355));
  INV_X1    g0155(.A(new_n265), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n213), .A2(G33), .A3(new_n214), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n354), .B1(new_n355), .B2(new_n356), .C1(new_n357), .C2(new_n252), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n275), .ZN(new_n359));
  INV_X1    g0159(.A(new_n275), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n206), .A2(G20), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n360), .A2(G50), .A3(new_n254), .A4(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G50), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n258), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT69), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(G50), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n364), .B(KEYINPUT69), .C1(new_n256), .C2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n359), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n349), .A2(new_n353), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(G190), .B1(new_n346), .B2(new_n347), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(KEYINPUT72), .B(G190), .C1(new_n346), .C2(new_n347), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n346), .A2(new_n347), .A3(new_n300), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT10), .B1(new_n376), .B2(KEYINPUT73), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n369), .A2(KEYINPUT9), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT9), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n359), .B(new_n379), .C1(new_n368), .C2(new_n365), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n348), .A2(G200), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n375), .A2(new_n377), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n377), .B1(new_n375), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n370), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n257), .A2(G68), .A3(new_n361), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT12), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n258), .B2(new_n202), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n254), .A2(KEYINPUT12), .A3(G68), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n265), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n357), .B2(new_n336), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n391), .A2(KEYINPUT11), .A3(new_n275), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT11), .B1(new_n391), .B2(new_n275), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n389), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n284), .A2(new_n333), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n221), .A2(G1698), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n398), .C1(new_n267), .C2(new_n268), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G97), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n338), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n283), .A2(G238), .A3(new_n293), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n292), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n396), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n283), .B1(new_n399), .B2(new_n400), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n292), .A2(new_n403), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT13), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n395), .B(G169), .C1(new_n405), .C2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n402), .A2(new_n404), .A3(new_n396), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT13), .B1(new_n406), .B2(new_n407), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G179), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n411), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n395), .B1(new_n414), .B2(G169), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT74), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n405), .A2(new_n408), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT14), .B1(new_n417), .B2(new_n318), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT74), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(new_n412), .A4(new_n409), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n394), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G190), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n394), .B1(new_n422), .B2(new_n414), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n417), .A2(new_n300), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n421), .A2(KEYINPUT75), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n384), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n215), .A2(G77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n428), .B1(new_n357), .B2(new_n429), .C1(new_n356), .C2(new_n252), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n275), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n336), .B1(new_n206), .B2(G20), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n257), .A2(new_n432), .B1(new_n336), .B2(new_n258), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT70), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n431), .A2(KEYINPUT70), .A3(new_n433), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n272), .A2(G232), .A3(new_n333), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n272), .A2(G238), .A3(G1698), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(new_n222), .C2(new_n272), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n338), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n341), .A2(G244), .B1(new_n343), .B2(new_n291), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n352), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n318), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n438), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(G200), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(G190), .A3(new_n443), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n436), .A2(new_n437), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n447), .A2(KEYINPUT71), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT71), .B1(new_n447), .B2(new_n450), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT75), .B1(new_n421), .B2(new_n425), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n332), .A2(new_n427), .A3(KEYINPUT81), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT81), .ZN(new_n457));
  INV_X1    g0257(.A(new_n370), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT72), .B1(new_n351), .B2(G190), .ZN(new_n459));
  INV_X1    g0259(.A(new_n374), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n381), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n377), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n375), .A2(new_n377), .A3(new_n381), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n416), .A2(new_n420), .ZN(new_n466));
  INV_X1    g0266(.A(new_n394), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT75), .ZN(new_n469));
  INV_X1    g0269(.A(new_n425), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n465), .A2(new_n471), .A3(new_n454), .A4(new_n453), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n327), .A2(new_n331), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n457), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n456), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT64), .A2(G20), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT64), .A2(G20), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(new_n272), .A3(G87), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT22), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n479), .A2(new_n272), .A3(KEYINPUT22), .A4(G87), .ZN(new_n483));
  OR2_X1    g0283(.A1(KEYINPUT23), .A2(G107), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n213), .B2(new_n214), .ZN(new_n485));
  AOI22_X1  g0285(.A1(KEYINPUT89), .A2(KEYINPUT24), .B1(KEYINPUT23), .B2(G107), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n486), .B1(G20), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n482), .A2(new_n483), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT89), .A2(KEYINPUT24), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n360), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n491), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n482), .A2(new_n489), .A3(new_n493), .A4(new_n483), .ZN(new_n494));
  OR3_X1    g0294(.A1(new_n254), .A2(KEYINPUT25), .A3(G107), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT25), .B1(new_n254), .B2(G107), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n206), .A2(G33), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n254), .A2(new_n497), .A3(new_n216), .A4(new_n255), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n495), .B(new_n496), .C1(new_n222), .C2(new_n498), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n499), .A2(KEYINPUT90), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(KEYINPUT90), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n492), .A2(new_n494), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G257), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(new_n333), .C1(new_n267), .C2(new_n268), .ZN(new_n504));
  AND2_X1   g0304(.A1(KEYINPUT91), .A2(G294), .ZN(new_n505));
  NOR2_X1   g0305(.A1(KEYINPUT91), .A2(G294), .ZN(new_n506));
  OAI21_X1  g0306(.A(G33), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT92), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n283), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT92), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n206), .A2(G45), .ZN(new_n513));
  OR2_X1    g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n343), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n516), .A2(new_n223), .A3(new_n338), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AND4_X1   g0319(.A1(new_n422), .A2(new_n512), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n518), .B1(new_n510), .B2(new_n511), .ZN(new_n521));
  AOI21_X1  g0321(.A(G200), .B1(new_n521), .B2(new_n517), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n502), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT93), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n502), .B(KEYINPUT93), .C1(new_n520), .C2(new_n522), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g0327(.A(KEYINPUT5), .B(G41), .ZN(new_n528));
  INV_X1    g0328(.A(new_n513), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(G257), .A3(new_n283), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n517), .ZN(new_n532));
  OAI211_X1 g0332(.A(G244), .B(new_n333), .C1(new_n267), .C2(new_n268), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n272), .A2(KEYINPUT4), .A3(G244), .A4(new_n333), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n535), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n532), .B1(new_n338), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n352), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n267), .A2(new_n268), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n270), .B1(new_n479), .B2(new_n542), .ZN(new_n543));
  NOR4_X1   g0343(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT7), .A4(G20), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n543), .A2(new_n544), .A3(new_n222), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n222), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  XNOR2_X1  g0346(.A(G97), .B(G107), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n549), .A2(new_n479), .B1(new_n336), .B2(new_n356), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n275), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n254), .A2(G97), .ZN(new_n552));
  INV_X1    g0352(.A(new_n498), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(G97), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n541), .B(new_n555), .C1(G169), .C2(new_n540), .ZN(new_n556));
  INV_X1    g0356(.A(new_n554), .ZN(new_n557));
  INV_X1    g0357(.A(new_n546), .ZN(new_n558));
  AND2_X1   g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  NOR2_X1   g0359(.A1(G97), .A2(G107), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n548), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(new_n215), .B1(G77), .B2(new_n265), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n277), .A2(new_n278), .A3(G107), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n557), .B1(new_n565), .B2(new_n275), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n539), .A2(new_n338), .ZN(new_n567));
  INV_X1    g0367(.A(new_n532), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(G190), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n540), .A2(G200), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n566), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR4_X1   g0372(.A1(KEYINPUT82), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G87), .A2(G97), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n222), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n400), .A2(new_n577), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n573), .A2(new_n576), .B1(new_n215), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G97), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n357), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n479), .A2(new_n272), .A3(G68), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT83), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n579), .A2(new_n581), .A3(new_n585), .A4(new_n582), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n275), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n498), .A2(new_n429), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n429), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n254), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n587), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G244), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n594));
  OAI211_X1 g0394(.A(G238), .B(new_n333), .C1(new_n267), .C2(new_n268), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G116), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n338), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n283), .A2(G274), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n513), .A2(G250), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n599), .A2(new_n513), .B1(new_n338), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n318), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n338), .B2(new_n597), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n352), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n593), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n598), .A2(new_n602), .A3(new_n422), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n605), .B2(G200), .ZN(new_n610));
  INV_X1    g0410(.A(G87), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n498), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n610), .A2(new_n587), .A3(new_n592), .A4(new_n613), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n556), .A2(new_n572), .A3(new_n608), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n490), .A2(new_n491), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n275), .A3(new_n494), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n500), .A2(new_n501), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n512), .A2(new_n517), .A3(new_n519), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n318), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n521), .A2(new_n352), .A3(new_n517), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n527), .A2(new_n615), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(G33), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G97), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n213), .A2(new_n626), .A3(new_n214), .A4(new_n537), .ZN(new_n627));
  INV_X1    g0427(.A(G116), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n255), .A2(new_n216), .B1(G20), .B2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n627), .A2(KEYINPUT20), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT20), .B1(new_n627), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n258), .A2(new_n628), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n498), .B2(new_n628), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT85), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n627), .A2(new_n629), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n627), .A2(KEYINPUT20), .A3(new_n629), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT85), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n318), .B1(new_n635), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT86), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(KEYINPUT21), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n338), .B1(new_n529), .B2(new_n528), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n647), .A2(G270), .B1(new_n343), .B2(new_n516), .ZN(new_n648));
  OAI211_X1 g0448(.A(G264), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n649));
  OAI211_X1 g0449(.A(G257), .B(new_n333), .C1(new_n267), .C2(new_n268), .ZN(new_n650));
  INV_X1    g0450(.A(G303), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n649), .B(new_n650), .C1(new_n651), .C2(new_n272), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n338), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n648), .A2(new_n653), .A3(KEYINPUT84), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT84), .B1(new_n648), .B2(new_n653), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n643), .A2(new_n646), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n648), .A2(new_n653), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n352), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n632), .A2(KEYINPUT85), .A3(new_n634), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n640), .A2(new_n641), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n646), .B1(new_n643), .B2(new_n656), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n298), .B1(new_n654), .B2(new_n655), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT84), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n658), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n648), .A2(new_n653), .A3(KEYINPUT84), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G200), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n640), .B(KEYINPUT85), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n666), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT87), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n666), .A2(new_n670), .A3(new_n671), .A4(KEYINPUT87), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n665), .A2(new_n676), .A3(KEYINPUT88), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT88), .B1(new_n665), .B2(new_n676), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n624), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n476), .A2(new_n679), .ZN(G372));
  NOR2_X1   g0480(.A1(new_n447), .A2(new_n425), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n329), .B1(new_n421), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n281), .A2(new_n319), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT18), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n281), .A2(new_n321), .A3(new_n319), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n463), .A2(new_n464), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n458), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(G169), .B1(new_n660), .B2(new_n661), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n668), .A2(new_n669), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n645), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(new_n662), .A3(new_n623), .A4(new_n657), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n527), .A2(new_n615), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n360), .B1(new_n583), .B2(KEYINPUT83), .ZN(new_n696));
  AOI211_X1 g0496(.A(new_n591), .B(new_n612), .C1(new_n696), .C2(new_n586), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n697), .A2(new_n610), .B1(new_n593), .B2(new_n607), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n567), .A2(new_n568), .A3(new_n352), .ZN(new_n699));
  AOI21_X1  g0499(.A(G169), .B1(new_n567), .B2(new_n568), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n699), .A2(new_n566), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT26), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n608), .A3(KEYINPUT26), .A4(new_n614), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n608), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n695), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n690), .B1(new_n476), .B2(new_n706), .ZN(G369));
  NAND3_X1  g0507(.A1(new_n479), .A2(new_n206), .A3(G13), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT27), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT27), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G213), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G343), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n671), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n677), .B2(new_n678), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n665), .A2(new_n716), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT94), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n722), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n623), .A2(new_n713), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n525), .A2(new_n526), .B1(new_n619), .B2(new_n713), .ZN(new_n728));
  INV_X1    g0528(.A(new_n623), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n730), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n665), .A2(new_n713), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT95), .B1(new_n735), .B2(new_n727), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT95), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n737), .B(new_n726), .C1(new_n733), .C2(new_n734), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n732), .B1(new_n736), .B2(new_n738), .ZN(G399));
  INV_X1    g0539(.A(KEYINPUT96), .ZN(new_n740));
  INV_X1    g0540(.A(new_n210), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(G41), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n210), .A2(KEYINPUT96), .A3(new_n289), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n573), .A2(new_n576), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n628), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(G1), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n219), .B2(new_n744), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  INV_X1    g0550(.A(new_n608), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT26), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n588), .B(new_n591), .C1(new_n696), .C2(new_n586), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n604), .A2(new_n606), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n614), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n752), .B1(new_n755), .B2(new_n556), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n751), .B1(new_n756), .B2(new_n703), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n527), .A2(new_n615), .A3(new_n694), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n713), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT29), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n569), .A2(new_n300), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n540), .A2(new_n422), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n555), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(KEYINPUT99), .B1(new_n701), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT99), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n572), .A2(new_n556), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n768), .A2(new_n527), .A3(new_n698), .A4(new_n694), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT98), .ZN(new_n770));
  AND3_X1   g0570(.A1(new_n593), .A2(new_n607), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n593), .B2(new_n607), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n756), .B2(new_n703), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n713), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n761), .B1(new_n760), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G330), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n624), .B(new_n714), .C1(new_n677), .C2(new_n678), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n659), .A2(new_n521), .A3(new_n540), .A4(new_n605), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT30), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(KEYINPUT97), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT97), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n779), .A2(new_n783), .A3(new_n780), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n658), .A2(new_n603), .A3(new_n352), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n785), .A2(KEYINPUT30), .A3(new_n521), .A4(new_n540), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n540), .A2(G179), .A3(new_n605), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n656), .A3(new_n620), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n782), .A2(new_n784), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(KEYINPUT31), .B1(new_n789), .B2(new_n713), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n713), .A2(KEYINPUT31), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n788), .A2(new_n786), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(new_n792), .B2(new_n781), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n777), .B1(new_n778), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n776), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n750), .B1(new_n796), .B2(G1), .ZN(G364));
  INV_X1    g0597(.A(new_n724), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n777), .ZN(new_n799));
  INV_X1    g0599(.A(new_n744), .ZN(new_n800));
  INV_X1    g0600(.A(G13), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n215), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G45), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G1), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n799), .A2(new_n725), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n210), .A2(new_n272), .ZN(new_n808));
  INV_X1    g0608(.A(G355), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n808), .A2(new_n809), .B1(G116), .B2(new_n210), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n741), .A2(new_n272), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n219), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(new_n290), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n246), .A2(G45), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n810), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G13), .A2(G33), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G20), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n216), .B1(G20), .B2(new_n318), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n805), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n215), .A2(new_n422), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT100), .ZN(new_n825));
  NOR2_X1   g0625(.A1(G179), .A2(G200), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G159), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT32), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n479), .A2(new_n352), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G200), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(G190), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n300), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(G190), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G68), .A2(new_n833), .B1(new_n835), .B2(G77), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n834), .A2(new_n297), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n836), .B1(new_n201), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n300), .A2(G179), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n825), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n222), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n841), .A2(new_n207), .A3(new_n422), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n542), .B1(new_n845), .B2(G87), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n215), .B1(new_n422), .B2(new_n827), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n832), .A2(new_n297), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n846), .B1(new_n580), .B2(new_n848), .C1(new_n850), .C2(new_n363), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n830), .A2(new_n839), .A3(new_n844), .A4(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n854));
  INV_X1    g0654(.A(new_n828), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n855), .A2(KEYINPUT102), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(KEYINPUT102), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(G329), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n849), .A2(G326), .ZN(new_n860));
  INV_X1    g0660(.A(new_n835), .ZN(new_n861));
  INV_X1    g0661(.A(G311), .ZN(new_n862));
  INV_X1    g0662(.A(new_n833), .ZN(new_n863));
  XOR2_X1   g0663(.A(KEYINPUT103), .B(KEYINPUT33), .Z(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(G317), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n860), .B1(new_n861), .B2(new_n862), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n837), .A2(G322), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n272), .B1(new_n845), .B2(G303), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n505), .A2(new_n506), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n848), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G283), .B2(new_n842), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n859), .A2(new_n867), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n854), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n823), .B1(new_n875), .B2(new_n820), .ZN(new_n876));
  INV_X1    g0676(.A(new_n819), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n724), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n807), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(G396));
  AOI22_X1  g0680(.A1(G50), .A2(new_n845), .B1(new_n847), .B2(G58), .ZN(new_n881));
  AOI22_X1  g0681(.A1(G143), .A2(new_n837), .B1(new_n835), .B2(G159), .ZN(new_n882));
  INV_X1    g0682(.A(G137), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n882), .B1(new_n883), .B2(new_n850), .C1(new_n355), .C2(new_n863), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT34), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n881), .B1(new_n202), .B2(new_n843), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n542), .B1(new_n858), .B2(G132), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT106), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n886), .B(new_n888), .C1(new_n885), .C2(new_n884), .ZN(new_n889));
  AOI22_X1  g0689(.A1(G283), .A2(new_n833), .B1(new_n849), .B2(G303), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n628), .B2(new_n861), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT104), .Z(new_n892));
  INV_X1    g0692(.A(new_n845), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n542), .B1(new_n848), .B2(new_n580), .C1(new_n222), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n843), .A2(new_n611), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n894), .B(new_n895), .C1(G294), .C2(new_n837), .ZN(new_n896));
  INV_X1    g0696(.A(new_n858), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n892), .B(new_n896), .C1(new_n862), .C2(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT105), .Z(new_n899));
  OAI21_X1  g0699(.A(new_n820), .B1(new_n889), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n820), .A2(new_n817), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n806), .B1(new_n336), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n438), .A2(new_n713), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n450), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n904), .A2(new_n447), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n447), .A2(new_n713), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n900), .B(new_n902), .C1(new_n818), .C2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n907), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n759), .B(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n795), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n805), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n911), .A2(new_n912), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n908), .B1(new_n914), .B2(new_n915), .ZN(G384));
  NOR2_X1   g0716(.A1(new_n802), .A2(new_n206), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n714), .A2(new_n394), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n468), .B2(new_n470), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n421), .A2(new_n425), .A3(new_n918), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n907), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n789), .A2(KEYINPUT31), .A3(new_n713), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(new_n790), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n778), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT38), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n479), .A2(new_n542), .A3(new_n270), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n927), .B(G68), .C1(new_n270), .C2(new_n269), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT16), .B1(new_n928), .B2(new_n266), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n259), .B1(new_n276), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n711), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n323), .B2(new_n326), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n314), .A2(new_n316), .A3(new_n931), .ZN(new_n934));
  INV_X1    g0734(.A(new_n281), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT37), .B1(new_n935), .B2(new_n311), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n320), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n306), .A2(new_n311), .A3(new_n259), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n930), .A2(new_n319), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n932), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT37), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n926), .B1(new_n933), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n932), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n330), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(KEYINPUT38), .A3(new_n942), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT40), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n925), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  INV_X1    g0750(.A(new_n934), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n938), .A2(new_n683), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT37), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n937), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n951), .B1(new_n686), .B2(new_n313), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n926), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n947), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n950), .B1(new_n925), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n949), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n778), .A2(new_n924), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n475), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(G330), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n962), .B2(new_n960), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT109), .Z(new_n965));
  NOR2_X1   g0765(.A1(new_n687), .A2(new_n931), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n920), .A2(new_n921), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n907), .B(new_n714), .C1(new_n695), .C2(new_n705), .ZN(new_n968));
  INV_X1    g0768(.A(new_n906), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n944), .A2(new_n947), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT108), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT39), .ZN(new_n974));
  AOI221_X4 g0774(.A(new_n926), .B1(new_n937), .B2(new_n941), .C1(new_n330), .C2(new_n945), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT38), .B1(new_n954), .B2(new_n955), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n944), .A2(KEYINPUT39), .A3(new_n947), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n468), .A2(new_n713), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n972), .A2(new_n973), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n973), .B1(new_n972), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n475), .A2(new_n776), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n690), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n983), .B(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n917), .B1(new_n965), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n965), .B2(new_n986), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n813), .A2(G77), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n262), .A2(new_n263), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n989), .A2(new_n990), .B1(G50), .B2(new_n202), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(G1), .A3(new_n801), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT107), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT36), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n628), .B(new_n218), .C1(new_n562), .C2(KEYINPUT35), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(KEYINPUT35), .B2(new_n562), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n993), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n994), .B2(new_n996), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n988), .A2(new_n998), .ZN(G367));
  INV_X1    g0799(.A(new_n735), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n768), .B1(new_n566), .B2(new_n714), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n701), .A2(new_n713), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT42), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1001), .A2(new_n623), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n713), .B1(new_n1006), .B2(new_n556), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n1004), .B2(KEYINPUT42), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n697), .A2(new_n714), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n751), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n755), .A2(new_n1010), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1016), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1009), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1005), .A2(new_n1008), .A3(new_n1017), .A4(new_n1016), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1003), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n732), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1023), .B(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n744), .B(KEYINPUT41), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n733), .A2(new_n734), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1000), .A2(KEYINPUT111), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(G330), .A3(new_n724), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1031), .B1(new_n724), .B2(G330), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1029), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n725), .A2(new_n1030), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1036), .A2(new_n1028), .A3(new_n1032), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n735), .A2(new_n727), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n737), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n735), .A2(KEYINPUT95), .A3(new_n727), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n1041), .A3(new_n1024), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT44), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(KEYINPUT44), .A3(new_n1041), .A4(new_n1024), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1003), .B1(new_n736), .B2(new_n738), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT45), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(KEYINPUT45), .B(new_n1003), .C1(new_n736), .C2(new_n738), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n731), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n732), .A2(new_n1046), .A3(new_n1051), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1038), .A2(new_n1053), .A3(new_n796), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1027), .B1(new_n1055), .B2(new_n796), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1026), .B1(new_n1056), .B2(new_n804), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n241), .A2(new_n812), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n821), .B1(new_n210), .B2(new_n429), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n805), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n848), .A2(new_n202), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n272), .B1(new_n893), .B2(new_n201), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G50), .C2(new_n835), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n842), .A2(G77), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n883), .C2(new_n855), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G143), .A2(new_n849), .B1(new_n837), .B2(G150), .ZN(new_n1066));
  INV_X1    g0866(.A(G159), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1066), .B1(new_n1067), .B2(new_n863), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n837), .A2(G303), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n835), .A2(G283), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n862), .B2(new_n850), .C1(new_n870), .C2(new_n863), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT46), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n893), .B2(new_n628), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n845), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n542), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G107), .B2(new_n847), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT112), .B(G317), .Z(new_n1078));
  NAND2_X1  g0878(.A1(new_n828), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n842), .A2(G97), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1065), .A2(new_n1068), .B1(new_n1072), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT47), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1060), .B1(new_n1083), .B2(new_n820), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1019), .B2(new_n877), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1057), .A2(new_n1085), .ZN(G387));
  AOI21_X1  g0886(.A(new_n744), .B1(new_n1038), .B2(new_n796), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n796), .B2(new_n1038), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n747), .A2(new_n808), .B1(G107), .B2(new_n210), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n237), .A2(G45), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT113), .ZN(new_n1091));
  AOI211_X1 g0891(.A(G45), .B(new_n746), .C1(G68), .C2(G77), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n252), .A2(G50), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT50), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n812), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1089), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n805), .B1(new_n1096), .B2(new_n822), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n733), .A2(new_n877), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n1067), .A2(new_n850), .B1(new_n863), .B2(new_n252), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G68), .B2(new_n835), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n828), .A2(G150), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n272), .B1(new_n848), .B2(new_n429), .C1(new_n336), .C2(new_n893), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G50), .B2(new_n837), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1100), .A2(new_n1080), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n272), .B1(new_n828), .B2(G326), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G322), .A2(new_n849), .B1(new_n837), .B2(new_n1078), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n651), .B2(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT48), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n870), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1111), .A2(new_n845), .B1(new_n847), .B2(G283), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT49), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1105), .B1(new_n628), .B2(new_n843), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1104), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1097), .B(new_n1098), .C1(new_n820), .C2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1038), .B2(new_n804), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1088), .A2(new_n1119), .ZN(G393));
  NAND3_X1  g0920(.A1(new_n1053), .A2(new_n804), .A3(new_n1054), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n821), .B1(new_n580), .B2(new_n210), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n811), .B2(new_n249), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n806), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n820), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G311), .A2(new_n837), .B1(new_n849), .B2(G317), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT52), .Z(new_n1127));
  INV_X1    g0927(.A(G283), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n542), .B1(new_n893), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G116), .B2(new_n847), .ZN(new_n1130));
  INV_X1    g0930(.A(G294), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n861), .C1(new_n651), .C2(new_n863), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n844), .B(new_n1132), .C1(G322), .C2(new_n828), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n272), .B1(new_n893), .B2(new_n202), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G77), .B2(new_n847), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n363), .B2(new_n863), .C1(new_n252), .C2(new_n861), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n895), .B(new_n1136), .C1(G143), .C2(new_n828), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G150), .A2(new_n849), .B1(new_n837), .B2(G159), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT51), .Z(new_n1139));
  AOI22_X1  g0939(.A1(new_n1127), .A2(new_n1133), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1124), .B1(new_n1003), .B2(new_n877), .C1(new_n1125), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1055), .A2(new_n800), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1038), .A2(new_n796), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1121), .B(new_n1141), .C1(new_n1142), .C2(new_n1143), .ZN(G390));
  NAND2_X1  g0944(.A1(new_n977), .A2(new_n978), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n979), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n906), .B1(new_n759), .B2(new_n907), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n967), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n778), .A2(new_n794), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n967), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1150), .A2(G330), .A3(new_n907), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n769), .A2(new_n774), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n905), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n714), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n967), .B1(new_n1155), .B2(new_n969), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1146), .B1(new_n975), .B2(new_n976), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1156), .A2(new_n1157), .A3(KEYINPUT114), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT114), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n713), .B(new_n905), .C1(new_n769), .C2(new_n774), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1151), .B1(new_n1160), .B2(new_n906), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n979), .B1(new_n957), .B2(new_n947), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1149), .B(new_n1152), .C1(new_n1158), .C2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(KEYINPUT114), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1165), .A2(new_n1166), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n777), .B(new_n922), .C1(new_n778), .C2(new_n924), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1164), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n968), .A2(new_n969), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1151), .B1(new_n795), .B2(new_n907), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n1168), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1160), .A2(new_n906), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n777), .B(new_n909), .C1(new_n778), .C2(new_n924), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1152), .C1(new_n1175), .C2(new_n1151), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n777), .B1(new_n778), .B2(new_n924), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n475), .A2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n984), .A2(new_n1179), .A3(new_n690), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(KEYINPUT115), .B(new_n800), .C1(new_n1170), .C2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1170), .A2(new_n1181), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1149), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1168), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1186), .A2(new_n1164), .A3(new_n1180), .A4(new_n1177), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT115), .B1(new_n1187), .B2(new_n800), .ZN(new_n1188));
  OAI21_X1  g0988(.A(KEYINPUT116), .B1(new_n1184), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n800), .B1(new_n1170), .B2(new_n1181), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT115), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT116), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n1183), .A4(new_n1182), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1189), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1186), .A2(new_n804), .A3(new_n1164), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1145), .A2(new_n817), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n222), .A2(new_n863), .B1(new_n850), .B2(new_n1128), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G116), .B2(new_n837), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n542), .B1(new_n848), .B2(new_n336), .C1(new_n611), .C2(new_n893), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G97), .B2(new_n835), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(new_n202), .C2(new_n843), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n897), .A2(new_n1131), .ZN(new_n1203));
  INV_X1    g1003(.A(G125), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n897), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n845), .A2(G150), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT53), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n542), .B(new_n1207), .C1(G159), .C2(new_n847), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G128), .A2(new_n849), .B1(new_n837), .B2(G132), .ZN(new_n1209));
  XOR2_X1   g1009(.A(KEYINPUT54), .B(G143), .Z(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT117), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G137), .A2(new_n833), .B1(new_n835), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n842), .A2(G50), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1208), .A2(new_n1209), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1202), .A2(new_n1203), .B1(new_n1205), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n820), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n806), .B1(new_n252), .B2(new_n901), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1197), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1196), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1195), .A2(new_n1220), .ZN(G378));
  NAND2_X1  g1021(.A1(new_n369), .A2(new_n931), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1222), .B(KEYINPUT55), .Z(new_n1223));
  XNOR2_X1  g1023(.A(new_n465), .B(new_n1223), .ZN(new_n1224));
  XOR2_X1   g1024(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1225));
  XOR2_X1   g1025(.A(new_n1224), .B(new_n1225), .Z(new_n1226));
  OAI21_X1  g1026(.A(G330), .B1(new_n949), .B2(new_n959), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT122), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1226), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n970), .A2(new_n971), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n966), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n980), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT108), .ZN(new_n1234));
  OAI211_X1 g1034(.A(KEYINPUT122), .B(G330), .C1(new_n949), .C2(new_n959), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n972), .A2(new_n973), .A3(new_n980), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1234), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1230), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n925), .A2(new_n958), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT40), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n925), .A2(new_n948), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n777), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(KEYINPUT122), .C1(new_n981), .C2(new_n982), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1229), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1239), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1226), .A2(new_n817), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n901), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n805), .B1(G50), .B2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n843), .A2(new_n201), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1061), .B(new_n1251), .C1(G97), .C2(new_n833), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n542), .A2(new_n289), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n845), .B2(G77), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT118), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n222), .A2(new_n838), .B1(new_n850), .B2(new_n628), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(new_n590), .C2(new_n835), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1252), .B(new_n1257), .C1(new_n1128), .C2(new_n897), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT58), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1253), .B(new_n363), .C1(G33), .C2(G41), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n861), .A2(new_n883), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G132), .B2(new_n833), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n849), .A2(G125), .B1(G150), .B2(new_n847), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n837), .A2(G128), .B1(new_n1211), .B2(new_n845), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT119), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1262), .B(new_n1263), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1268), .A2(KEYINPUT59), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(KEYINPUT59), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n625), .B(new_n289), .C1(new_n843), .C2(new_n1067), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G124), .B2(new_n828), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1259), .B(new_n1260), .C1(new_n1269), .C2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT120), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1125), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1250), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1247), .A2(new_n804), .B1(new_n1248), .B2(new_n1278), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1244), .A2(new_n1229), .A3(new_n1245), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1229), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1180), .B1(new_n1170), .B2(new_n1181), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT57), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n800), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT57), .B1(new_n1247), .B2(new_n1283), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1279), .B1(new_n1285), .B2(new_n1286), .ZN(G375));
  OR2_X1    g1087(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1027), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1181), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n967), .A2(new_n817), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n805), .B1(G68), .B2(new_n1249), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n897), .A2(new_n651), .ZN(new_n1293));
  OAI22_X1  g1093(.A1(new_n222), .A2(new_n861), .B1(new_n850), .B2(new_n1131), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(G116), .B2(new_n833), .ZN(new_n1295));
  OAI221_X1 g1095(.A(new_n542), .B1(new_n848), .B2(new_n429), .C1(new_n580), .C2(new_n893), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(G283), .B2(new_n837), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1064), .A3(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n858), .A2(G128), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1251), .ZN(new_n1300));
  OAI221_X1 g1100(.A(new_n272), .B1(new_n848), .B2(new_n363), .C1(new_n1067), .C2(new_n893), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(G150), .B2(new_n835), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n833), .A2(new_n1211), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(G132), .A2(new_n849), .B1(new_n837), .B2(G137), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .A4(new_n1304), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n1293), .A2(new_n1298), .B1(new_n1299), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1292), .B1(new_n1306), .B2(new_n820), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1177), .A2(new_n804), .B1(new_n1291), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1290), .A2(new_n1308), .ZN(G381));
  NAND3_X1  g1109(.A1(new_n1088), .A2(new_n879), .A3(new_n1119), .ZN(new_n1310));
  NOR4_X1   g1110(.A1(G390), .A2(new_n1310), .A3(G384), .A4(G381), .ZN(new_n1311));
  INV_X1    g1111(.A(G387), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n804), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1278), .A2(new_n1248), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1283), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT57), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1187), .B2(new_n1180), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n744), .B1(new_n1247), .B2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1315), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1322), .A2(new_n1219), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1311), .A2(new_n1312), .A3(new_n1321), .A4(new_n1323), .ZN(G407));
  NAND2_X1  g1124(.A1(new_n712), .A2(G213), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1321), .A2(new_n1323), .A3(new_n1326), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1327), .B(KEYINPUT123), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(G213), .A3(G407), .ZN(G409));
  OAI21_X1  g1129(.A(new_n1279), .B1(new_n1027), .B2(new_n1316), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1323), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1219), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT124), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(G375), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(KEYINPUT124), .B1(G378), .B2(new_n1321), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1331), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1325), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1181), .A2(KEYINPUT60), .ZN(new_n1338));
  OR2_X1    g1138(.A1(new_n1338), .A2(new_n1288), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1288), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1339), .A2(new_n800), .A3(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1308), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(G384), .ZN(new_n1343));
  AND2_X1   g1143(.A1(new_n1326), .A2(G2897), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1343), .B(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT61), .B1(new_n1337), .B2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(G378), .A2(KEYINPUT124), .A3(new_n1321), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1333), .B1(G375), .B2(new_n1332), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1326), .B1(new_n1349), .B2(new_n1331), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1350), .A2(KEYINPUT62), .A3(new_n1343), .ZN(new_n1351));
  AOI21_X1  g1151(.A(KEYINPUT62), .B1(new_n1350), .B2(new_n1343), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1346), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(G390), .B1(new_n1057), .B2(new_n1085), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(G393), .A2(G396), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1310), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1057), .A2(G390), .A3(new_n1085), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1355), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1359), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1357), .B1(new_n1361), .B2(new_n1354), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1360), .A2(new_n1362), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1363), .B(KEYINPUT126), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1353), .A2(new_n1364), .ZN(new_n1365));
  AND2_X1   g1165(.A1(new_n1343), .A2(KEYINPUT63), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1336), .A2(new_n1325), .A3(new_n1366), .ZN(new_n1367));
  AND2_X1   g1167(.A1(new_n1360), .A2(new_n1362), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(KEYINPUT63), .B1(new_n1350), .B2(new_n1343), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  AOI21_X1  g1171(.A(KEYINPUT125), .B1(new_n1371), .B2(new_n1346), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1363), .B1(new_n1350), .B2(new_n1366), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1336), .A2(new_n1325), .A3(new_n1343), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT63), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  AND4_X1   g1176(.A1(KEYINPUT125), .A2(new_n1346), .A3(new_n1373), .A4(new_n1376), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1365), .B1(new_n1372), .B2(new_n1377), .ZN(G405));
  XNOR2_X1  g1178(.A(new_n1363), .B(new_n1343), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(G375), .A2(new_n1323), .ZN(new_n1380));
  XNOR2_X1  g1180(.A(new_n1380), .B(KEYINPUT127), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1381), .A2(new_n1349), .ZN(new_n1382));
  XNOR2_X1  g1182(.A(new_n1379), .B(new_n1382), .ZN(G402));
endmodule


