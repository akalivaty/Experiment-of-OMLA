//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G146), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G143), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n189), .B(G146), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n196), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(G143), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(new_n193), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n190), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n195), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G137), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n211), .B2(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(G134), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(new_n214), .ZN(new_n219));
  AOI211_X1 g033(.A(G131), .B(new_n213), .C1(new_n216), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n219), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n210), .A2(new_n212), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n201), .B(new_n208), .C1(new_n220), .C2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT67), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n194), .A2(new_n200), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n230), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n190), .A2(G146), .ZN(new_n234));
  OAI21_X1  g048(.A(G128), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n206), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n221), .B1(new_n217), .B2(new_n212), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n213), .B1(new_n216), .B2(new_n219), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n238), .B1(new_n239), .B2(new_n221), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT68), .B(G119), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G119), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G116), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT2), .B(G113), .Z(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n242), .A2(new_n243), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(new_n246), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n225), .A2(new_n241), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT69), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n225), .A2(new_n241), .A3(new_n256), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n225), .A2(new_n241), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n249), .A2(new_n252), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n225), .A2(new_n241), .A3(KEYINPUT30), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G953), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G237), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(G210), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT27), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT27), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n269), .A2(new_n273), .A3(G210), .A4(new_n270), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT26), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n272), .A2(new_n277), .A3(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G101), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n276), .A2(new_n278), .A3(G101), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n258), .A2(new_n264), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT31), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n258), .A2(new_n264), .A3(new_n284), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n253), .B1(new_n225), .B2(new_n241), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n201), .A2(new_n208), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n218), .B1(new_n217), .B2(new_n214), .ZN(new_n293));
  AOI211_X1 g107(.A(KEYINPUT66), .B(KEYINPUT11), .C1(new_n209), .C2(G134), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n223), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G131), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n239), .A2(new_n221), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n292), .A2(new_n298), .B1(new_n237), .B2(new_n240), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n256), .B1(new_n299), .B2(new_n253), .ZN(new_n300));
  INV_X1    g114(.A(new_n257), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n291), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT28), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n254), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n284), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n188), .B1(new_n289), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n305), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(new_n302), .B2(KEYINPUT28), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n286), .B(new_n288), .C1(new_n311), .C2(new_n284), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT32), .A3(new_n188), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G472), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n283), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n290), .B1(new_n255), .B2(new_n257), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n305), .B(new_n317), .C1(new_n318), .C2(new_n304), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  INV_X1    g134(.A(G902), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n319), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n305), .B1(new_n318), .B2(new_n304), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n284), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n258), .A2(new_n264), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n283), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n316), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n315), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n187), .B1(new_n314), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n319), .A2(new_n321), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT71), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT29), .B1(new_n326), .B2(new_n328), .ZN(new_n337));
  OAI21_X1  g151(.A(G472), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n338), .A2(KEYINPUT72), .A3(new_n309), .A4(new_n313), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G217), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(G234), .B2(new_n321), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G125), .ZN(new_n345));
  INV_X1    g159(.A(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G140), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n347), .A3(KEYINPUT16), .ZN(new_n348));
  OR3_X1    g162(.A1(new_n346), .A2(KEYINPUT16), .A3(G140), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(G146), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n345), .A2(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n193), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT68), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G119), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n226), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n245), .A2(G128), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT73), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT73), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n242), .B2(new_n226), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(KEYINPUT24), .A2(G110), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT24), .A2(G110), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(KEYINPUT74), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT74), .ZN(new_n366));
  AND2_X1   g180(.A1(KEYINPUT24), .A2(G110), .ZN(new_n367));
  NOR2_X1   g181(.A1(KEYINPUT24), .A2(G110), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT23), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G128), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G119), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(G128), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n375), .B(new_n376), .C1(new_n242), .C2(new_n374), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n377), .A2(G110), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n353), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n348), .A2(new_n349), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n193), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT75), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n350), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n359), .A2(new_n370), .A3(new_n361), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT75), .A4(G146), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n377), .A2(G110), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n388), .A2(new_n389), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n380), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT22), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n209), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n393), .A2(KEYINPUT22), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(KEYINPUT22), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(G137), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n392), .A2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n348), .A2(G146), .A3(new_n349), .ZN(new_n401));
  AOI21_X1  g215(.A(G146), .B1(new_n348), .B2(new_n349), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT75), .ZN(new_n403));
  INV_X1    g217(.A(new_n386), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n405), .A2(KEYINPUT76), .A3(new_n385), .A4(new_n387), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n388), .A2(new_n389), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n399), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n380), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n321), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT25), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n400), .A2(KEYINPUT25), .A3(new_n410), .A4(new_n321), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n343), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n409), .B1(new_n408), .B2(new_n380), .ZN(new_n416));
  AOI211_X1 g230(.A(new_n379), .B(new_n399), .C1(new_n406), .C2(new_n407), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n342), .A2(G902), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n340), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT77), .ZN(new_n423));
  INV_X1    g237(.A(new_n421), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n332), .B2(new_n339), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT77), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g241(.A(KEYINPUT9), .B(G234), .Z(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G221), .B1(new_n429), .B2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G469), .ZN(new_n432));
  XOR2_X1   g246(.A(G110), .B(G140), .Z(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT78), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n269), .A2(G227), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G107), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT79), .B1(new_n437), .B2(G104), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n439));
  INV_X1    g253(.A(G104), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(G107), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT3), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n440), .B2(G107), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(KEYINPUT3), .A3(G104), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n438), .A2(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT80), .B1(new_n445), .B2(new_n280), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n438), .A2(new_n441), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n444), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT80), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(G101), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n280), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n446), .A2(new_n451), .A3(KEYINPUT4), .A4(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(G101), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n292), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT82), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n453), .A2(new_n292), .A3(new_n458), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT83), .B1(new_n437), .B2(G104), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n440), .B2(G107), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n437), .A2(KEYINPUT83), .A3(G104), .ZN(new_n463));
  OAI21_X1  g277(.A(G101), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n452), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n194), .A2(new_n200), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n227), .B1(new_n192), .B2(new_n193), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n226), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n465), .B1(new_n468), .B2(new_n232), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT84), .B(KEYINPUT10), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n465), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT10), .A3(new_n237), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n460), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n298), .ZN(new_n475));
  INV_X1    g289(.A(new_n298), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n460), .A2(new_n471), .A3(new_n476), .A4(new_n473), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n436), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n472), .A2(new_n237), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n298), .B1(new_n479), .B2(new_n469), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT12), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(KEYINPUT12), .B(new_n298), .C1(new_n479), .C2(new_n469), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n477), .A2(new_n484), .A3(new_n436), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n432), .B(new_n321), .C1(new_n478), .C2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n477), .A3(new_n436), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n477), .A2(new_n484), .ZN(new_n489));
  INV_X1    g303(.A(new_n436), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G469), .B1(new_n492), .B2(G902), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n487), .B1(new_n493), .B2(KEYINPUT85), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n495), .B(G469), .C1(new_n492), .C2(G902), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n431), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n269), .A2(G214), .A3(new_n270), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n192), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n269), .A2(new_n190), .A3(G214), .A4(new_n270), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(G131), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT89), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n499), .A2(new_n503), .A3(G131), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n499), .A2(new_n500), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n221), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT91), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n502), .A2(new_n504), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n405), .B1(new_n511), .B2(KEYINPUT17), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n505), .A2(new_n513), .A3(new_n506), .A4(new_n508), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n507), .A2(KEYINPUT88), .ZN(new_n516));
  NAND2_X1  g330(.A1(KEYINPUT18), .A2(G131), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n516), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n351), .B(G146), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G113), .B(G122), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n440), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n515), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n524), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n351), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n528), .B(KEYINPUT19), .Z(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n350), .B1(new_n530), .B2(G146), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n508), .B2(new_n505), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n526), .B1(new_n532), .B2(new_n521), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(G475), .A2(G902), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT20), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT20), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(new_n538), .A3(new_n535), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n515), .A2(new_n524), .A3(new_n522), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n524), .B1(new_n515), .B2(new_n522), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n321), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n537), .A2(new_n539), .B1(G475), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n544));
  OAI21_X1  g358(.A(G128), .B1(new_n198), .B2(new_n199), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n190), .A2(G128), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G134), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n211), .A3(new_n547), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n243), .A2(G122), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n437), .B1(new_n552), .B2(KEYINPUT14), .ZN(new_n553));
  XNOR2_X1  g367(.A(G116), .B(G122), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT13), .B(new_n547), .C1(new_n192), .C2(new_n226), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n557), .B(G134), .C1(new_n545), .C2(KEYINPUT13), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n554), .B(new_n437), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n550), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n428), .A2(G217), .A3(new_n265), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n564));
  INV_X1    g378(.A(new_n562), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n556), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n556), .A2(new_n560), .A3(KEYINPUT92), .A4(new_n565), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n321), .ZN(new_n569));
  INV_X1    g383(.A(G478), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT15), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n544), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n569), .A2(new_n571), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(KEYINPUT93), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n567), .A2(new_n568), .A3(new_n575), .A4(new_n321), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n573), .B1(new_n577), .B2(new_n571), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n572), .B1(new_n578), .B2(new_n544), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G214), .B1(G237), .B2(G902), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n244), .A2(KEYINPUT5), .A3(new_n247), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n583), .B(G113), .C1(KEYINPUT5), .C2(new_n244), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n249), .A3(new_n472), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n453), .A2(new_n262), .A3(new_n455), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(G110), .B(G122), .Z(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(KEYINPUT6), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT6), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n587), .A2(new_n593), .A3(new_n588), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n237), .A2(G125), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n346), .B1(new_n201), .B2(new_n208), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n595), .A2(KEYINPUT86), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(G224), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(G953), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT86), .B1(new_n595), .B2(new_n596), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n600), .B1(new_n598), .B2(new_n601), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n592), .B(new_n594), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n588), .B(KEYINPUT8), .Z(new_n605));
  INV_X1    g419(.A(new_n585), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n472), .B1(new_n584), .B2(new_n249), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n595), .A2(new_n596), .ZN(new_n609));
  INV_X1    g423(.A(new_n600), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT7), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n609), .A2(new_n611), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n608), .B(new_n591), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n604), .A2(new_n321), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G210), .B1(G237), .B2(G902), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT87), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n617), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n604), .A2(new_n321), .A3(new_n619), .A4(new_n614), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n582), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(G234), .A2(G237), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n622), .A2(G952), .A3(new_n265), .ZN(new_n623));
  INV_X1    g437(.A(new_n269), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(G902), .A3(new_n622), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n625), .B(KEYINPUT95), .Z(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT21), .B(G898), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AND4_X1   g445(.A1(new_n497), .A2(new_n543), .A3(new_n580), .A4(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n423), .A2(new_n427), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  NAND2_X1  g448(.A1(new_n493), .A2(KEYINPUT85), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n496), .A3(new_n486), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n430), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n312), .A2(new_n321), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(G472), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n307), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n637), .A2(new_n424), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n542), .A2(G475), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n538), .B1(new_n534), .B2(new_n535), .ZN(new_n643));
  INV_X1    g457(.A(new_n535), .ZN(new_n644));
  AOI211_X1 g458(.A(KEYINPUT20), .B(new_n644), .C1(new_n525), .C2(new_n533), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n642), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n574), .A2(new_n570), .A3(new_n576), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n566), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n563), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n566), .A2(new_n648), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT33), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n567), .A2(new_n568), .ZN(new_n653));
  OAI211_X1 g467(.A(G478), .B(new_n652), .C1(new_n653), .C2(KEYINPUT33), .ZN(new_n654));
  NAND2_X1  g468(.A1(G478), .A2(G902), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n647), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT97), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n647), .A2(new_n654), .A3(new_n658), .A4(new_n655), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n646), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n630), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n641), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT98), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT34), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n440), .ZN(G6));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n537), .A2(new_n666), .A3(new_n539), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n645), .A2(KEYINPUT99), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n667), .A2(new_n579), .A3(new_n642), .A4(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n630), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n641), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  INV_X1    g487(.A(new_n640), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT25), .B1(new_n418), .B2(new_n321), .ZN(new_n675));
  INV_X1    g489(.A(new_n414), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n342), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n399), .A2(KEYINPUT36), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n392), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n419), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT100), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n680), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n415), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n632), .A2(new_n674), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT37), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G110), .ZN(G12));
  OAI21_X1  g504(.A(new_n621), .B1(new_n681), .B2(new_n685), .ZN(new_n691));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n626), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n623), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n542), .B2(G475), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n667), .A2(new_n579), .A3(new_n668), .A4(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n340), .A2(new_n697), .A3(new_n497), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XNOR2_X1  g513(.A(new_n694), .B(KEYINPUT39), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n637), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n618), .A2(new_n620), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT38), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n646), .A2(new_n579), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n705), .A2(new_n582), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n701), .A2(new_n702), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n302), .A2(new_n284), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n283), .B1(new_n258), .B2(new_n264), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n318), .A2(new_n283), .ZN(new_n713));
  OAI211_X1 g527(.A(KEYINPUT101), .B(new_n713), .C1(new_n327), .C2(new_n283), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n714), .A3(new_n321), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G472), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n309), .A2(new_n716), .A3(new_n313), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n677), .A2(new_n680), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n703), .A2(new_n707), .A3(new_n708), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n192), .ZN(G45));
  INV_X1    g536(.A(new_n691), .ZN(new_n723));
  INV_X1    g537(.A(new_n694), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n646), .A2(new_n657), .A3(new_n659), .A4(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n340), .A2(new_n497), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  NOR2_X1   g542(.A1(new_n478), .A2(new_n485), .ZN(new_n729));
  OAI21_X1  g543(.A(G469), .B1(new_n729), .B2(G902), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n430), .A3(new_n486), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n340), .A2(new_n421), .A3(new_n661), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  NAND4_X1  g549(.A1(new_n340), .A2(new_n421), .A3(new_n670), .A4(new_n732), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  NOR2_X1   g551(.A1(new_n691), .A2(new_n731), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n646), .A2(new_n579), .A3(new_n628), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n340), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  NAND2_X1  g555(.A1(new_n325), .A2(KEYINPUT103), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n743), .B(new_n305), .C1(new_n318), .C2(new_n304), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n742), .A2(new_n283), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n188), .B1(new_n745), .B2(new_n289), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n421), .A3(new_n639), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT104), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n746), .A2(new_n639), .A3(new_n421), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n704), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n706), .A2(new_n582), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n751), .A2(new_n629), .A3(new_n753), .A4(new_n732), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G122), .ZN(G24));
  NAND3_X1  g569(.A1(new_n746), .A2(new_n719), .A3(new_n639), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n725), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n621), .A3(new_n732), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G125), .ZN(G27));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n488), .A2(new_n491), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT106), .B1(new_n489), .B2(new_n490), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n763), .A3(G469), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(G469), .A2(G902), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT105), .Z(new_n768));
  AND2_X1   g582(.A1(new_n486), .A2(new_n763), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n432), .B(new_n764), .C1(new_n761), .C2(KEYINPUT106), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n766), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n431), .A2(new_n582), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n752), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n314), .A2(new_n331), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n775), .B2(new_n424), .ZN(new_n776));
  OAI211_X1 g590(.A(KEYINPUT108), .B(new_n421), .C1(new_n314), .C2(new_n331), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n760), .B1(new_n778), .B2(new_n726), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n771), .A2(new_n752), .A3(new_n772), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n425), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n726), .A2(new_n760), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G131), .ZN(G33));
  NOR3_X1   g599(.A1(new_n422), .A2(new_n696), .A3(new_n773), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n211), .ZN(G36));
  NAND3_X1  g601(.A1(new_n762), .A2(KEYINPUT45), .A3(new_n765), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n788), .B(G469), .C1(KEYINPUT45), .C2(new_n492), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n768), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n487), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n768), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n431), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n700), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n618), .A2(new_n581), .A3(new_n620), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n657), .A2(new_n659), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n646), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT43), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n640), .A3(new_n719), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n799), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n794), .A2(KEYINPUT109), .A3(new_n795), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n803), .A2(new_n804), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n798), .A2(new_n805), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT47), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n794), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n810), .A2(KEYINPUT47), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n811), .B1(new_n794), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n340), .A2(new_n421), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n725), .A2(new_n799), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n812), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT111), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n344), .ZN(G42));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  INV_X1    g634(.A(new_n727), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n698), .A2(new_n758), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n698), .A2(KEYINPUT114), .A3(new_n758), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n415), .A2(new_n683), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n694), .B(KEYINPUT115), .Z(new_n828));
  AND4_X1   g642(.A1(new_n430), .A2(new_n717), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n753), .A3(new_n771), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n820), .B1(new_n826), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n727), .A2(new_n698), .A3(new_n830), .A4(new_n758), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n754), .A2(new_n733), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n736), .A2(new_n740), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n733), .A2(new_n754), .A3(new_n736), .A4(new_n740), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT112), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n779), .A2(new_n783), .A3(new_n786), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n667), .A2(new_n668), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n682), .B2(new_n686), .ZN(new_n845));
  INV_X1    g659(.A(new_n799), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n846), .A2(new_n580), .A3(new_n695), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n340), .A2(new_n497), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n757), .A2(new_n752), .A3(new_n772), .A4(new_n771), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n660), .B1(new_n646), .B2(new_n580), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT113), .B1(new_n580), .B2(new_n646), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n631), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT113), .B1(new_n660), .B2(new_n630), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n641), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n633), .A2(new_n850), .A3(new_n688), .A4(new_n856), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n835), .A2(new_n842), .A3(new_n843), .A4(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n698), .A2(KEYINPUT114), .A3(new_n758), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT114), .B1(new_n698), .B2(new_n758), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n727), .B(new_n830), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT52), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n863));
  INV_X1    g677(.A(new_n833), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n834), .A2(new_n858), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n776), .A2(new_n777), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n726), .A3(new_n780), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT42), .ZN(new_n869));
  INV_X1    g683(.A(new_n786), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n869), .B(new_n870), .C1(new_n781), .C2(new_n782), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n633), .A2(new_n850), .A3(new_n688), .A4(new_n856), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n864), .A3(new_n842), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT53), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n866), .A2(KEYINPUT54), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n840), .A2(new_n835), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n857), .A2(new_n843), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n834), .A2(new_n865), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n875), .A2(new_n835), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n877), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n802), .A2(new_n623), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n731), .A2(new_n799), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(new_n867), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT48), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(KEYINPUT48), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n731), .B1(new_n748), .B2(new_n750), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(new_n621), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(G952), .A3(new_n265), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n886), .A2(new_n582), .A3(new_n705), .A4(new_n892), .ZN(new_n896));
  NOR2_X1   g710(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n888), .A2(new_n639), .A3(new_n719), .A4(new_n746), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n887), .A2(new_n421), .A3(new_n718), .A4(new_n623), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n543), .A3(new_n800), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT51), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n886), .A2(new_n751), .A3(new_n846), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n812), .A2(new_n814), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n730), .A2(new_n431), .A3(new_n486), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n890), .B(new_n895), .C1(new_n904), .C2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n905), .ZN(new_n910));
  INV_X1    g724(.A(new_n906), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n907), .B(KEYINPUT117), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT51), .B1(new_n903), .B2(new_n913), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n885), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n900), .A2(new_n660), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n915), .A2(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n421), .A2(new_n705), .A3(new_n718), .A4(new_n772), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n730), .A2(new_n486), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT49), .Z(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n801), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n917), .A2(new_n921), .ZN(G75));
  NAND2_X1  g736(.A1(new_n592), .A2(new_n594), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT119), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n321), .B(new_n619), .C1(new_n881), .C2(new_n882), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n602), .A2(new_n603), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n926), .A2(KEYINPUT56), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n321), .B1(new_n881), .B2(new_n882), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n617), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n925), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n269), .A2(G952), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n929), .B1(new_n926), .B2(KEYINPUT56), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n933), .A3(new_n928), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n938), .A3(new_n924), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(G51));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n768), .B(KEYINPUT57), .Z(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n863), .B1(new_n862), .B2(new_n864), .ZN(new_n944));
  AOI211_X1 g758(.A(KEYINPUT116), .B(new_n833), .C1(new_n861), .C2(KEYINPUT52), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n945), .A3(new_n879), .ZN(new_n946));
  AND4_X1   g760(.A1(new_n842), .A2(new_n857), .A3(new_n843), .A4(new_n874), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT53), .B1(new_n947), .B2(new_n864), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT54), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n943), .B1(new_n949), .B2(new_n884), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n941), .B1(new_n950), .B2(new_n729), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n881), .A2(new_n883), .A3(new_n882), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n883), .B1(new_n881), .B2(new_n882), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n942), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n729), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(KEYINPUT120), .A3(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n931), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(new_n789), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n951), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(new_n936), .ZN(G54));
  NAND3_X1  g774(.A1(new_n931), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  INV_X1    g775(.A(new_n534), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n963), .A2(new_n936), .A3(new_n964), .ZN(G60));
  XOR2_X1   g779(.A(new_n655), .B(KEYINPUT59), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n885), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT122), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n653), .A2(KEYINPUT33), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n650), .A2(new_n651), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(KEYINPUT33), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n968), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n966), .B1(new_n877), .B2(new_n884), .ZN(new_n974));
  INV_X1    g788(.A(new_n972), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT122), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n975), .B(new_n967), .C1(new_n952), .C2(new_n953), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT121), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n966), .B1(new_n949), .B2(new_n884), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(KEYINPUT121), .A3(new_n975), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n977), .A2(new_n983), .A3(new_n936), .ZN(G63));
  NAND2_X1  g798(.A1(new_n881), .A2(new_n882), .ZN(new_n985));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT60), .Z(new_n987));
  NAND3_X1  g801(.A1(new_n985), .A2(new_n679), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n985), .A2(new_n987), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n936), .B(new_n988), .C1(new_n989), .C2(new_n418), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g805(.A(G953), .B1(new_n627), .B2(new_n599), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n633), .A2(new_n688), .A3(new_n856), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n842), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n995), .B2(new_n624), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n924), .B1(G898), .B2(new_n269), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT123), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n996), .B(new_n998), .ZN(G69));
  NAND2_X1  g813(.A1(new_n261), .A2(new_n263), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(new_n530), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n826), .A2(new_n721), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n826), .A2(KEYINPUT62), .A3(new_n721), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n808), .A2(new_n817), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n423), .A2(new_n427), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1008), .A2(new_n701), .A3(new_n846), .A4(new_n851), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT124), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1006), .A2(new_n1007), .A3(KEYINPUT124), .A4(new_n1009), .ZN(new_n1013));
  AOI211_X1 g827(.A(new_n624), .B(new_n1001), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(G900), .B1(new_n1001), .B2(G227), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n624), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n808), .A2(new_n817), .A3(new_n826), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n798), .A2(new_n753), .A3(new_n867), .A4(new_n806), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n843), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n269), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n1001), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n269), .A2(G227), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1016), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n1014), .A2(new_n1023), .ZN(G72));
  NAND3_X1  g838(.A1(new_n1012), .A2(new_n995), .A3(new_n1013), .ZN(new_n1025));
  XNOR2_X1  g839(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n315), .A2(new_n321), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(new_n711), .ZN(new_n1030));
  INV_X1    g844(.A(new_n711), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1028), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(new_n327), .B2(new_n283), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n866), .A2(new_n876), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n328), .B(KEYINPUT126), .Z(new_n1035));
  NOR3_X1   g849(.A1(new_n1017), .A2(new_n1019), .A3(new_n994), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1035), .B1(new_n1036), .B2(new_n1032), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1030), .A2(new_n936), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT127), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n1030), .A2(KEYINPUT127), .A3(new_n936), .A4(new_n1038), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1041), .A2(new_n1042), .ZN(G57));
endmodule


