

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  AND2_X1 U325 ( .A1(n563), .A2(n513), .ZN(n402) );
  XOR2_X1 U326 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n293) );
  AND2_X1 U327 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U328 ( .A(n386), .B(n385), .Z(n295) );
  AND2_X1 U329 ( .A1(n562), .A2(n576), .ZN(n452) );
  XNOR2_X1 U330 ( .A(KEYINPUT25), .B(KEYINPUT98), .ZN(n403) );
  XNOR2_X1 U331 ( .A(n404), .B(n403), .ZN(n409) );
  XNOR2_X1 U332 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(n465) );
  INV_X1 U334 ( .A(G176GAT), .ZN(n389) );
  XNOR2_X1 U335 ( .A(n422), .B(n294), .ZN(n423) );
  XNOR2_X1 U336 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U337 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U338 ( .A(n392), .B(n391), .ZN(n396) );
  NOR2_X1 U339 ( .A1(n540), .A2(n555), .ZN(n587) );
  XOR2_X1 U340 ( .A(n400), .B(n399), .Z(n563) );
  XNOR2_X1 U341 ( .A(n470), .B(G218GAT), .ZN(n471) );
  XNOR2_X1 U342 ( .A(n449), .B(G43GAT), .ZN(n450) );
  XNOR2_X1 U343 ( .A(n472), .B(n471), .ZN(G1355GAT) );
  XNOR2_X1 U344 ( .A(n451), .B(n450), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT7), .B(G50GAT), .Z(n297) );
  XNOR2_X1 U346 ( .A(G36GAT), .B(G29GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U348 ( .A(KEYINPUT8), .B(n298), .ZN(n445) );
  INV_X1 U349 ( .A(n445), .ZN(n317) );
  XOR2_X1 U350 ( .A(KEYINPUT79), .B(KEYINPUT76), .Z(n300) );
  XNOR2_X1 U351 ( .A(G190GAT), .B(KEYINPUT9), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U353 ( .A(KEYINPUT10), .B(KEYINPUT75), .Z(n302) );
  XNOR2_X1 U354 ( .A(G106GAT), .B(KEYINPUT64), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U356 ( .A(n304), .B(n303), .Z(n315) );
  XOR2_X1 U357 ( .A(KEYINPUT77), .B(G162GAT), .Z(n306) );
  XNOR2_X1 U358 ( .A(G134GAT), .B(G99GAT), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n313) );
  XOR2_X1 U360 ( .A(G85GAT), .B(G92GAT), .Z(n416) );
  XOR2_X1 U361 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n308) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(G218GAT), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U364 ( .A(n416), .B(n309), .Z(n311) );
  NAND2_X1 U365 ( .A1(G232GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U369 ( .A(n317), .B(n316), .Z(n473) );
  INV_X1 U370 ( .A(n473), .ZN(n572) );
  XOR2_X1 U371 ( .A(n572), .B(KEYINPUT36), .Z(n469) );
  XOR2_X1 U372 ( .A(G64GAT), .B(G78GAT), .Z(n319) );
  XNOR2_X1 U373 ( .A(G22GAT), .B(G71GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U375 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n321) );
  XNOR2_X1 U376 ( .A(KEYINPUT82), .B(KEYINPUT81), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n333) );
  XNOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n324), .B(KEYINPUT69), .ZN(n425) );
  XOR2_X1 U381 ( .A(KEYINPUT80), .B(G211GAT), .Z(n326) );
  XNOR2_X1 U382 ( .A(G8GAT), .B(G183GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n365) );
  XOR2_X1 U384 ( .A(KEYINPUT14), .B(n365), .Z(n328) );
  NAND2_X1 U385 ( .A1(G231GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U387 ( .A(n425), .B(n329), .Z(n331) );
  XOR2_X1 U388 ( .A(G15GAT), .B(G127GAT), .Z(n385) );
  XOR2_X1 U389 ( .A(G1GAT), .B(G155GAT), .Z(n339) );
  XNOR2_X1 U390 ( .A(n385), .B(n339), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U392 ( .A(n333), .B(n332), .Z(n459) );
  INV_X1 U393 ( .A(n459), .ZN(n586) );
  XOR2_X1 U394 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n335) );
  XNOR2_X1 U395 ( .A(G127GAT), .B(G57GAT), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n343) );
  XOR2_X1 U397 ( .A(G148GAT), .B(G120GAT), .Z(n337) );
  XNOR2_X1 U398 ( .A(G141GAT), .B(G113GAT), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U400 ( .A(n338), .B(G85GAT), .Z(n341) );
  XNOR2_X1 U401 ( .A(G29GAT), .B(n339), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n353) );
  XOR2_X1 U404 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n345) );
  NAND2_X1 U405 ( .A1(G225GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U407 ( .A(n346), .B(KEYINPUT4), .Z(n351) );
  XNOR2_X1 U408 ( .A(G134GAT), .B(KEYINPUT85), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n347), .B(KEYINPUT0), .ZN(n398) );
  XOR2_X1 U410 ( .A(KEYINPUT3), .B(KEYINPUT93), .Z(n349) );
  XNOR2_X1 U411 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n380) );
  XNOR2_X1 U413 ( .A(n398), .B(n380), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U415 ( .A(n353), .B(n352), .Z(n511) );
  INV_X1 U416 ( .A(n511), .ZN(n489) );
  XOR2_X1 U417 ( .A(G176GAT), .B(G64GAT), .Z(n417) );
  XOR2_X1 U418 ( .A(G92GAT), .B(G204GAT), .Z(n355) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(G36GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U421 ( .A(n417), .B(n356), .Z(n358) );
  NAND2_X1 U422 ( .A1(G226GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U424 ( .A(n359), .B(KEYINPUT96), .Z(n363) );
  XOR2_X1 U425 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n361) );
  XNOR2_X1 U426 ( .A(G197GAT), .B(G218GAT), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n375), .B(KEYINPUT95), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n367) );
  XNOR2_X1 U430 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n293), .B(n364), .ZN(n386) );
  XOR2_X1 U432 ( .A(n386), .B(n365), .Z(n366) );
  XOR2_X1 U433 ( .A(n367), .B(n366), .Z(n513) );
  XOR2_X1 U434 ( .A(KEYINPUT27), .B(n513), .Z(n407) );
  NOR2_X1 U435 ( .A1(n489), .A2(n407), .ZN(n541) );
  XOR2_X1 U436 ( .A(G141GAT), .B(G22GAT), .Z(n432) );
  XOR2_X1 U437 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n369) );
  XNOR2_X1 U438 ( .A(G50GAT), .B(G155GAT), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U440 ( .A(n432), .B(n370), .Z(n372) );
  NAND2_X1 U441 ( .A1(G228GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n372), .B(n371), .ZN(n384) );
  XOR2_X1 U443 ( .A(G211GAT), .B(KEYINPUT90), .Z(n374) );
  XNOR2_X1 U444 ( .A(KEYINPUT22), .B(KEYINPUT91), .ZN(n373) );
  XNOR2_X1 U445 ( .A(n374), .B(n373), .ZN(n376) );
  XOR2_X1 U446 ( .A(n376), .B(n375), .Z(n382) );
  XOR2_X1 U447 ( .A(G148GAT), .B(G106GAT), .Z(n378) );
  XNOR2_X1 U448 ( .A(G204GAT), .B(G78GAT), .ZN(n377) );
  XNOR2_X1 U449 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U450 ( .A(KEYINPUT71), .B(n379), .Z(n427) );
  XNOR2_X1 U451 ( .A(n427), .B(n380), .ZN(n381) );
  XNOR2_X1 U452 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U453 ( .A(n384), .B(n383), .ZN(n556) );
  XNOR2_X1 U454 ( .A(KEYINPUT28), .B(n556), .ZN(n518) );
  INV_X1 U455 ( .A(n518), .ZN(n496) );
  NAND2_X1 U456 ( .A1(n541), .A2(n496), .ZN(n524) );
  NAND2_X1 U457 ( .A1(G227GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n295), .B(n387), .ZN(n392) );
  XNOR2_X1 U459 ( .A(G99GAT), .B(G71GAT), .ZN(n388) );
  XNOR2_X1 U460 ( .A(n388), .B(G120GAT), .ZN(n428) );
  XNOR2_X1 U461 ( .A(n428), .B(G183GAT), .ZN(n390) );
  XOR2_X1 U462 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n394) );
  XNOR2_X1 U463 ( .A(KEYINPUT88), .B(KEYINPUT86), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U465 ( .A(n396), .B(n395), .Z(n400) );
  XNOR2_X1 U466 ( .A(G169GAT), .B(G43GAT), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n397), .B(G113GAT), .ZN(n431) );
  XNOR2_X1 U468 ( .A(n431), .B(n398), .ZN(n399) );
  XOR2_X1 U469 ( .A(KEYINPUT89), .B(n563), .Z(n401) );
  NOR2_X1 U470 ( .A1(n524), .A2(n401), .ZN(n412) );
  OR2_X1 U471 ( .A1(n556), .A2(n402), .ZN(n404) );
  XOR2_X1 U472 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n406) );
  INV_X1 U473 ( .A(n563), .ZN(n558) );
  NAND2_X1 U474 ( .A1(n558), .A2(n556), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n540) );
  NOR2_X1 U476 ( .A1(n540), .A2(n407), .ZN(n408) );
  NOR2_X1 U477 ( .A1(n409), .A2(n408), .ZN(n410) );
  NOR2_X1 U478 ( .A1(n410), .A2(n511), .ZN(n411) );
  NOR2_X1 U479 ( .A1(n412), .A2(n411), .ZN(n477) );
  NOR2_X1 U480 ( .A1(n586), .A2(n477), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n413), .B(KEYINPUT101), .ZN(n414) );
  NOR2_X1 U482 ( .A1(n469), .A2(n414), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n415), .B(KEYINPUT37), .ZN(n510) );
  XOR2_X1 U484 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n419) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n424) );
  XOR2_X1 U487 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n421) );
  XNOR2_X1 U488 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n420) );
  XOR2_X1 U489 ( .A(n421), .B(n420), .Z(n422) );
  XNOR2_X1 U490 ( .A(n426), .B(n425), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n580) );
  XOR2_X1 U493 ( .A(G15GAT), .B(n431), .Z(n434) );
  XNOR2_X1 U494 ( .A(n432), .B(G197GAT), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U496 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n436) );
  NAND2_X1 U497 ( .A1(G229GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U499 ( .A(n438), .B(n437), .Z(n443) );
  XOR2_X1 U500 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n440) );
  XNOR2_X1 U501 ( .A(G8GAT), .B(G1GAT), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n441), .B(KEYINPUT66), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U505 ( .A(n445), .B(n444), .Z(n576) );
  INV_X1 U506 ( .A(n576), .ZN(n498) );
  XOR2_X1 U507 ( .A(KEYINPUT68), .B(n498), .Z(n559) );
  NAND2_X1 U508 ( .A1(n580), .A2(n559), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n446), .B(KEYINPUT74), .ZN(n480) );
  NOR2_X1 U510 ( .A1(n510), .A2(n480), .ZN(n448) );
  XOR2_X1 U511 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n447) );
  XNOR2_X1 U512 ( .A(n448), .B(n447), .ZN(n495) );
  NOR2_X1 U513 ( .A1(n495), .A2(n558), .ZN(n451) );
  XNOR2_X1 U514 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n449) );
  INV_X1 U515 ( .A(n513), .ZN(n493) );
  XOR2_X1 U516 ( .A(KEYINPUT110), .B(n459), .Z(n570) );
  XOR2_X1 U517 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n453) );
  XNOR2_X1 U518 ( .A(KEYINPUT41), .B(n580), .ZN(n562) );
  XNOR2_X1 U519 ( .A(n453), .B(n452), .ZN(n454) );
  NOR2_X1 U520 ( .A1(n570), .A2(n454), .ZN(n455) );
  XNOR2_X1 U521 ( .A(KEYINPUT112), .B(n455), .ZN(n456) );
  NAND2_X1 U522 ( .A1(n456), .A2(n473), .ZN(n458) );
  NOR2_X1 U523 ( .A1(n459), .A2(n469), .ZN(n460) );
  XNOR2_X1 U524 ( .A(KEYINPUT45), .B(n460), .ZN(n461) );
  NAND2_X1 U525 ( .A1(n461), .A2(n580), .ZN(n462) );
  XOR2_X1 U526 ( .A(KEYINPUT114), .B(n462), .Z(n463) );
  INV_X1 U527 ( .A(n559), .ZN(n526) );
  NAND2_X1 U528 ( .A1(n463), .A2(n526), .ZN(n464) );
  NAND2_X1 U529 ( .A1(n465), .A2(n464), .ZN(n466) );
  XOR2_X1 U530 ( .A(n466), .B(KEYINPUT48), .Z(n539) );
  NOR2_X1 U531 ( .A1(n493), .A2(n539), .ZN(n467) );
  XNOR2_X1 U532 ( .A(n467), .B(KEYINPUT54), .ZN(n468) );
  NAND2_X1 U533 ( .A1(n468), .A2(n489), .ZN(n555) );
  INV_X1 U534 ( .A(n587), .ZN(n581) );
  NOR2_X1 U535 ( .A1(n469), .A2(n581), .ZN(n472) );
  XNOR2_X1 U536 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n470) );
  XOR2_X1 U537 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n482) );
  NAND2_X1 U538 ( .A1(n473), .A2(n586), .ZN(n476) );
  XNOR2_X1 U539 ( .A(KEYINPUT16), .B(KEYINPUT84), .ZN(n474) );
  XNOR2_X1 U540 ( .A(n474), .B(KEYINPUT83), .ZN(n475) );
  XNOR2_X1 U541 ( .A(n476), .B(n475), .ZN(n479) );
  INV_X1 U542 ( .A(n477), .ZN(n478) );
  NAND2_X1 U543 ( .A1(n479), .A2(n478), .ZN(n499) );
  NOR2_X1 U544 ( .A1(n480), .A2(n499), .ZN(n487) );
  NAND2_X1 U545 ( .A1(n487), .A2(n511), .ZN(n481) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n487), .A2(n513), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U551 ( .A1(n487), .A2(n563), .ZN(n485) );
  XNOR2_X1 U552 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U553 ( .A1(n487), .A2(n518), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U555 ( .A1(n489), .A2(n495), .ZN(n492) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT100), .ZN(n490) );
  XNOR2_X1 U557 ( .A(n490), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U558 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n493), .A2(n495), .ZN(n494) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  NOR2_X1 U561 ( .A1(n496), .A2(n495), .ZN(n497) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n497), .Z(G1331GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n501) );
  NAND2_X1 U564 ( .A1(n498), .A2(n562), .ZN(n509) );
  NOR2_X1 U565 ( .A1(n509), .A2(n499), .ZN(n505) );
  NAND2_X1 U566 ( .A1(n505), .A2(n511), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U568 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NAND2_X1 U569 ( .A1(n505), .A2(n513), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n503), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n563), .A2(n505), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U574 ( .A1(n505), .A2(n518), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U576 ( .A(G78GAT), .B(n508), .Z(G1335GAT) );
  NOR2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n519) );
  NAND2_X1 U578 ( .A1(n519), .A2(n511), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(KEYINPUT106), .ZN(n515) );
  NAND2_X1 U581 ( .A1(n513), .A2(n519), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT107), .Z(n517) );
  NAND2_X1 U584 ( .A1(n519), .A2(n563), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(G1338GAT) );
  XNOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n523) );
  XOR2_X1 U587 ( .A(G106GAT), .B(KEYINPUT108), .Z(n521) );
  NAND2_X1 U588 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n539), .A2(n524), .ZN(n525) );
  NAND2_X1 U592 ( .A1(n525), .A2(n563), .ZN(n529) );
  NOR2_X1 U593 ( .A1(n526), .A2(n529), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1340GAT) );
  INV_X1 U596 ( .A(n529), .ZN(n535) );
  AND2_X1 U597 ( .A1(n562), .A2(n535), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n533) );
  NAND2_X1 U601 ( .A1(n535), .A2(n570), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U603 ( .A(G127GAT), .B(n534), .Z(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U605 ( .A1(n535), .A2(n572), .ZN(n536) );
  XNOR2_X1 U606 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U607 ( .A(G134GAT), .B(n538), .Z(G1343GAT) );
  XOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT119), .Z(n545) );
  NOR2_X1 U609 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(n543), .Z(n552) );
  NAND2_X1 U612 ( .A1(n552), .A2(n576), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n547) );
  NAND2_X1 U615 ( .A1(n552), .A2(n562), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n548), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n550) );
  NAND2_X1 U619 ( .A1(n586), .A2(n552), .ZN(n549) );
  XNOR2_X1 U620 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n552), .A2(n572), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n553), .B(KEYINPUT122), .ZN(n554) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  XOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT123), .Z(n561) );
  NOR2_X1 U626 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n557), .B(KEYINPUT55), .ZN(n564) );
  NOR2_X1 U628 ( .A1(n558), .A2(n564), .ZN(n573) );
  NAND2_X1 U629 ( .A1(n573), .A2(n559), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n563), .A2(n562), .ZN(n565) );
  OR2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n573), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1351GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n578) );
  NAND2_X1 U643 ( .A1(n587), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
endmodule

