//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT72), .B(G71gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G99gat), .ZN(new_n205));
  XOR2_X1   g004(.A(G15gat), .B(G43gat), .Z(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G227gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n211), .A2(KEYINPUT26), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n212), .A2(KEYINPUT26), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT64), .B(KEYINPUT28), .Z(new_n219));
  INV_X1    g018(.A(G183gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT27), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT27), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT28), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G190gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n221), .A3(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT65), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT27), .B(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(new_n227), .ZN(new_n232));
  AOI221_X4 g031(.A(new_n218), .B1(new_n219), .B2(new_n225), .C1(new_n229), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n232), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n225), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT66), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n217), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n212), .B(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n211), .B1(new_n242), .B2(new_n215), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n220), .A2(new_n224), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT24), .A3(new_n214), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(KEYINPUT67), .B(new_n217), .C1(new_n233), .C2(new_n236), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n239), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  OR2_X1    g050(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(KEYINPUT70), .A2(G113gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(G113gat), .A2(G120gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G127gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G134gat), .ZN(new_n259));
  INV_X1    g058(.A(G134gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G127gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n254), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n260), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(G127gat), .B(G134gat), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n267), .B2(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g067(.A1(G113gat), .A2(G120gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n255), .A2(new_n256), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n265), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n266), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT68), .ZN(new_n273));
  AND4_X1   g072(.A1(new_n265), .A2(new_n270), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n264), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n268), .A2(new_n265), .A3(new_n270), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n263), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT71), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n250), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n283), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n285), .A2(new_n248), .A3(new_n239), .A4(new_n249), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n208), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n207), .B1(new_n287), .B2(KEYINPUT33), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT32), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n284), .A2(new_n286), .A3(new_n208), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT34), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n284), .A2(new_n286), .ZN(new_n295));
  INV_X1    g094(.A(new_n208), .ZN(new_n296));
  AOI221_X4 g095(.A(new_n289), .B1(KEYINPUT33), .B2(new_n207), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n291), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n288), .A2(new_n290), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n293), .B1(new_n300), .B2(new_n297), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n203), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n300), .A2(new_n297), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT73), .B1(new_n303), .B2(new_n294), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n202), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n301), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT36), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g108(.A1(G197gat), .A2(G204gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(G197gat), .A2(G204gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT22), .ZN(new_n312));
  NAND2_X1  g111(.A1(G211gat), .A2(G218gat), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n310), .A2(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(KEYINPUT74), .A3(new_n315), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n250), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n325));
  INV_X1    g124(.A(new_n217), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n231), .B1(new_n230), .B2(new_n227), .ZN(new_n327));
  AND4_X1   g126(.A1(new_n231), .A2(new_n227), .A3(new_n221), .A4(new_n223), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n235), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n218), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n234), .A2(KEYINPUT66), .A3(new_n235), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n326), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n246), .B(KEYINPUT25), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n325), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n237), .A2(KEYINPUT75), .A3(new_n248), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n322), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n324), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n334), .A2(new_n335), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n323), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n323), .A2(KEYINPUT29), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n250), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n345), .A3(new_n321), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n324), .A2(new_n338), .A3(KEYINPUT76), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G8gat), .B(G36gat), .Z(new_n349));
  XNOR2_X1  g148(.A(G64gat), .B(G92gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT30), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n341), .A2(new_n346), .A3(new_n347), .A4(new_n353), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G57gat), .B(G85gat), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT86), .ZN(new_n360));
  XOR2_X1   g159(.A(G1gat), .B(G29gat), .Z(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G155gat), .B(G162gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G141gat), .B(G148gat), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(KEYINPUT2), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(KEYINPUT81), .A2(G148gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(KEYINPUT81), .A2(G148gat), .ZN(new_n370));
  INV_X1    g169(.A(G141gat), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G148gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(G141gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n365), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(KEYINPUT82), .A2(G155gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(KEYINPUT82), .A2(G155gat), .ZN(new_n377));
  OAI21_X1  g176(.A(G162gat), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n378), .A2(KEYINPUT2), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n368), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n281), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT5), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(KEYINPUT2), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n373), .ZN(new_n387));
  NAND2_X1  g186(.A1(KEYINPUT81), .A2(G148gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(G141gat), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n374), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n385), .A2(new_n391), .A3(new_n365), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n384), .B1(new_n392), .B2(new_n368), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n281), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n384), .A3(new_n368), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT83), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n397));
  AND4_X1   g196(.A1(KEYINPUT83), .A2(new_n397), .A3(new_n395), .A4(new_n275), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n382), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n380), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n277), .A2(new_n282), .A3(KEYINPUT4), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n281), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT84), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n401), .A2(new_n404), .ZN(new_n407));
  INV_X1    g206(.A(new_n382), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n394), .A2(KEYINPUT83), .A3(new_n395), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n397), .A2(new_n275), .A3(new_n395), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n408), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n407), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n383), .B1(new_n406), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n402), .A2(new_n403), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n277), .A2(new_n282), .A3(new_n400), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(new_n403), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n413), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n364), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT87), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n415), .ZN(new_n424));
  INV_X1    g223(.A(new_n383), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n364), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT6), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT87), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n429), .B(new_n364), .C1(new_n416), .C2(new_n421), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT6), .B(new_n364), .C1(new_n416), .C2(new_n421), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n357), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n347), .A2(new_n346), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n435), .A2(KEYINPUT79), .A3(new_n341), .A4(new_n353), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n436), .A3(new_n356), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n434), .A2(new_n436), .A3(KEYINPUT80), .A4(new_n356), .ZN(new_n440));
  AOI221_X4 g239(.A(new_n358), .B1(new_n431), .B2(new_n432), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(G22gat), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(KEYINPUT31), .B(G50gat), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n395), .A2(new_n336), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n321), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n319), .A2(new_n320), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n316), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n319), .A2(KEYINPUT89), .A3(new_n320), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT3), .B1(new_n455), .B2(new_n336), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n449), .B1(new_n456), .B2(new_n400), .ZN(new_n457));
  NAND2_X1  g256(.A1(G228gat), .A2(G233gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n458), .B(KEYINPUT88), .Z(new_n459));
  AOI21_X1  g258(.A(new_n447), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n447), .A3(new_n459), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n458), .B1(new_n448), .B2(new_n321), .ZN(new_n464));
  INV_X1    g263(.A(new_n321), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT3), .B1(new_n465), .B2(new_n336), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n466), .B2(new_n400), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n446), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n457), .A2(new_n447), .A3(new_n459), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n446), .B(new_n467), .C1(new_n469), .C2(new_n460), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n444), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n469), .B2(new_n460), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n445), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(new_n443), .A3(new_n470), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT91), .B1(new_n472), .B2(new_n475), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n309), .B1(new_n441), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT93), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n409), .A2(new_n412), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n419), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n408), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT92), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(KEYINPUT92), .A3(new_n408), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n490), .B1(new_n381), .B2(new_n382), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n487), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n427), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT40), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT40), .A4(new_n427), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n422), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n439), .A2(new_n440), .ZN(new_n499));
  INV_X1    g298(.A(new_n358), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n432), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n422), .B2(new_n428), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n354), .B1(new_n348), .B2(KEYINPUT37), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT37), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(new_n435), .B2(new_n341), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT38), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n434), .A2(new_n436), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n323), .A2(new_n342), .B1(new_n250), .B2(new_n344), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n505), .B1(new_n509), .B2(new_n465), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n465), .B1(new_n250), .B2(new_n323), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n338), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT38), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n513), .B(new_n354), .C1(new_n348), .C2(KEYINPUT37), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n503), .A2(new_n507), .A3(new_n508), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n476), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n482), .B1(new_n501), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n500), .ZN(new_n519));
  INV_X1    g318(.A(new_n498), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n515), .A2(new_n516), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(KEYINPUT93), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n481), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n358), .B1(new_n439), .B2(new_n440), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n431), .A2(new_n432), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n476), .A2(new_n306), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n474), .A2(new_n443), .A3(new_n470), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n443), .B1(new_n474), .B2(new_n470), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT35), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n428), .A2(new_n422), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n432), .ZN(new_n535));
  INV_X1    g334(.A(new_n304), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n530), .A2(new_n533), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT94), .B1(new_n537), .B2(new_n519), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n476), .A2(new_n503), .A3(KEYINPUT35), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n302), .A2(new_n304), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n539), .A2(new_n525), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n529), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n524), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n478), .A2(new_n479), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n525), .A2(new_n526), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n546), .A2(new_n547), .B1(new_n305), .B2(new_n308), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT93), .B1(new_n521), .B2(new_n522), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n501), .A2(new_n517), .A3(new_n482), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n529), .A2(new_n538), .A3(new_n542), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT95), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(G29gat), .A2(G36gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT14), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G29gat), .A2(G36gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G43gat), .B(G50gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(KEYINPUT15), .A3(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n558), .B(KEYINPUT96), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n562), .A2(new_n557), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT97), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT16), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(G1gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(G1gat), .B2(new_n570), .ZN(new_n573));
  INV_X1    g372(.A(G8gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n566), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(KEYINPUT17), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n569), .A2(new_n578), .B1(new_n576), .B2(new_n566), .ZN(new_n579));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT18), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT99), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n582), .ZN(new_n586));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587));
  INV_X1    g386(.A(G197gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT11), .B(G169gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT12), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n575), .B(new_n577), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n580), .B(KEYINPUT13), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n586), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n585), .A2(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n586), .A2(KEYINPUT98), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n586), .A2(KEYINPUT98), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n596), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n592), .B1(new_n601), .B2(new_n584), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n554), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n526), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT7), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(KEYINPUT8), .A2(new_n614), .B1(new_n608), .B2(new_n609), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G99gat), .B(G106gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n566), .ZN(new_n619));
  NAND3_X1  g418(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n619), .B(new_n620), .C1(KEYINPUT104), .C2(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n618), .B1(KEYINPUT17), .B2(new_n577), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n569), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(KEYINPUT104), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n630), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G71gat), .A2(G78gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(KEYINPUT9), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637));
  NOR2_X1   g436(.A1(G71gat), .A2(G78gat), .ZN(new_n638));
  OAI22_X1  g437(.A1(new_n636), .A2(new_n637), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G57gat), .B(G64gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(KEYINPUT21), .ZN(new_n643));
  XOR2_X1   g442(.A(G127gat), .B(G155gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n576), .B1(KEYINPUT21), .B2(new_n642), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  NAND2_X1  g446(.A1(G231gat), .A2(G233gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT101), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G183gat), .B(G211gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT102), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n651), .B(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n647), .A2(new_n654), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n633), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n618), .B(new_n642), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT10), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n642), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G120gat), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(G176gat), .B(G204gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  NAND3_X1  g469(.A1(new_n665), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n663), .A2(KEYINPUT105), .A3(new_n664), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n673), .A2(new_n674), .B1(new_n660), .B2(new_n666), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n671), .B1(new_n675), .B2(new_n670), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n607), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT106), .B(G1gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1324gat));
  NOR4_X1   g480(.A1(new_n554), .A2(new_n678), .A3(new_n604), .A4(new_n525), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT107), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT107), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n683), .B(new_n684), .C1(new_n685), .C2(G8gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT16), .B(G8gat), .ZN(new_n687));
  NOR2_X1   g486(.A1(KEYINPUT108), .A2(KEYINPUT42), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n682), .B2(new_n685), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n678), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n605), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n693), .B2(new_n309), .ZN(new_n694));
  INV_X1    g493(.A(new_n540), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(G15gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n693), .B2(new_n696), .ZN(G1326gat));
  NAND3_X1  g496(.A1(new_n605), .A2(new_n692), .A3(new_n546), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND3_X1  g499(.A1(new_n677), .A2(new_n658), .A3(new_n633), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n607), .A2(G29gat), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(KEYINPUT45), .ZN(new_n704));
  INV_X1    g503(.A(G29gat), .ZN(new_n705));
  INV_X1    g504(.A(new_n633), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n545), .B2(new_n553), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n524), .A2(new_n543), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n707), .B1(new_n710), .B2(new_n706), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n657), .B(KEYINPUT109), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n604), .A2(new_n714), .A3(new_n676), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n712), .A2(new_n526), .A3(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n717), .ZN(G1328gat));
  OAI21_X1  g517(.A(new_n544), .B1(new_n524), .B2(new_n543), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n551), .A2(KEYINPUT95), .A3(new_n552), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n701), .A2(G36gat), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n721), .A2(new_n603), .A3(new_n519), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT46), .ZN(new_n724));
  INV_X1    g523(.A(G36gat), .ZN(new_n725));
  INV_X1    g524(.A(new_n708), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n719), .B2(new_n720), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n551), .A2(new_n552), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n728), .B2(new_n633), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n727), .A2(new_n729), .A3(new_n716), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n725), .B1(new_n730), .B2(new_n519), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n724), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT110), .ZN(G1329gat));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  INV_X1    g533(.A(new_n309), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  OR3_X1    g535(.A1(new_n695), .A2(new_n701), .A3(G43gat), .ZN(new_n737));
  AOI211_X1 g536(.A(new_n604), .B(new_n737), .C1(new_n719), .C2(new_n720), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT112), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n738), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT47), .B1(new_n740), .B2(KEYINPUT111), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n709), .A2(new_n735), .A3(new_n711), .A4(new_n715), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(new_n744), .A3(new_n740), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n739), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n741), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n744), .B1(new_n743), .B2(new_n740), .ZN(new_n748));
  AOI211_X1 g547(.A(KEYINPUT112), .B(new_n738), .C1(new_n742), .C2(G43gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n746), .A2(new_n750), .ZN(G1330gat));
  NAND2_X1  g550(.A1(new_n730), .A2(new_n546), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G50gat), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n701), .A2(G50gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n721), .A2(new_n603), .A3(new_n546), .A4(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n709), .A2(new_n476), .A3(new_n711), .A4(new_n715), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G50gat), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n762), .A2(new_n755), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n759), .B(new_n760), .C1(new_n756), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n756), .B1(new_n762), .B2(new_n755), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n757), .B1(new_n752), .B2(G50gat), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT113), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(G1331gat));
  AND4_X1   g567(.A1(new_n659), .A2(new_n728), .A3(new_n676), .A4(new_n604), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n606), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT114), .B(G57gat), .Z(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1332gat));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n519), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT49), .B(G64gat), .Z(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(G1333gat));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n735), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n695), .A2(G71gat), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n777), .A2(G71gat), .B1(new_n769), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1334gat));
  NAND2_X1  g580(.A1(new_n769), .A2(new_n546), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n603), .A2(new_n657), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n676), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n712), .A2(new_n526), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n728), .A2(new_n633), .A3(new_n784), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT51), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n606), .A2(new_n608), .A3(new_n676), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n786), .A2(new_n608), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT116), .ZN(G1336gat));
  NOR2_X1   g590(.A1(new_n712), .A2(new_n785), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n609), .B1(new_n792), .B2(new_n519), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n519), .A2(new_n609), .A3(new_n676), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(KEYINPUT117), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(KEYINPUT117), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n788), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n793), .A2(new_n797), .A3(KEYINPUT52), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT52), .B1(new_n793), .B2(new_n797), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1337gat));
  NOR3_X1   g599(.A1(new_n712), .A2(new_n309), .A3(new_n785), .ZN(new_n801));
  INV_X1    g600(.A(G99gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n540), .A2(new_n802), .A3(new_n676), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n801), .A2(new_n802), .B1(new_n788), .B2(new_n803), .ZN(G1338gat));
  INV_X1    g603(.A(G106gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n792), .B2(new_n546), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n787), .B(KEYINPUT51), .Z(new_n807));
  NOR3_X1   g606(.A1(new_n516), .A2(new_n677), .A3(G106gat), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n805), .B1(new_n792), .B2(new_n476), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n810), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n813), .ZN(G1339gat));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n673), .A2(new_n815), .A3(new_n674), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n663), .B2(new_n664), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n661), .A2(new_n666), .A3(new_n662), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n670), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n671), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n603), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n816), .A2(new_n819), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n579), .A2(new_n580), .B1(new_n594), .B2(new_n595), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n585), .A2(new_n597), .B1(new_n591), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n676), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n633), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n827), .A2(new_n633), .A3(new_n830), .A4(new_n821), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n713), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n678), .B2(new_n603), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n606), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n837), .A2(new_n525), .A3(new_n527), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n838), .A2(new_n252), .A3(new_n253), .A4(new_n603), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n546), .A2(new_n695), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n525), .A2(new_n606), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n604), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n839), .A2(new_n845), .ZN(G1340gat));
  AOI21_X1  g645(.A(G120gat), .B1(new_n838), .B2(new_n676), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n677), .A2(new_n251), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n843), .B2(new_n848), .ZN(G1341gat));
  AND3_X1   g648(.A1(new_n838), .A2(new_n258), .A3(new_n657), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n258), .B1(new_n843), .B2(new_n714), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1342gat));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n260), .A3(new_n633), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n844), .B2(new_n706), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n857), .B(new_n858), .C1(new_n861), .C2(new_n862), .ZN(G1343gat));
  NOR2_X1   g662(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n836), .A2(new_n865), .A3(new_n476), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n735), .A2(new_n842), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT121), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n822), .A2(new_n825), .B1(new_n676), .B2(new_n830), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n833), .B1(new_n869), .B2(new_n633), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n870), .A2(new_n658), .B1(new_n692), .B2(new_n604), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT57), .B1(new_n871), .B2(new_n480), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n866), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n604), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n735), .A2(new_n516), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n603), .A2(new_n371), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT122), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n837), .A2(new_n525), .A3(new_n875), .A4(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n864), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g678(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n879), .B(new_n880), .ZN(G1344gat));
  NAND3_X1  g680(.A1(new_n836), .A2(KEYINPUT57), .A3(new_n476), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n865), .B1(new_n871), .B2(new_n480), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n676), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT59), .B(G148gat), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n837), .A2(new_n525), .A3(new_n875), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n676), .A2(new_n387), .A3(new_n388), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n873), .A2(new_n677), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n387), .B2(new_n388), .ZN(new_n893));
  OAI221_X1 g692(.A(new_n889), .B1(new_n890), .B2(new_n891), .C1(KEYINPUT59), .C2(new_n893), .ZN(G1345gat));
  OR2_X1    g693(.A1(new_n376), .A2(new_n377), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n873), .B2(new_n713), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n658), .A2(new_n895), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n890), .B2(new_n897), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n873), .B2(new_n706), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n706), .A2(G162gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n890), .B2(new_n900), .ZN(G1347gat));
  AND2_X1   g700(.A1(new_n836), .A2(new_n526), .ZN(new_n902));
  INV_X1    g701(.A(new_n527), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT125), .B1(new_n903), .B2(new_n525), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n903), .A2(new_n525), .A3(KEYINPUT125), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n603), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n525), .A2(new_n606), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n836), .A2(new_n840), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n604), .A2(new_n209), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(G1348gat));
  XNOR2_X1  g712(.A(new_n909), .B(KEYINPUT126), .ZN(new_n914));
  OAI21_X1  g713(.A(G176gat), .B1(new_n914), .B2(new_n677), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n906), .A2(new_n210), .A3(new_n676), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1349gat));
  OAI21_X1  g716(.A(G183gat), .B1(new_n914), .B2(new_n713), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n906), .A2(new_n657), .A3(new_n230), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT60), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n224), .A3(new_n633), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n633), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(G190gat), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT61), .B(new_n224), .C1(new_n911), .C2(new_n633), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(G1351gat));
  INV_X1    g729(.A(new_n908), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n931), .A2(new_n735), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(new_n884), .B2(new_n886), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n933), .A2(new_n588), .A3(new_n604), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n902), .A2(new_n519), .A3(new_n875), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n603), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n934), .A2(new_n936), .ZN(G1352gat));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n938));
  AOI21_X1  g737(.A(G204gat), .B1(new_n938), .B2(KEYINPUT62), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n676), .A3(new_n939), .ZN(new_n940));
  OR3_X1    g739(.A1(new_n940), .A2(new_n938), .A3(KEYINPUT62), .ZN(new_n941));
  OAI21_X1  g740(.A(G204gat), .B1(new_n933), .B2(new_n677), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n938), .B2(KEYINPUT62), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G1353gat));
  INV_X1    g743(.A(G211gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n935), .A2(new_n945), .A3(new_n657), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n657), .B(new_n932), .C1(new_n884), .C2(new_n886), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n947), .B2(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(G1354gat));
  OAI21_X1  g749(.A(G218gat), .B1(new_n933), .B2(new_n706), .ZN(new_n951));
  INV_X1    g750(.A(G218gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n952), .A3(new_n633), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1355gat));
endmodule


