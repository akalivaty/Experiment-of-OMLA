//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n621, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G2104), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(G137), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n469), .A2(new_n465), .A3(G125), .ZN(new_n470));
  AND2_X1   g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n463), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n477));
  AND4_X1   g052(.A1(KEYINPUT68), .A2(new_n462), .A3(new_n464), .A4(new_n465), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n467), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  MUX2_X1   g058(.A(G100), .B(G112), .S(G2105), .Z(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2104), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n462), .A2(new_n464), .A3(new_n467), .A4(new_n465), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n469), .A2(new_n465), .A3(G138), .A4(new_n467), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n492));
  NOR2_X1   g067(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G102), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2104), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n499), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n503));
  AND2_X1   g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n502), .A2(new_n503), .B1(new_n466), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n508), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(new_n509), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT71), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n517), .B2(new_n509), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(G651), .B1(G50), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n522), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n527), .A2(G51), .B1(new_n519), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n516), .A2(G89), .A3(new_n520), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT72), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n534), .A2(KEYINPUT72), .A3(new_n536), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n533), .B1(new_n538), .B2(new_n539), .ZN(G168));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n515), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(new_n545), .B2(new_n544), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n521), .A2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n527), .A2(G52), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(new_n521), .A2(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n515), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G651), .B1(G43), .B2(new_n527), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n527), .A2(G53), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n527), .B(G53), .C1(new_n566), .C2(new_n567), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n515), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n569), .A2(new_n570), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n516), .A2(G91), .A3(new_n520), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n574), .A2(KEYINPUT75), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT75), .B1(new_n574), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(new_n539), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n532), .B1(new_n579), .B2(new_n537), .ZN(G286));
  OR2_X1    g155(.A1(new_n519), .A2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n527), .B2(G49), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n516), .A2(new_n520), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(G288));
  AND3_X1   g160(.A1(new_n516), .A2(G86), .A3(new_n520), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n527), .A2(G48), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(new_n541), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n527), .A2(G47), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n583), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT76), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n541), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(KEYINPUT77), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G290));
  NAND3_X1  g177(.A1(new_n521), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n583), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n515), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g189(.A(new_n613), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  XOR2_X1   g191(.A(G299), .B(KEYINPUT78), .Z(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  XOR2_X1   g193(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g194(.A(G860), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n612), .B1(G559), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT80), .ZN(G148));
  OR2_X1    g197(.A1(new_n612), .A2(G559), .ZN(new_n623));
  MUX2_X1   g198(.A(new_n557), .B(new_n623), .S(G868), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  MUX2_X1   g200(.A(G99), .B(G111), .S(G2105), .Z(new_n626));
  AOI22_X1  g201(.A1(new_n482), .A2(G123), .B1(G2104), .B2(new_n626), .ZN(new_n627));
  AND3_X1   g202(.A1(new_n480), .A2(KEYINPUT81), .A3(G135), .ZN(new_n628));
  AOI21_X1  g203(.A(KEYINPUT81), .B1(new_n480), .B2(G135), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(G2096), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT82), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT84), .Z(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n640), .B2(new_n641), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT85), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n647), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n656), .A3(G14), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT86), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT17), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n663), .B1(new_n660), .B2(new_n662), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n661), .B2(new_n662), .ZN(new_n666));
  INV_X1    g241(.A(new_n662), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n667), .A2(new_n663), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n664), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT87), .Z(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  MUX2_X1   g270(.A(G24), .B(G290), .S(G16), .Z(new_n696));
  INV_X1    g271(.A(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G22), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G166), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT91), .B(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G6), .A2(G16), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n590), .B2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(G288), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT33), .B(G1976), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n702), .A2(new_n706), .A3(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n482), .A2(G119), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT90), .B1(G95), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NOR3_X1   g293(.A1(KEYINPUT90), .A2(G95), .A3(G2105), .ZN(new_n719));
  OAI221_X1 g294(.A(G2104), .B1(G107), .B2(new_n467), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n480), .A2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n698), .A2(new_n714), .A3(new_n715), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT36), .ZN(new_n728));
  NOR2_X1   g303(.A1(G27), .A2(G29), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G164), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2078), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n482), .A2(G129), .ZN(new_n732));
  NAND3_X1  g307(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT26), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n735), .A2(new_n736), .B1(G105), .B2(new_n473), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n480), .A2(G141), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n742), .B2(G32), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n731), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n707), .A2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G168), .B2(new_n707), .ZN(new_n748));
  INV_X1    g323(.A(G1966), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2090), .ZN(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G35), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G162), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT29), .Z(new_n754));
  OAI211_X1 g329(.A(new_n746), .B(new_n750), .C1(new_n751), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n480), .A2(G139), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n469), .A2(new_n465), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n757), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  AOI21_X1  g333(.A(KEYINPUT25), .B1(new_n473), .B2(G103), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n473), .A2(KEYINPUT25), .A3(G103), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n756), .B1(new_n467), .B2(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G33), .B(new_n761), .S(G29), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2072), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n755), .B(new_n764), .C1(new_n751), .C2(new_n754), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n742), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT94), .B1(G104), .B2(G2105), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g344(.A1(KEYINPUT94), .A2(G104), .A3(G2105), .ZN(new_n770));
  OAI221_X1 g345(.A(G2104), .B1(G116), .B2(new_n467), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n482), .A2(KEYINPUT93), .A3(G128), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(KEYINPUT93), .B1(new_n482), .B2(G128), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n477), .A2(new_n478), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(new_n467), .ZN(new_n778));
  INV_X1    g353(.A(G140), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n480), .A2(KEYINPUT92), .A3(G140), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n767), .B1(new_n783), .B2(new_n742), .ZN(new_n784));
  INV_X1    g359(.A(G2067), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G4), .A2(G16), .ZN(new_n787));
  INV_X1    g362(.A(new_n612), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1348), .Z(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n744), .B2(new_n745), .ZN(new_n791));
  NAND2_X1  g366(.A1(G299), .A2(G16), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n707), .A2(G20), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT23), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1956), .ZN(new_n796));
  NOR2_X1   g371(.A1(G16), .A2(G19), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n558), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1341), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n707), .A2(G5), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G171), .B2(new_n707), .ZN(new_n801));
  INV_X1    g376(.A(G1961), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT31), .B(G11), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT97), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT30), .B(G28), .Z(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(G29), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT24), .B(G34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(new_n742), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n475), .B2(new_n742), .ZN(new_n812));
  INV_X1    g387(.A(G2084), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n808), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI221_X1 g389(.A(new_n814), .B1(new_n813), .B2(new_n812), .C1(new_n630), .C2(new_n742), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n791), .A2(new_n796), .A3(new_n804), .A4(new_n815), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n728), .A2(new_n765), .A3(new_n786), .A4(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  NAND2_X1  g393(.A1(new_n527), .A2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  OAI221_X1 g396(.A(new_n819), .B1(new_n541), .B2(new_n820), .C1(new_n583), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  XOR2_X1   g399(.A(new_n557), .B(new_n822), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n788), .A2(G559), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n825), .B(new_n826), .Z(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT99), .Z(new_n832));
  OAI21_X1  g407(.A(new_n620), .B1(new_n830), .B2(KEYINPUT39), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n824), .B1(new_n832), .B2(new_n833), .ZN(G145));
  INV_X1    g409(.A(G37), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n506), .B1(new_n775), .B2(new_n782), .ZN(new_n836));
  INV_X1    g411(.A(new_n771), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n777), .A2(G2105), .ZN(new_n839));
  INV_X1    g414(.A(G128), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n837), .B1(new_n841), .B2(new_n772), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n780), .A2(new_n781), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(G164), .A3(new_n843), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n836), .A2(new_n740), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n740), .B1(new_n836), .B2(new_n844), .ZN(new_n846));
  OAI211_X1 g421(.A(KEYINPUT100), .B(new_n761), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n836), .A2(new_n844), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n741), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n836), .A2(new_n740), .A3(new_n844), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n761), .A2(KEYINPUT100), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n761), .A2(KEYINPUT100), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n634), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n723), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n480), .A2(G142), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n482), .A2(G130), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT101), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(KEYINPUT101), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n859), .B(new_n860), .C1(G118), .C2(new_n467), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n721), .A2(new_n634), .A3(new_n722), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n855), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n855), .B2(new_n863), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n847), .A2(new_n853), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n486), .B(G160), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n630), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n847), .A2(new_n853), .ZN(new_n871));
  INV_X1    g446(.A(new_n866), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT102), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n874));
  AOI211_X1 g449(.A(new_n874), .B(new_n866), .C1(new_n847), .C2(new_n853), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n870), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n872), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n874), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n871), .A2(KEYINPUT102), .A3(new_n872), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n867), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n847), .A2(new_n853), .A3(KEYINPUT103), .A4(new_n866), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n878), .A2(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n835), .B(new_n876), .C1(new_n883), .C2(new_n869), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g460(.A1(new_n822), .A2(G868), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n709), .B1(new_n600), .B2(new_n601), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n600), .A2(new_n709), .A3(new_n601), .ZN(new_n889));
  XNOR2_X1  g464(.A(G305), .B(G303), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n888), .B2(new_n889), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT42), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT104), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n892), .A2(new_n893), .ZN(new_n897));
  XOR2_X1   g472(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT106), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n788), .B1(new_n577), .B2(new_n576), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(G299), .A2(new_n612), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n902), .B2(new_n904), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n901), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n825), .B(new_n623), .ZN(new_n911));
  MUX2_X1   g486(.A(new_n905), .B(new_n910), .S(new_n911), .Z(new_n912));
  OR3_X1    g487(.A1(new_n896), .A2(new_n900), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n896), .B2(new_n900), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n886), .B1(new_n915), .B2(G868), .ZN(G295));
  AOI21_X1  g491(.A(new_n886), .B1(new_n915), .B2(G868), .ZN(G331));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n918));
  XNOR2_X1  g493(.A(G286), .B(G171), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n825), .ZN(new_n920));
  INV_X1    g495(.A(new_n825), .ZN(new_n921));
  XNOR2_X1  g496(.A(G286), .B(G301), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n907), .A3(new_n908), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n905), .A2(new_n923), .A3(new_n920), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n918), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n897), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n835), .B1(new_n897), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n925), .A2(new_n926), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT107), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n894), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n928), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT44), .B1(new_n938), .B2(new_n935), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n937), .B(new_n939), .ZN(G397));
  INV_X1    g515(.A(KEYINPUT126), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n491), .A2(new_n494), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT67), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(G138), .A3(new_n467), .A4(new_n464), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n947), .B2(KEYINPUT4), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n464), .A3(new_n504), .ZN(new_n949));
  INV_X1    g524(.A(new_n503), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT69), .B1(new_n499), .B2(G2104), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n942), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(KEYINPUT109), .B(G40), .Z(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  AND4_X1   g532(.A1(new_n468), .A2(new_n472), .A3(new_n474), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n783), .A2(new_n785), .ZN(new_n961));
  OAI21_X1  g536(.A(G2067), .B1(new_n775), .B2(new_n782), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n740), .B(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n723), .B(new_n725), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(G290), .B(new_n697), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n960), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n955), .A2(new_n958), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n974), .B2(G2078), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n496), .B2(new_n505), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  AOI211_X1 g553(.A(new_n978), .B(G1384), .C1(new_n496), .C2(new_n505), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n958), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n802), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n974), .A2(new_n972), .A3(G2078), .ZN(new_n983));
  OAI21_X1  g558(.A(G171), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n976), .A2(new_n958), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n582), .B(G1976), .C1(new_n584), .C2(new_n583), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(G8), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT52), .ZN(new_n988));
  INV_X1    g563(.A(G8), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n976), .B2(new_n958), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT110), .B(G1976), .Z(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n986), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(KEYINPUT111), .A2(KEYINPUT49), .ZN(new_n994));
  NAND2_X1  g569(.A1(G73), .A2(G543), .ZN(new_n995));
  INV_X1    g570(.A(G61), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n515), .B2(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n997), .A2(G651), .B1(G48), .B2(new_n527), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n516), .A2(G86), .A3(new_n520), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(new_n998), .B2(new_n999), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n994), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(G1981), .B1(new_n586), .B2(new_n589), .ZN(new_n1005));
  INV_X1    g580(.A(new_n994), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1001), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n990), .A3(new_n1007), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n988), .A2(new_n993), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1971), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n974), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n751), .B(new_n958), .C1(new_n977), .C2(new_n979), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n989), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G303), .A2(G8), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1009), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n506), .B2(new_n942), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n954), .B(G1384), .C1(new_n496), .C2(new_n505), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1971), .B1(new_n1020), .B2(new_n958), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n953), .A2(new_n978), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1023));
  AOI211_X1 g598(.A(G2090), .B(new_n959), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1016), .B(G8), .C1(new_n1021), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n984), .A2(new_n1017), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT118), .B1(G168), .B2(new_n989), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n1029));
  NAND3_X1  g604(.A1(G286), .A2(new_n1029), .A3(G8), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(KEYINPUT119), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n974), .A2(new_n749), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n813), .B(new_n958), .C1(new_n977), .C2(new_n979), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1033), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n989), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1032), .B(new_n1031), .C1(new_n1041), .C2(new_n1038), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1027), .A2(new_n1045), .A3(KEYINPUT122), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT62), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT122), .B1(new_n1027), .B2(new_n1045), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1009), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G288), .A2(G1976), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1008), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n990), .B1(new_n1054), .B2(new_n1002), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT112), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1052), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1009), .B(new_n1061), .C1(new_n1013), .C2(new_n1016), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n989), .B(G286), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1014), .B(KEYINPUT55), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n959), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n751), .A2(new_n1068), .B1(new_n974), .B2(new_n1010), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1069), .B2(new_n989), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1061), .B1(new_n1070), .B2(new_n1009), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1070), .A2(new_n1063), .A3(new_n1025), .A4(new_n1009), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1073), .A2(new_n1064), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1060), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1017), .A2(new_n1026), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1047), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n976), .A2(new_n785), .A3(new_n958), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1068), .B2(G1348), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1079), .A2(KEYINPUT60), .A3(new_n612), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n1081));
  INV_X1    g656(.A(new_n974), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G2072), .ZN(new_n1083));
  INV_X1    g658(.A(G1956), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1082), .A2(new_n1083), .B1(new_n980), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n569), .A2(new_n570), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n573), .A2(G651), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(new_n575), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT115), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n574), .A2(new_n1092), .A3(new_n575), .A4(new_n1089), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1088), .A2(KEYINPUT114), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1095), .A3(new_n1093), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1081), .B1(new_n1085), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n955), .A2(new_n958), .A3(new_n973), .A4(new_n1083), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1068), .B2(G1956), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1080), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1079), .A2(new_n788), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1078), .B(new_n612), .C1(new_n1068), .C2(G1348), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n955), .A2(new_n964), .A3(new_n958), .A4(new_n973), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT58), .B(G1341), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT116), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n985), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n558), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1116), .A3(new_n558), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1108), .A2(KEYINPUT60), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1104), .A2(KEYINPUT117), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1102), .A2(new_n1103), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1119), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1105), .B(new_n1118), .C1(new_n1123), .C2(KEYINPUT61), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1119), .A2(new_n1106), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1103), .B2(new_n1102), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1077), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n982), .A2(G171), .ZN(new_n1128));
  INV_X1    g703(.A(G2078), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1129), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1020), .A2(G160), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n984), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n975), .A2(new_n981), .A3(new_n1131), .A4(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n975), .A2(new_n981), .A3(new_n1131), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT120), .ZN(new_n1139));
  INV_X1    g714(.A(new_n983), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1137), .A2(new_n1139), .B1(new_n1140), .B2(new_n1128), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1134), .B1(new_n1141), .B2(new_n1133), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1075), .B1(new_n1127), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1051), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1077), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1075), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT121), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n971), .B1(new_n1145), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n963), .A2(new_n965), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT123), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n961), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n960), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n967), .A2(new_n960), .ZN(new_n1158));
  NOR2_X1   g733(.A1(G290), .A2(G1986), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n960), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT124), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1162), .A3(new_n960), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(KEYINPUT48), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT48), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1157), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n961), .A2(new_n962), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n960), .B1(new_n1168), .B2(new_n740), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n960), .A2(new_n964), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT46), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT47), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT125), .B1(new_n1167), .B2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1172), .B(KEYINPUT47), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1166), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1177), .A2(new_n1158), .A3(new_n1164), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .A4(new_n1157), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n941), .B1(new_n1152), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1148), .A2(new_n1144), .A3(new_n1149), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1051), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n970), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1187), .A2(KEYINPUT126), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1182), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g765(.A1(new_n694), .A2(new_n657), .A3(G319), .A4(new_n674), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1192), .B1(new_n931), .B2(new_n936), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n878), .A2(new_n879), .ZN(new_n1194));
  NAND2_X1  g768(.A1(new_n881), .A2(new_n882), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n869), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n876), .A2(new_n835), .ZN(new_n1197));
  OAI211_X1 g771(.A(new_n1193), .B(KEYINPUT127), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g772(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g773(.A(KEYINPUT127), .B1(new_n884), .B2(new_n1193), .ZN(new_n1200));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1200), .ZN(G308));
  NAND2_X1  g775(.A1(new_n884), .A2(new_n1193), .ZN(G225));
endmodule


