//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(G58), .A2(G68), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n222), .A2(G50), .A3(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n204), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n209), .A2(new_n220), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n219), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n226), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n203), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G226), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G45), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n262), .A3(new_n253), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1698), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G222), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G77), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n270), .A2(new_n271), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n273), .B(new_n277), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n229), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n257), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n267), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n228), .A2(new_n229), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G150), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n204), .A2(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n204), .B1(new_n221), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n290), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n228), .A2(new_n299), .A3(new_n229), .A4(new_n289), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n204), .A2(G1), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(G50), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n299), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n296), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n298), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n288), .B(new_n307), .C1(G169), .C2(new_n286), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n293), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n310), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n294), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G77), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n313), .A2(new_n290), .B1(new_n314), .B2(new_n305), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n301), .A2(G77), .A3(new_n303), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n266), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n258), .A2(G244), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n272), .A2(G232), .ZN(new_n320));
  INV_X1    g0120(.A(G107), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n320), .B1(new_n321), .B2(new_n278), .C1(new_n212), .C2(new_n279), .ZN(new_n322));
  AOI211_X1 g0122(.A(new_n318), .B(new_n319), .C1(new_n322), .C2(new_n285), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n317), .B1(new_n323), .B2(G190), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n323), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n287), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n327), .B(new_n317), .C1(G169), .C2(new_n323), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT9), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n286), .A2(G190), .B1(new_n307), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n286), .A2(new_n325), .B1(new_n330), .B2(new_n307), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT10), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n333), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT10), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n336), .A3(new_n331), .ZN(new_n337));
  AOI211_X1 g0137(.A(new_n309), .B(new_n329), .C1(new_n334), .C2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT13), .ZN(new_n339));
  INV_X1    g0139(.A(G226), .ZN(new_n340));
  INV_X1    g0140(.A(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n342), .B1(G232), .B2(new_n341), .C1(new_n274), .C2(new_n275), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G97), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(new_n285), .B1(KEYINPUT68), .B2(new_n266), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT68), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n318), .A2(new_n347), .B1(G238), .B2(new_n258), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n339), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(new_n348), .A3(new_n339), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G190), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n299), .A2(G68), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT12), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT11), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n291), .A2(G50), .B1(G20), .B2(new_n211), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n314), .B2(new_n294), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n290), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n301), .A2(G68), .A3(new_n303), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(new_n357), .C2(new_n360), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n325), .B1(new_n350), .B2(new_n351), .ZN(new_n364));
  OR3_X1    g0164(.A1(new_n354), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  INV_X1    g0166(.A(new_n351), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n366), .B(G169), .C1(new_n367), .C2(new_n349), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n287), .B2(new_n352), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n366), .B1(new_n352), .B2(G169), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n363), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n300), .A2(new_n310), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n299), .B1(new_n293), .B2(new_n302), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(KEYINPUT69), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT69), .B1(new_n375), .B2(new_n376), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT7), .B1(new_n276), .B2(new_n204), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  NOR4_X1   g0181(.A1(new_n274), .A2(new_n275), .A3(new_n381), .A4(G20), .ZN(new_n382));
  OAI21_X1  g0182(.A(G68), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G58), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n384), .A2(new_n211), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n385), .B2(new_n221), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n291), .A2(G159), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT16), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n270), .A2(new_n204), .A3(new_n271), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n381), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n211), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n386), .A2(KEYINPUT16), .A3(new_n387), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n290), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n379), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n280), .A2(new_n341), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n340), .A2(G1698), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n274), .C2(new_n275), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n284), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n256), .A2(new_n257), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(G232), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n266), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(G169), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n266), .A2(new_n405), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n401), .A2(new_n398), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n285), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n407), .B1(new_n411), .B2(new_n287), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n374), .B1(new_n397), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n397), .A2(new_n374), .A3(new_n412), .ZN(new_n415));
  INV_X1    g0215(.A(new_n290), .ZN(new_n416));
  INV_X1    g0216(.A(new_n395), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n383), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n394), .B2(new_n388), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n408), .A2(new_n410), .A3(new_n353), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n325), .B1(new_n402), .B2(new_n406), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(new_n424), .A3(new_n379), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n375), .A2(new_n376), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT69), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n375), .A2(KEYINPUT69), .A3(new_n376), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n420), .B2(new_n418), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(KEYINPUT17), .A3(new_n424), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n414), .A2(new_n415), .A3(new_n427), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n338), .A2(new_n373), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n278), .A2(G244), .A3(G1698), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G33), .A2(G116), .ZN(new_n439));
  OAI211_X1 g0239(.A(G238), .B(new_n341), .C1(new_n274), .C2(new_n275), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n285), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n254), .A2(new_n264), .A3(G1), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n254), .A2(G1), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n214), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n444), .A2(new_n445), .B1(new_n403), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(G190), .A3(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(KEYINPUT72), .A2(G87), .ZN(new_n450));
  NOR2_X1   g0250(.A1(G97), .A2(G107), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT72), .A2(G87), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT19), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n204), .B1(new_n344), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n278), .A2(new_n204), .A3(G68), .ZN(new_n457));
  INV_X1    g0257(.A(G97), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n454), .B1(new_n294), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n460), .A2(new_n290), .B1(new_n305), .B2(new_n312), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n300), .B1(new_n203), .B2(G33), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G87), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n325), .B1(new_n442), .B2(new_n448), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G169), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n442), .A2(new_n448), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n312), .B(KEYINPUT73), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n467), .A2(new_n468), .B1(new_n461), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n442), .A2(new_n287), .A3(new_n448), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n449), .A2(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  OAI211_X1 g0274(.A(G250), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(new_n341), .C1(new_n274), .C2(new_n275), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n474), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT4), .B1(new_n272), .B2(G244), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n285), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(G274), .A3(new_n446), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n481), .A2(new_n446), .B1(new_n256), .B2(new_n257), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(G257), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n480), .A2(new_n485), .A3(G179), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n467), .B1(new_n480), .B2(new_n485), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  AND2_X1   g0288(.A1(G97), .A2(G107), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(new_n451), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT70), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT6), .A2(G97), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(G107), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n321), .A2(KEYINPUT70), .A3(KEYINPUT6), .A4(G97), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(G20), .B1(G77), .B2(new_n291), .ZN(new_n496));
  OAI21_X1  g0296(.A(G107), .B1(new_n380), .B2(new_n382), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n416), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n305), .A2(new_n458), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n301), .B1(G1), .B2(new_n269), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n458), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n486), .A2(new_n487), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n498), .A2(new_n501), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n480), .A2(new_n485), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G200), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n480), .A2(new_n485), .A3(G190), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n204), .B(G87), .C1(new_n274), .C2(new_n275), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT22), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n278), .A2(new_n510), .A3(new_n204), .A4(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n439), .A2(G20), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT23), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n204), .B2(G107), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n321), .A2(KEYINPUT23), .A3(G20), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n512), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n513), .B1(new_n512), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n290), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT25), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n299), .B2(G107), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n305), .A2(KEYINPUT25), .A3(new_n321), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n462), .A2(G107), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G257), .B(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n526));
  OAI211_X1 g0326(.A(G250), .B(new_n341), .C1(new_n274), .C2(new_n275), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G294), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(new_n285), .B1(new_n484), .B2(G264), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n530), .A2(new_n353), .A3(new_n482), .ZN(new_n531));
  AOI21_X1  g0331(.A(G200), .B1(new_n530), .B2(new_n482), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n521), .B(new_n525), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n473), .A2(new_n502), .A3(new_n507), .A4(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G13), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(G1), .ZN(new_n536));
  INV_X1    g0336(.A(G116), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(G20), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(G20), .B1(G33), .B2(G283), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n269), .A2(G97), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n539), .A2(new_n540), .B1(G20), .B2(new_n537), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n541), .A2(new_n290), .A3(KEYINPUT20), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT20), .B1(new_n541), .B2(new_n290), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n538), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT74), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n500), .B2(new_n537), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n462), .A2(KEYINPUT74), .A3(G116), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT21), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n483), .B1(G270), .B2(new_n484), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n278), .A2(G264), .A3(G1698), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n278), .A2(G257), .A3(new_n341), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n276), .A2(G303), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n285), .ZN(new_n556));
  AOI211_X1 g0356(.A(new_n550), .B(new_n467), .C1(new_n551), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n551), .A2(new_n556), .A3(G179), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n549), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n551), .A2(new_n556), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G169), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n550), .B1(new_n548), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n521), .A2(new_n525), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n530), .A2(new_n482), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n467), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(G179), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n561), .A2(new_n353), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(G200), .B2(new_n561), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n548), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n437), .A2(new_n534), .A3(new_n574), .ZN(G372));
  AOI21_X1  g0375(.A(KEYINPUT77), .B1(new_n334), .B2(new_n337), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n334), .A2(KEYINPUT77), .A3(new_n337), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n434), .A2(new_n427), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n365), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n371), .B2(new_n328), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n397), .A2(new_n374), .A3(new_n412), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n413), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n579), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n586), .A2(new_n308), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n468), .A2(new_n467), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n461), .A2(new_n470), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(new_n472), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT75), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n468), .A2(G200), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n592), .A2(new_n461), .A3(new_n449), .A4(new_n463), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n521), .A2(new_n525), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n531), .A2(new_n532), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n593), .B(new_n590), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n502), .A2(new_n507), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n560), .B(new_n563), .C1(new_n565), .C2(new_n568), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n591), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n502), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n473), .A2(KEYINPUT26), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT76), .B1(new_n486), .B2(new_n487), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n504), .A2(G169), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT76), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n480), .A2(new_n485), .A3(G179), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n503), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n603), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n593), .A2(new_n590), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n602), .B1(new_n611), .B2(KEYINPUT26), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n600), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n587), .B1(new_n437), .B2(new_n614), .ZN(G369));
  NAND2_X1  g0415(.A1(new_n536), .A2(new_n204), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n616), .A2(KEYINPUT27), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(KEYINPUT27), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(G213), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(G343), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n548), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n564), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n573), .ZN(new_n625));
  INV_X1    g0425(.A(G330), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n533), .B1(new_n565), .B2(new_n622), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n594), .B(new_n567), .C1(G179), .C2(new_n566), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n569), .A2(new_n622), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT78), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT78), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n631), .A2(new_n635), .A3(new_n632), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n628), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n564), .A2(new_n622), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n634), .B2(new_n636), .ZN(new_n641));
  INV_X1    g0441(.A(new_n632), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n639), .A2(new_n643), .ZN(G399));
  INV_X1    g0444(.A(new_n207), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(G41), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n453), .A2(G116), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G1), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n224), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT28), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n473), .A2(new_n652), .A3(new_n601), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n600), .B(new_n653), .C1(new_n652), .C2(new_n611), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(KEYINPUT29), .A3(new_n622), .ZN(new_n655));
  XOR2_X1   g0455(.A(new_n655), .B(KEYINPUT82), .Z(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT79), .B1(new_n614), .B2(new_n621), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT79), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n613), .A2(new_n658), .A3(new_n622), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(KEYINPUT80), .B(KEYINPUT29), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT81), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT81), .ZN(new_n664));
  AOI211_X1 g0464(.A(new_n664), .B(new_n661), .C1(new_n657), .C2(new_n659), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n656), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n570), .A2(new_n598), .A3(new_n573), .A4(new_n622), .ZN(new_n667));
  INV_X1    g0467(.A(new_n530), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n468), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n559), .A2(new_n669), .A3(new_n480), .A4(new_n485), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT30), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n561), .A2(new_n287), .A3(new_n468), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n504), .A2(new_n566), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n670), .A2(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR4_X1   g0474(.A1(new_n558), .A2(new_n504), .A3(new_n468), .A4(new_n668), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT30), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n622), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT31), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n667), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n677), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT31), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n626), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n666), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n651), .B1(new_n686), .B2(G1), .ZN(G364));
  NOR2_X1   g0487(.A1(new_n535), .A2(G20), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n203), .B1(new_n688), .B2(G45), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n646), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n625), .A2(new_n626), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n628), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT83), .Z(new_n695));
  NOR2_X1   g0495(.A1(G13), .A2(G33), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G20), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n625), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n645), .A2(new_n278), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n260), .A2(new_n262), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n225), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n254), .B2(new_n251), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n645), .A2(new_n276), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n705), .A2(G355), .B1(new_n537), .B2(new_n645), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n231), .B1(G20), .B2(new_n467), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n698), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n692), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n708), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n204), .A2(new_n287), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT84), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(KEYINPUT84), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n325), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n353), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n287), .A2(new_n325), .A3(KEYINPUT85), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT85), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(G179), .B2(G200), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n353), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n204), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n716), .A2(G322), .B1(G294), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G311), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n715), .A2(G190), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n723), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n712), .A2(G200), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G190), .ZN(new_n729));
  INV_X1    g0529(.A(G317), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT33), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n730), .A2(KEYINPUT33), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G303), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n204), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G190), .A3(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n728), .A2(new_n353), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT87), .B(G326), .ZN(new_n739));
  OAI221_X1 g0539(.A(new_n733), .B1(new_n734), .B2(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n717), .A2(new_n719), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n204), .A2(G190), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(G329), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n735), .A2(new_n353), .A3(G200), .ZN(new_n745));
  INV_X1    g0545(.A(G283), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n276), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR4_X1   g0547(.A1(new_n727), .A2(new_n740), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n729), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n749), .A2(new_n211), .B1(new_n738), .B2(new_n296), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n743), .A2(G159), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n716), .A2(G58), .B1(KEYINPUT32), .B2(new_n751), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n752), .B1(KEYINPUT32), .B2(new_n751), .C1(new_n458), .C2(new_n721), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n750), .B(new_n753), .C1(G77), .C2(new_n725), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n736), .B1(new_n450), .B2(new_n452), .ZN(new_n755));
  INV_X1    g0555(.A(new_n745), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n276), .B(new_n755), .C1(G107), .C2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT86), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n748), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n699), .B(new_n710), .C1(new_n711), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n695), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(G396));
  NAND2_X1  g0563(.A1(new_n317), .A2(new_n621), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n326), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n328), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n328), .A2(new_n621), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n697), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n745), .A2(new_n213), .B1(new_n736), .B2(new_n321), .ZN(new_n772));
  INV_X1    g0572(.A(new_n743), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n276), .B1(new_n749), .B2(new_n746), .C1(new_n773), .C2(new_n724), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n772), .B(new_n774), .C1(G303), .C2(new_n737), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n725), .A2(G116), .B1(G97), .B2(new_n722), .ZN(new_n776));
  INV_X1    g0576(.A(G294), .ZN(new_n777));
  INV_X1    g0577(.A(new_n716), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n775), .B(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n729), .A2(G150), .B1(new_n737), .B2(G137), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  INV_X1    g0581(.A(G143), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n780), .B1(new_n726), .B2(new_n781), .C1(new_n782), .C2(new_n778), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT34), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n278), .B1(new_n736), .B2(new_n296), .C1(new_n211), .C2(new_n745), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G132), .B2(new_n743), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n785), .B(new_n787), .C1(new_n384), .C2(new_n721), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n783), .A2(new_n784), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n779), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n708), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n711), .A2(new_n697), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT88), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n791), .B1(G77), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n691), .B1(new_n771), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n660), .A2(new_n769), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n326), .A2(new_n328), .A3(new_n622), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n591), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n570), .B2(new_n534), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n610), .A2(new_n652), .A3(new_n502), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n473), .A2(new_n608), .A3(new_n607), .A4(new_n603), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(new_n802), .B2(new_n652), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n798), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT89), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT89), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n613), .A2(new_n806), .A3(new_n798), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n796), .A2(new_n684), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n692), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n684), .B1(new_n796), .B2(new_n808), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n795), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT90), .Z(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G384));
  OR2_X1    g0614(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n815), .A2(G116), .A3(new_n232), .A4(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT36), .Z(new_n818));
  OR3_X1    g0618(.A1(new_n224), .A2(new_n314), .A3(new_n385), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n296), .A2(G68), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n203), .B(G13), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n437), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n656), .B(new_n823), .C1(new_n663), .C2(new_n665), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n587), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT96), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n363), .A2(new_n621), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n372), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n365), .A2(new_n371), .A3(new_n827), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT91), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n808), .B2(new_n768), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n806), .B1(new_n613), .B2(new_n798), .ZN(new_n834));
  AOI211_X1 g0634(.A(KEYINPUT89), .B(new_n797), .C1(new_n600), .C2(new_n612), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n832), .B(new_n768), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n831), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n428), .B1(new_n390), .B2(new_n396), .ZN(new_n840));
  INV_X1    g0640(.A(new_n619), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n433), .A2(new_n424), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n412), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n397), .A2(new_n412), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n619), .B(KEYINPUT92), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n397), .A2(new_n846), .ZN(new_n847));
  AND4_X1   g0647(.A1(new_n839), .A2(new_n845), .A3(new_n847), .A4(new_n425), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT93), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n424), .ZN(new_n850));
  INV_X1    g0650(.A(new_n428), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n418), .B2(new_n420), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n397), .A2(new_n850), .B1(new_n852), .B2(new_n619), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n840), .A2(new_n412), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT93), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n845), .A2(new_n847), .A3(new_n839), .A4(new_n425), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n852), .A2(new_n619), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n435), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n849), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n849), .A2(KEYINPUT38), .A3(new_n860), .A4(new_n858), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n838), .A2(new_n866), .B1(new_n584), .B2(new_n846), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n371), .A2(new_n621), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n863), .B2(new_n864), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n845), .A2(new_n847), .A3(new_n425), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(new_n839), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n847), .B1(new_n580), .B2(new_n584), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n862), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n864), .A2(new_n874), .A3(new_n869), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT94), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n870), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n855), .A2(new_n857), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n878), .A2(KEYINPUT93), .B1(new_n435), .B2(new_n859), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n879), .B2(new_n858), .ZN(new_n880));
  AND4_X1   g0680(.A1(KEYINPUT38), .A2(new_n849), .A3(new_n858), .A4(new_n860), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT39), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n882), .A2(KEYINPUT94), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT95), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n864), .A2(new_n874), .A3(new_n869), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(KEYINPUT94), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT95), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n870), .A2(new_n876), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n868), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n867), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n826), .B(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT97), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n680), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n681), .B1(new_n677), .B2(KEYINPUT97), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n678), .B(new_n667), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n769), .B1(new_n829), .B2(new_n830), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT40), .B1(new_n863), .B2(new_n864), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n864), .A2(new_n874), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT40), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n823), .A2(new_n896), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n626), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n892), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n203), .B2(new_n688), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n892), .A2(new_n907), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n822), .B1(new_n909), .B2(new_n910), .ZN(G367));
  AND2_X1   g0711(.A1(new_n700), .A2(new_n243), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n709), .B1(new_n207), .B2(new_n312), .ZN(new_n913));
  INV_X1    g0713(.A(new_n736), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT46), .B1(new_n914), .B2(G116), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n278), .B1(new_n729), .B2(G294), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n737), .A2(G311), .B1(new_n756), .B2(G97), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n916), .B(new_n917), .C1(new_n778), .C2(new_n734), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n726), .A2(new_n746), .B1(new_n321), .B2(new_n721), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n914), .A2(KEYINPUT46), .A3(G116), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n773), .B2(new_n730), .ZN(new_n921));
  OR4_X1    g0721(.A1(new_n915), .A2(new_n918), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n736), .A2(new_n384), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n749), .A2(new_n781), .B1(new_n738), .B2(new_n782), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n923), .B(new_n924), .C1(G137), .C2(new_n743), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n278), .B1(new_n745), .B2(new_n314), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n925), .B1(KEYINPUT104), .B2(new_n926), .C1(new_n211), .C2(new_n721), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n725), .A2(G50), .B1(KEYINPUT104), .B2(new_n926), .ZN(new_n928));
  INV_X1    g0728(.A(G150), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n929), .B2(new_n778), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n922), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT47), .Z(new_n932));
  OAI221_X1 g0732(.A(new_n691), .B1(new_n912), .B2(new_n913), .C1(new_n932), .C2(new_n711), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT105), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n464), .A2(new_n621), .ZN(new_n935));
  MUX2_X1   g0735(.A(new_n799), .B(new_n610), .S(new_n935), .Z(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n698), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT106), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n503), .A2(new_n622), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n609), .A2(new_n622), .B1(new_n597), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT98), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT101), .B1(new_n643), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT101), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n945), .B(new_n942), .C1(new_n641), .C2(new_n642), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n641), .A2(new_n642), .A3(new_n942), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT45), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n944), .A2(KEYINPUT44), .A3(new_n946), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n638), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT102), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n949), .A2(new_n639), .A3(new_n951), .A4(new_n952), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n953), .A2(KEYINPUT102), .A3(new_n638), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT103), .B1(new_n637), .B2(new_n640), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n628), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n634), .A2(new_n636), .ZN(new_n962));
  INV_X1    g0762(.A(new_n640), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n627), .B1(new_n964), .B2(KEYINPUT103), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n641), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n961), .A2(new_n641), .A3(new_n965), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n959), .A2(new_n686), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n686), .B1(new_n958), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n646), .B(KEYINPUT41), .Z(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n690), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n943), .A2(new_n641), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT42), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n502), .B1(new_n942), .B2(new_n630), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n622), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT43), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n936), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n981), .A2(KEYINPUT99), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n978), .A2(new_n983), .A3(new_n980), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT99), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n936), .B(new_n982), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n984), .B(new_n987), .C1(new_n981), .C2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT100), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n638), .A2(new_n943), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n990), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n939), .B1(new_n975), .B2(new_n996), .ZN(G387));
  INV_X1    g0797(.A(new_n240), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n700), .B1(new_n998), .B2(new_n702), .ZN(new_n999));
  INV_X1    g0799(.A(new_n705), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n648), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n310), .A2(KEYINPUT50), .A3(new_n296), .ZN(new_n1003));
  AOI21_X1  g0803(.A(KEYINPUT50), .B1(new_n310), .B2(new_n296), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n648), .B(new_n1002), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1001), .A2(new_n1005), .B1(new_n321), .B2(new_n645), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n709), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n691), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n729), .A2(G311), .B1(new_n737), .B2(G322), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n726), .B2(new_n734), .C1(new_n730), .C2(new_n778), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n722), .A2(G283), .B1(G294), .B2(new_n914), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT49), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n276), .B1(new_n537), .B2(new_n745), .C1(new_n773), .C2(new_n739), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n781), .A2(new_n738), .B1(new_n749), .B2(new_n293), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n278), .B1(new_n458), .B2(new_n745), .C1(new_n773), .C2(new_n929), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G77), .C2(new_n914), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n469), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(new_n721), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G50), .B2(new_n716), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1023), .B(new_n1026), .C1(new_n211), .C2(new_n726), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n711), .B1(new_n1020), .B2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1008), .B(new_n1028), .C1(new_n637), .C2(new_n698), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n970), .B2(new_n690), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n970), .A2(new_n666), .A3(new_n684), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(KEYINPUT107), .A3(new_n646), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n686), .B2(new_n970), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT107), .B1(new_n1031), .B2(new_n646), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(G393));
  INV_X1    g0835(.A(new_n971), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n957), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n955), .B2(new_n954), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n647), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT108), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n954), .A2(new_n1040), .A3(new_n957), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n953), .A2(KEYINPUT108), .A3(new_n638), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n1031), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n942), .A2(new_n698), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n716), .A2(G311), .B1(G317), .B2(new_n737), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT52), .Z(new_n1046));
  AOI22_X1  g0846(.A1(new_n722), .A2(G116), .B1(G303), .B2(new_n729), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n726), .B2(new_n777), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT111), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n276), .B1(new_n736), .B2(new_n746), .C1(new_n321), .C2(new_n745), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G322), .B2(new_n743), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1046), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT112), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n716), .A2(G159), .B1(G150), .B2(new_n737), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n276), .B1(new_n756), .B2(G87), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n211), .B2(new_n736), .C1(new_n749), .C2(new_n296), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G143), .B2(new_n743), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n725), .A2(new_n310), .B1(G77), .B2(new_n722), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1053), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1052), .A2(KEYINPUT112), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n708), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1007), .B1(G97), .B2(new_n645), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n701), .A2(new_n248), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n692), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1039), .A2(new_n1043), .B1(new_n1044), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT109), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n689), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(G390));
  NAND3_X1  g0875(.A1(new_n683), .A2(new_n770), .A3(new_n831), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT115), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n831), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n896), .A2(G330), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1079), .A2(KEYINPUT117), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n770), .B1(new_n1079), .B2(KEYINPUT117), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n654), .A2(new_n622), .A3(new_n766), .ZN(new_n1083));
  AND3_X1   g0883(.A1(new_n1083), .A2(KEYINPUT113), .A3(new_n768), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT113), .B1(new_n1083), .B2(new_n768), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1077), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1078), .B1(new_n684), .B2(new_n769), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n896), .A2(new_n897), .A3(G330), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT116), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n768), .B1(new_n834), .B2(new_n835), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(KEYINPUT91), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n836), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1090), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1091), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1087), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n823), .A2(new_n896), .A3(G330), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n824), .A2(new_n587), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n901), .A2(new_n868), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n1086), .B2(new_n1078), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n884), .A2(new_n889), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n868), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n1094), .B2(new_n831), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1104), .B(new_n1077), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1102), .B1(new_n1109), .B2(new_n831), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n838), .A2(new_n868), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(KEYINPUT114), .B(new_n1108), .C1(new_n1115), .C2(new_n1089), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1078), .B1(new_n1093), .B2(new_n836), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n884), .B(new_n889), .C1(new_n1117), .C2(new_n1106), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n1104), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT114), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1089), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1101), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(new_n647), .ZN(new_n1124));
  AOI211_X1 g0924(.A(KEYINPUT114), .B(new_n1089), .C1(new_n1118), .C2(new_n1104), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1120), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n1108), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT118), .B1(new_n1127), .B2(new_n1101), .ZN(new_n1128));
  AND4_X1   g0928(.A1(KEYINPUT118), .A2(new_n1116), .A3(new_n1122), .A4(new_n1101), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1127), .A2(new_n689), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1113), .A2(new_n696), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n793), .A2(new_n310), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n738), .A2(new_n746), .B1(new_n213), .B2(new_n736), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n278), .B(new_n1134), .C1(G68), .C2(new_n756), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n716), .A2(G116), .B1(G77), .B2(new_n722), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(new_n777), .C2(new_n773), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n725), .A2(G97), .B1(G107), .B2(new_n729), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT119), .Z(new_n1139));
  AOI22_X1  g0939(.A1(new_n729), .A2(G137), .B1(new_n737), .B2(G128), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n743), .A2(G125), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n276), .B1(new_n756), .B2(G50), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT54), .B(G143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G132), .A2(new_n716), .B1(new_n725), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n736), .A2(new_n929), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(new_n781), .C2(new_n721), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n1137), .A2(new_n1139), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n692), .B(new_n1133), .C1(new_n1150), .C2(new_n708), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1131), .B1(new_n1132), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1130), .A2(new_n1152), .ZN(G378));
  INV_X1    g0953(.A(KEYINPUT121), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n307), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n619), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n579), .B2(new_n308), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n309), .B(new_n1156), .C1(new_n577), .C2(new_n578), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT120), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n578), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n308), .B1(new_n1161), .B2(new_n576), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1156), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n579), .A2(new_n308), .A3(new_n1157), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT120), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  NAND3_X1  g0967(.A1(new_n1160), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1158), .A2(new_n1159), .A3(KEYINPUT120), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1165), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n898), .A2(new_n899), .B1(new_n902), .B2(KEYINPUT40), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1168), .B(new_n1172), .C1(new_n1173), .C2(new_n626), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1168), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n904), .A2(new_n1175), .A3(G330), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1177), .A2(new_n867), .A3(new_n890), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n584), .A2(new_n846), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1117), .B2(new_n865), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1179), .A2(new_n1181), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1154), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1177), .B1(new_n867), .B2(new_n890), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1179), .A2(new_n1181), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n1185), .A3(KEYINPUT121), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1123), .B2(new_n1099), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT57), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1123), .B2(new_n1099), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT122), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT122), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1194), .B(new_n1191), .C1(new_n1123), .C2(new_n1099), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1190), .A2(new_n1193), .A3(new_n646), .A4(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n691), .B1(new_n793), .B2(G50), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n721), .A2(new_n929), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n725), .A2(G137), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n729), .A2(G132), .B1(new_n737), .B2(G125), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n736), .C2(new_n1144), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1198), .B(new_n1201), .C1(G128), .C2(new_n716), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n269), .B(new_n253), .C1(new_n745), .C2(new_n781), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G124), .B2(new_n743), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n716), .A2(G107), .B1(G68), .B2(new_n722), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1024), .B2(new_n726), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n745), .A2(new_n384), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G116), .B2(new_n737), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n458), .B2(new_n749), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n773), .A2(new_n746), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n253), .B(new_n276), .C1(new_n736), .C2(new_n314), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n1210), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G50), .B1(new_n269), .B2(new_n253), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n278), .B2(G41), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1208), .A2(new_n1217), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1197), .B1(new_n1221), .B2(new_n708), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1175), .B2(new_n697), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1187), .B2(new_n690), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1196), .A2(new_n1225), .ZN(G375));
  NAND2_X1  g1026(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT116), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1090), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1099), .A3(new_n1087), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1101), .A2(new_n1231), .A3(new_n974), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT123), .Z(new_n1233));
  NAND2_X1  g1033(.A1(new_n1078), .A2(new_n696), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n691), .B1(new_n793), .B2(G68), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1025), .B1(G107), .B2(new_n725), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n746), .B2(new_n778), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n276), .B1(new_n745), .B2(new_n314), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G303), .B2(new_n743), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n729), .A2(G116), .B1(new_n737), .B2(G294), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1239), .B(new_n1240), .C1(new_n458), .C2(new_n736), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G137), .A2(new_n716), .B1(new_n725), .B2(G150), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n296), .B2(new_n721), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n276), .B(new_n1211), .C1(G128), .C2(new_n743), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n737), .A2(G132), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n729), .A2(new_n1145), .B1(new_n914), .B2(G159), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1237), .A2(new_n1241), .B1(new_n1243), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1235), .B1(new_n1248), .B2(new_n708), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1097), .A2(new_n690), .B1(new_n1234), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1233), .A2(new_n1250), .ZN(G381));
  NOR2_X1   g1051(.A1(G375), .A2(G378), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(G407));
  INV_X1    g1055(.A(G213), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(G343), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1252), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G407), .A2(G213), .A3(new_n1258), .ZN(G409));
  NAND3_X1  g1059(.A1(new_n1196), .A2(G378), .A3(new_n1225), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1224), .B1(new_n1261), .B2(new_n690), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1188), .B2(new_n973), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n1130), .A3(new_n1152), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1260), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1257), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1231), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1230), .A2(KEYINPUT60), .A3(new_n1099), .A4(new_n1087), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1269), .A2(new_n646), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1250), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(G384), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n813), .A3(new_n1250), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1265), .A2(new_n1266), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT62), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1271), .A2(new_n813), .A3(new_n1250), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n813), .B1(new_n1271), .B2(new_n1250), .ZN(new_n1280));
  INV_X1    g1080(.A(G2897), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n1279), .A2(new_n1280), .B1(new_n1281), .B2(new_n1266), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1266), .A2(new_n1281), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1273), .A2(new_n1274), .A3(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1278), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1257), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1275), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1277), .A2(new_n1286), .A3(new_n1287), .A4(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(G393), .B(new_n762), .ZN(new_n1292));
  AND2_X1   g1092(.A1(G387), .A2(G390), .ZN(new_n1293));
  OAI211_X1 g1093(.A(KEYINPUT126), .B(new_n1292), .C1(new_n1293), .C2(new_n1253), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n685), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n689), .B1(new_n1295), .B2(new_n973), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n994), .A2(new_n995), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1298), .A2(new_n939), .A3(new_n1074), .A4(new_n1070), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1292), .A2(KEYINPUT126), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G387), .A2(G390), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(G393), .B(G396), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .A4(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1294), .A2(KEYINPUT127), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT127), .B1(new_n1294), .B2(new_n1305), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1291), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1294), .A2(new_n1287), .A3(new_n1305), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1276), .B2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1288), .A2(KEYINPUT63), .A3(new_n1275), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1282), .A2(new_n1284), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(KEYINPUT124), .B2(new_n1288), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1288), .A2(KEYINPUT124), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1312), .B(new_n1313), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1309), .A2(new_n1320), .ZN(G405));
  NAND3_X1  g1121(.A1(G375), .A2(new_n1130), .A3(new_n1152), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1260), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1275), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1306), .A2(new_n1307), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1303), .B(new_n1302), .C1(new_n1299), .C2(new_n1301), .ZN(new_n1327));
  AND4_X1   g1127(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .A4(new_n1304), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1326), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1294), .A2(KEYINPUT127), .A3(new_n1305), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1275), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1323), .B1(new_n1325), .B2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1324), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1329), .A2(new_n1330), .A3(new_n1275), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1333), .A2(new_n1334), .A3(new_n1260), .A4(new_n1322), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1332), .A2(new_n1335), .ZN(G402));
endmodule


