//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT27), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT64), .B1(new_n193), .B2(G137), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  OAI211_X1 g011(.A(KEYINPUT64), .B(new_n197), .C1(new_n193), .C2(G137), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G137), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(KEYINPUT65), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n193), .A2(G137), .ZN(new_n205));
  OAI211_X1 g019(.A(G131), .B(new_n203), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n208), .B(new_n210), .C1(KEYINPUT1), .C2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT1), .B1(new_n209), .B2(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n209), .A2(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n207), .A2(G143), .ZN(new_n215));
  OAI211_X1 g029(.A(G128), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AND4_X1   g030(.A1(new_n200), .A2(new_n206), .A3(new_n212), .A4(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n195), .A2(new_n198), .A3(new_n199), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n200), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n208), .A2(new_n210), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G143), .B(G146), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT0), .B(G128), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT69), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n222), .B(new_n227), .C1(new_n223), .C2(new_n224), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n217), .B1(new_n220), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n231));
  INV_X1    g045(.A(G113), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT2), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G113), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n233), .A2(new_n235), .B1(new_n236), .B2(G119), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT67), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n241), .A3(G116), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n237), .A2(KEYINPUT68), .A3(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n236), .A2(G119), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n233), .A2(new_n235), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n245), .A2(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n230), .A2(new_n231), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n228), .ZN(new_n252));
  INV_X1    g066(.A(new_n221), .ZN(new_n253));
  OR2_X1    g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n253), .B(new_n254), .C1(new_n214), .C2(new_n215), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n227), .B1(new_n255), .B2(new_n222), .ZN(new_n256));
  AND4_X1   g070(.A1(new_n196), .A2(new_n195), .A3(new_n198), .A4(new_n199), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n202), .A2(G134), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n194), .B2(KEYINPUT11), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n196), .B1(new_n259), .B2(new_n198), .ZN(new_n260));
  OAI22_X1  g074(.A1(new_n252), .A2(new_n256), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n216), .A2(new_n212), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n200), .A3(new_n206), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n250), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n251), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n225), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n257), .B2(new_n260), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n263), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n248), .A2(new_n249), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n237), .A2(KEYINPUT68), .A3(new_n242), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT68), .B1(new_n237), .B2(new_n242), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n192), .B1(new_n266), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n225), .B1(new_n219), .B2(new_n200), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT66), .B(new_n277), .C1(new_n278), .C2(new_n217), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n261), .A2(KEYINPUT30), .A3(new_n263), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT66), .B1(new_n269), .B2(new_n277), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n281), .A2(new_n282), .A3(new_n250), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n264), .A2(new_n192), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n276), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n277), .B1(new_n278), .B2(new_n217), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n288), .A2(new_n273), .A3(new_n280), .A4(new_n279), .ZN(new_n289));
  INV_X1    g103(.A(new_n284), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(KEYINPUT31), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n275), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n187), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n187), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT70), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n230), .A2(new_n250), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n265), .B2(new_n251), .ZN(new_n300));
  INV_X1    g114(.A(new_n192), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(G902), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n266), .A2(new_n274), .A3(new_n192), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n302), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n192), .B1(new_n289), .B2(new_n264), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G472), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n289), .A2(KEYINPUT31), .A3(new_n290), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT31), .B1(new_n289), .B2(new_n290), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n266), .A2(new_n274), .ZN(new_n312));
  OAI22_X1  g126(.A1(new_n310), .A2(new_n311), .B1(new_n312), .B2(new_n192), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n296), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n295), .A2(new_n298), .A3(new_n309), .A4(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT22), .B(G137), .ZN(new_n317));
  INV_X1    g131(.A(G953), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(G221), .A3(G234), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n317), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT67), .B(G119), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(G128), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n238), .A2(new_n211), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n323), .B2(new_n211), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n326), .B2(new_n322), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G110), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT24), .B(G110), .Z(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT16), .ZN(new_n331));
  INV_X1    g145(.A(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(G125), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n333), .B1(new_n337), .B2(new_n331), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n207), .ZN(new_n339));
  OAI211_X1 g153(.A(G146), .B(new_n333), .C1(new_n337), .C2(new_n331), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n328), .A2(new_n330), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n334), .A2(new_n336), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(new_n207), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n337), .A2(KEYINPUT72), .A3(G146), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G110), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n324), .C1(new_n326), .C2(new_n322), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n326), .A2(new_n329), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n321), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n351), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n354), .B(new_n340), .C1(new_n347), .C2(new_n346), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n342), .A3(new_n320), .ZN(new_n356));
  INV_X1    g170(.A(G902), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT25), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n353), .A2(new_n356), .A3(new_n360), .A4(new_n357), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT71), .B(G217), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(G234), .B2(new_n357), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n359), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n353), .A2(new_n356), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n363), .A2(G902), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(KEYINPUT73), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n353), .A2(new_n356), .A3(new_n366), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n316), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G469), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT3), .A3(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT75), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n379), .B2(G104), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(KEYINPUT75), .A3(G107), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n381), .A2(new_n382), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n377), .A2(G107), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n379), .A2(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n386), .A2(new_n212), .A3(new_n216), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT10), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n262), .A2(new_n392), .A3(new_n386), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n257), .A2(new_n260), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n378), .A2(new_n380), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n384), .A2(new_n385), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT76), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n381), .A2(new_n399), .A3(new_n384), .A4(new_n385), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(G101), .A3(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n382), .A2(KEYINPUT4), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n229), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n394), .B(new_n395), .C1(new_n403), .C2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(G110), .B(G140), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n318), .A2(G227), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n386), .A2(new_n389), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n216), .A2(new_n212), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n390), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n416), .A2(KEYINPUT12), .A3(new_n220), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT12), .B1(new_n416), .B2(new_n220), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n412), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n394), .B1(new_n403), .B2(new_n406), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n220), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n411), .B1(new_n422), .B2(new_n407), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n375), .B(new_n357), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n407), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n410), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n407), .A2(new_n427), .A3(new_n411), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n422), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n427), .B1(new_n407), .B2(new_n411), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n426), .B(G469), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(G469), .A2(G902), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n424), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT9), .B(G234), .ZN(new_n434));
  OAI21_X1  g248(.A(G221), .B1(new_n434), .B2(G902), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT74), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n439), .B(KEYINPUT78), .Z(new_n440));
  OAI21_X1  g254(.A(G210), .B1(G237), .B2(G902), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n245), .A2(new_n246), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n386), .A2(new_n389), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n242), .A2(KEYINPUT5), .A3(new_n247), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n445), .B(G113), .C1(KEYINPUT5), .C2(new_n242), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G122), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n273), .A2(new_n405), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n447), .B(new_n448), .C1(new_n403), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n401), .A2(new_n402), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n273), .A3(new_n405), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT79), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n447), .A4(new_n448), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n448), .B1(new_n453), .B2(new_n447), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(KEYINPUT80), .B(KEYINPUT6), .Z(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT81), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n457), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n225), .A2(G125), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n414), .A2(new_n335), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n225), .A2(new_n469), .A3(G125), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G224), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G953), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n471), .B(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n460), .A2(new_n463), .A3(new_n465), .A4(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n451), .A2(new_n455), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n468), .A2(new_n466), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(new_n479), .B2(new_n473), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n473), .A2(new_n479), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n467), .A2(new_n468), .A3(new_n470), .A4(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n448), .B(KEYINPUT8), .Z(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n445), .ZN(new_n486));
  OAI21_X1  g300(.A(G113), .B1(new_n242), .B2(KEYINPUT5), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n271), .A2(new_n272), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(new_n413), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n444), .B1(new_n443), .B2(new_n446), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n413), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n484), .B1(new_n494), .B2(new_n447), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n480), .A2(new_n482), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT83), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(KEYINPUT84), .B(new_n357), .C1(new_n477), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n476), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n456), .A2(new_n497), .A3(new_n493), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT84), .B1(new_n501), .B2(new_n357), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n442), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n357), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT84), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n506), .A2(new_n441), .A3(new_n476), .A4(new_n499), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n440), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n211), .A2(G143), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n211), .A2(G143), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(KEYINPUT13), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT86), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n193), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n209), .A2(G128), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT13), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT86), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n513), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n510), .A3(new_n193), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT87), .ZN(new_n519));
  XNOR2_X1  g333(.A(G116), .B(G122), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(new_n379), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n379), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n523), .A2(KEYINPUT88), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n236), .A2(KEYINPUT14), .A3(G122), .ZN(new_n525));
  INV_X1    g339(.A(new_n520), .ZN(new_n526));
  OAI211_X1 g340(.A(G107), .B(new_n525), .C1(new_n526), .C2(KEYINPUT14), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n514), .A2(new_n510), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G134), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n518), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n523), .A2(KEYINPUT88), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n524), .A2(new_n527), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n362), .A2(new_n434), .A3(G953), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n522), .A2(new_n532), .A3(new_n534), .ZN(new_n537));
  AOI21_X1  g351(.A(G902), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G478), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n538), .B(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n544));
  OAI21_X1  g358(.A(G131), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n544), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n196), .A3(new_n542), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n542), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT17), .A3(G131), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n549), .A2(new_n339), .A3(new_n340), .A4(new_n551), .ZN(new_n552));
  OAI22_X1  g366(.A1(new_n346), .A2(new_n347), .B1(new_n207), .B2(new_n345), .ZN(new_n553));
  NAND2_X1  g367(.A1(KEYINPUT18), .A2(G131), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n542), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n550), .A2(KEYINPUT18), .A3(G131), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(G113), .B(G122), .Z(new_n558));
  XOR2_X1   g372(.A(KEYINPUT85), .B(G104), .Z(new_n559));
  XOR2_X1   g373(.A(new_n558), .B(new_n559), .Z(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n552), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n561), .B1(new_n552), .B2(new_n557), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n357), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G475), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT20), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT19), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT19), .B1(new_n334), .B2(new_n336), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n207), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n340), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n545), .B2(new_n547), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n560), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n562), .ZN(new_n575));
  NOR2_X1   g389(.A1(G475), .A2(G902), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n567), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n576), .ZN(new_n578));
  AOI211_X1 g392(.A(KEYINPUT20), .B(new_n578), .C1(new_n574), .C2(new_n562), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n566), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(G234), .A2(G237), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(G952), .A3(new_n318), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT21), .B(G898), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(G902), .A3(G953), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n541), .A2(new_n580), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n374), .A2(new_n438), .A3(new_n508), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  OAI21_X1  g404(.A(G472), .B1(new_n292), .B2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n313), .A2(new_n293), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n372), .A2(new_n433), .A3(new_n437), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT89), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT91), .ZN(new_n598));
  INV_X1    g412(.A(new_n537), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n534), .B1(new_n522), .B2(new_n532), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n598), .B(KEYINPUT33), .C1(new_n599), .C2(new_n600), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(G478), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n539), .A2(new_n357), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n538), .B2(new_n539), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n606), .B1(new_n605), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n580), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT90), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n503), .A2(new_n507), .ZN(new_n614));
  INV_X1    g428(.A(new_n440), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI211_X1 g430(.A(KEYINPUT90), .B(new_n440), .C1(new_n503), .C2(new_n507), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n586), .B(new_n612), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n597), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT34), .B(G104), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  XNOR2_X1  g435(.A(new_n508), .B(new_n613), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n538), .B(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n624), .A2(new_n580), .A3(new_n587), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n596), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G107), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NAND2_X1  g443(.A1(new_n355), .A2(new_n342), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n321), .A2(KEYINPUT36), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n366), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n359), .A2(new_n361), .A3(new_n363), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n433), .A2(new_n437), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n593), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n508), .A2(new_n638), .A3(new_n588), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  XOR2_X1   g455(.A(new_n582), .B(KEYINPUT94), .Z(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(G900), .B2(new_n585), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n624), .A2(new_n580), .A3(new_n644), .ZN(new_n645));
  AND4_X1   g459(.A1(new_n316), .A2(new_n438), .A3(new_n636), .A4(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(new_n616), .B2(new_n617), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT95), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n646), .B(KEYINPUT95), .C1(new_n616), .C2(new_n617), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  AND2_X1   g466(.A1(new_n298), .A2(new_n315), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n301), .B1(new_n289), .B2(new_n264), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n264), .A2(new_n301), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n357), .B1(new_n299), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n659), .A2(new_n660), .B1(new_n592), .B2(new_n187), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT98), .Z(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n643), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n438), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT40), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT101), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n614), .B(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n580), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n636), .A2(new_n672), .A3(new_n440), .A4(new_n624), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT99), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  AND4_X1   g489(.A1(new_n663), .A2(new_n668), .A3(new_n669), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n209), .ZN(G45));
  OAI211_X1 g491(.A(new_n580), .B(new_n643), .C1(new_n609), .C2(new_n610), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n616), .B2(new_n617), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT102), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n316), .A2(new_n438), .A3(new_n636), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n684), .B(new_n679), .C1(new_n616), .C2(new_n617), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NAND2_X1  g501(.A1(new_n422), .A2(new_n407), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n405), .A2(new_n229), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n689), .A2(new_n452), .B1(new_n391), .B2(new_n393), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n410), .B1(new_n690), .B2(new_n395), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n395), .B1(new_n390), .B2(new_n415), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT12), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n688), .A2(new_n410), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(G469), .B1(new_n694), .B2(G902), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(KEYINPUT103), .A3(new_n424), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(G469), .C1(new_n694), .C2(G902), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT104), .B1(new_n699), .B2(new_n437), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n701), .B(new_n436), .C1(new_n696), .C2(new_n698), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n374), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n618), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT41), .B(G113), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NOR3_X1   g521(.A1(new_n373), .A2(new_n700), .A3(new_n702), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n622), .A2(new_n625), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  AND3_X1   g524(.A1(new_n316), .A2(new_n588), .A3(new_n636), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n622), .A2(new_n703), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT105), .B(G119), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G21));
  NOR2_X1   g528(.A1(new_n672), .A2(new_n624), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n716), .B1(new_n364), .B2(new_n371), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n635), .A2(KEYINPUT106), .A3(new_n370), .A4(new_n367), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI22_X1  g533(.A1(new_n310), .A2(new_n311), .B1(new_n192), .B2(new_n300), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n293), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n719), .A2(new_n591), .A3(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n700), .A2(new_n702), .A3(new_n587), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n622), .A2(new_n715), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NAND3_X1  g539(.A1(new_n591), .A2(new_n636), .A3(new_n721), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n678), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n703), .B(new_n727), .C1(new_n616), .C2(new_n617), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  NAND3_X1  g543(.A1(new_n503), .A2(new_n615), .A3(new_n507), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n429), .B2(new_n430), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n412), .A2(KEYINPUT77), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(KEYINPUT107), .A3(new_n422), .A4(new_n428), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(G469), .A3(new_n426), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n424), .A2(new_n432), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n437), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n424), .A2(new_n432), .ZN(new_n742));
  INV_X1    g556(.A(new_n426), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n733), .B2(new_n735), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n742), .B1(G469), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT108), .B1(new_n745), .B2(new_n436), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n731), .A2(new_n741), .A3(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n295), .A2(new_n309), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n313), .A2(new_n296), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n679), .A3(new_n719), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT42), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n740), .B1(new_n739), .B2(new_n437), .ZN(new_n753));
  AOI211_X1 g567(.A(KEYINPUT108), .B(new_n436), .C1(new_n737), .C2(new_n738), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n753), .A2(new_n754), .A3(new_n730), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n374), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n196), .ZN(G33));
  NOR2_X1   g573(.A1(new_n753), .A2(new_n730), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(new_n374), .A3(new_n645), .A4(new_n741), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND2_X1  g576(.A1(new_n593), .A2(new_n636), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT109), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n672), .B1(new_n609), .B2(new_n610), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT43), .Z(new_n766));
  AND2_X1   g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n767), .A2(KEYINPUT44), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n744), .A2(KEYINPUT45), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n429), .A2(new_n430), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n743), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n770), .B(G469), .C1(KEYINPUT45), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT46), .B1(new_n773), .B2(new_n432), .ZN(new_n774));
  INV_X1    g588(.A(new_n424), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n432), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n436), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n665), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n768), .A2(new_n769), .A3(new_n779), .A4(new_n730), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n202), .ZN(G39));
  NOR4_X1   g595(.A1(new_n730), .A2(new_n316), .A3(new_n372), .A4(new_n678), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n778), .A2(KEYINPUT47), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NOR2_X1   g602(.A1(new_n636), .A2(new_n644), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n375), .B(new_n743), .C1(new_n733), .C2(new_n735), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n789), .B(new_n437), .C1(new_n790), .C2(new_n742), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n653), .B2(new_n661), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n792), .B(new_n715), .C1(new_n616), .C2(new_n617), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n728), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n686), .A2(new_n794), .A3(new_n651), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT52), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n724), .A2(new_n709), .A3(new_n712), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n541), .A2(new_n580), .A3(new_n644), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n503), .A2(new_n507), .A3(new_n615), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n682), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n755), .B2(new_n727), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n752), .A3(new_n757), .A4(new_n761), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT113), .B1(new_n624), .B2(new_n580), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n577), .A2(new_n579), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n541), .A3(new_n805), .A4(new_n566), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n587), .B1(new_n807), .B2(new_n611), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n508), .A3(new_n595), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(new_n639), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n810), .B(new_n589), .C1(new_n618), .C2(new_n704), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n797), .A2(new_n802), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n686), .A2(new_n794), .A3(new_n651), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n796), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n796), .A2(new_n812), .A3(KEYINPUT53), .A4(new_n814), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n819), .A2(new_n818), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT54), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n817), .A2(new_n823), .A3(new_n819), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n817), .A2(new_n819), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT115), .B1(new_n827), .B2(KEYINPUT54), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n822), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n642), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n766), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(new_n722), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n731), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT116), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n783), .A2(new_n784), .ZN(new_n835));
  INV_X1    g649(.A(new_n699), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n437), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(KEYINPUT116), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n834), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n615), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n671), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n832), .A2(new_n703), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n840), .A2(new_n841), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n703), .A2(new_n731), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n831), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(new_n726), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n844), .A2(new_n845), .ZN(new_n852));
  INV_X1    g666(.A(new_n372), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n663), .A2(new_n847), .A3(new_n853), .A4(new_n582), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n609), .A2(new_n610), .A3(new_n580), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n839), .A2(new_n851), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n832), .A2(new_n622), .A3(new_n703), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(G952), .A3(new_n318), .ZN(new_n862));
  INV_X1    g676(.A(new_n719), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n748), .B2(new_n749), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n831), .A2(new_n848), .A3(new_n864), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT48), .Z(new_n866));
  AOI211_X1 g680(.A(new_n862), .B(new_n866), .C1(new_n612), .C2(new_n854), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n839), .A2(new_n851), .A3(KEYINPUT51), .A4(new_n857), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n860), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n829), .A2(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n863), .A2(new_n765), .A3(new_n436), .A4(new_n440), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT111), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n836), .A2(KEYINPUT49), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(KEYINPUT111), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT112), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n671), .B1(KEYINPUT49), .B2(new_n836), .ZN(new_n878));
  OR3_X1    g692(.A1(new_n877), .A2(new_n663), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n870), .A2(new_n879), .ZN(G75));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n357), .B1(new_n817), .B2(new_n819), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(G210), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n460), .A2(new_n463), .A3(new_n465), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n475), .ZN(new_n887));
  XOR2_X1   g701(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n885), .A2(new_n889), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n318), .A2(G952), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G51));
  XOR2_X1   g707(.A(new_n432), .B(KEYINPUT57), .Z(new_n894));
  AOI21_X1  g708(.A(new_n823), .B1(new_n817), .B2(new_n819), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n824), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n689), .A2(new_n452), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n395), .B1(new_n899), .B2(new_n394), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n410), .B1(new_n425), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n691), .A2(new_n693), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(KEYINPUT119), .B(new_n894), .C1(new_n824), .C2(new_n895), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n773), .B(KEYINPUT120), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n882), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n892), .B1(new_n905), .B2(new_n907), .ZN(G54));
  INV_X1    g722(.A(new_n575), .ZN(new_n909));
  NAND2_X1  g723(.A1(KEYINPUT58), .A2(G475), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n909), .B1(new_n883), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n892), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .A4(new_n575), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n911), .A2(KEYINPUT121), .A3(new_n912), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(G60));
  NAND2_X1  g732(.A1(new_n603), .A2(new_n604), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n607), .B(KEYINPUT59), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n829), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n824), .A2(new_n895), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n919), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n912), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n922), .A2(new_n925), .ZN(G63));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT60), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n827), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n365), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n892), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT61), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n632), .B2(new_n929), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI221_X1 g749(.A(new_n931), .B1(new_n932), .B2(KEYINPUT61), .C1(new_n632), .C2(new_n929), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(G66));
  OAI21_X1  g751(.A(G953), .B1(new_n583), .B2(new_n472), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT123), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n797), .A2(new_n811), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(G953), .ZN(new_n941));
  MUX2_X1   g755(.A(new_n939), .B(KEYINPUT123), .S(new_n941), .Z(new_n942));
  OAI21_X1  g756(.A(new_n886), .B1(G898), .B2(new_n318), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  AOI211_X1 g758(.A(new_n666), .B(new_n730), .C1(new_n611), .C2(new_n807), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n780), .B1(new_n374), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n686), .A2(new_n651), .A3(new_n728), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT62), .B1(new_n676), .B2(new_n947), .ZN(new_n948));
  OR3_X1    g762(.A1(new_n676), .A2(new_n947), .A3(KEYINPUT62), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n946), .A2(new_n787), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n318), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n281), .A2(new_n282), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n569), .A2(new_n570), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n954), .B1(G900), .B2(G953), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n622), .A2(new_n715), .A3(new_n864), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n779), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n780), .A2(new_n947), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n752), .A2(new_n757), .A3(new_n761), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT125), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n787), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n957), .B1(new_n963), .B2(G953), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n955), .A2(new_n956), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n318), .B1(G227), .B2(G900), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n955), .A2(new_n956), .A3(new_n968), .A4(new_n964), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(G72));
  NOR2_X1   g784(.A1(new_n283), .A2(new_n655), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n960), .A2(new_n787), .A3(new_n940), .A4(new_n962), .ZN(new_n972));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  AND3_X1   g788(.A1(new_n972), .A2(KEYINPUT126), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT126), .B1(new_n972), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n283), .A2(new_n284), .ZN(new_n978));
  OAI221_X1 g792(.A(new_n974), .B1(new_n978), .B2(new_n307), .C1(new_n820), .C2(new_n821), .ZN(new_n979));
  INV_X1    g793(.A(new_n940), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n974), .B1(new_n950), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n892), .B1(new_n981), .B2(new_n654), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n977), .A2(new_n979), .A3(new_n982), .ZN(G57));
endmodule


