//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n639,
    new_n640, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  OR2_X1    g034(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(KEYINPUT3), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G2104), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n462), .A2(new_n467), .A3(G137), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n460), .A2(new_n461), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n464), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  INV_X1    g051(.A(G113), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n472), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(G2105), .B2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n462), .A2(new_n467), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n484), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n483), .A2(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n462), .A2(new_n467), .A3(KEYINPUT4), .A4(G138), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n462), .A2(new_n467), .A3(G126), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n484), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n473), .A2(new_n474), .A3(G138), .A4(new_n484), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n493), .A2(new_n496), .A3(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT72), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT72), .A3(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT71), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n511), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(new_n506), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n514), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n510), .B1(new_n519), .B2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND2_X1  g097(.A1(new_n516), .A2(G51), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n513), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XOR2_X1   g100(.A(new_n525), .B(KEYINPUT7), .Z(new_n526));
  INV_X1    g101(.A(new_n506), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n523), .A2(new_n524), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n506), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n516), .A2(G52), .B1(new_n509), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n513), .A2(G90), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(KEYINPUT74), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT74), .B1(new_n535), .B2(new_n536), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(new_n513), .A2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n516), .A2(G43), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n506), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(new_n509), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND3_X1  g129(.A1(new_n516), .A2(KEYINPUT9), .A3(G53), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT9), .B1(new_n516), .B2(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT75), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n557), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n559), .A2(new_n560), .A3(new_n555), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT76), .B(G65), .Z(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n563), .B2(new_n506), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n513), .A2(G91), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n558), .A2(new_n561), .A3(new_n565), .ZN(G299));
  NAND2_X1  g141(.A1(G49), .A2(G543), .ZN(new_n567));
  OR3_X1    g142(.A1(new_n512), .A2(KEYINPUT77), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT77), .B1(new_n512), .B2(new_n567), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n506), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n513), .A2(G87), .B1(G651), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G48), .A2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n512), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n513), .A2(new_n577), .A3(G86), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n579));
  OR2_X1    g154(.A1(KEYINPUT71), .A2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(KEYINPUT71), .A2(G651), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n527), .B(G86), .C1(new_n582), .C2(new_n511), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT80), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n576), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n503), .A2(new_n505), .A3(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(new_n509), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(KEYINPUT78), .A3(new_n509), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n586), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT78), .B1(new_n589), .B2(new_n509), .ZN(new_n595));
  AND2_X1   g170(.A1(KEYINPUT71), .A2(G651), .ZN(new_n596));
  NOR2_X1   g171(.A1(KEYINPUT71), .A2(G651), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI211_X1 g173(.A(new_n591), .B(new_n598), .C1(new_n587), .C2(new_n588), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n595), .A2(new_n599), .A3(KEYINPUT79), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n585), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(new_n516), .A2(G47), .ZN(new_n605));
  INV_X1    g180(.A(new_n512), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n527), .ZN(new_n607));
  INV_X1    g182(.A(G85), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT83), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G72), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G60), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n506), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n509), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT82), .Z(new_n616));
  OAI211_X1 g191(.A(new_n605), .B(KEYINPUT83), .C1(new_n608), .C2(new_n607), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n611), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(KEYINPUT84), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n611), .A2(new_n616), .A3(new_n620), .A4(new_n617), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(G290));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n607), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n513), .A2(KEYINPUT10), .A3(G92), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(G79), .A2(G543), .ZN(new_n628));
  INV_X1    g203(.A(G66), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n506), .B2(new_n629), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n516), .A2(G54), .B1(G651), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  MUX2_X1   g207(.A(new_n632), .B(G301), .S(G868), .Z(G284));
  XOR2_X1   g208(.A(G284), .B(KEYINPUT85), .Z(G321));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(G299), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(G168), .ZN(G297));
  OAI21_X1  g212(.A(new_n636), .B1(new_n635), .B2(G168), .ZN(G280));
  AND2_X1   g213(.A1(new_n627), .A2(new_n631), .ZN(new_n639));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G860), .ZN(G148));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G868), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n485), .A2(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(G99), .A2(G2105), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(new_n484), .B2(G111), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n481), .A2(KEYINPUT88), .A3(G135), .ZN(new_n649));
  AOI21_X1  g224(.A(KEYINPUT88), .B1(new_n481), .B2(G135), .ZN(new_n650));
  OAI221_X1 g225(.A(new_n646), .B1(new_n647), .B2(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT3), .B(G2104), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n469), .A2(new_n653), .A3(new_n484), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n654), .B(new_n655), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT87), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n652), .A2(new_n659), .ZN(G156));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(KEYINPUT14), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1341), .B(G1348), .Z(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2443), .B(G2446), .Z(new_n672));
  XNOR2_X1  g247(.A(G2451), .B(G2454), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(G14), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n675), .B2(new_n671), .ZN(G401));
  XNOR2_X1  g252(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(KEYINPUT17), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2072), .B(G2078), .Z(new_n685));
  AOI21_X1  g260(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n684), .B2(new_n685), .ZN(new_n688));
  XOR2_X1   g263(.A(G2096), .B(G2100), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT91), .ZN(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT20), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n695), .A2(new_n696), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n701), .C1(new_n692), .C2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT92), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1991), .B(G1996), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1981), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n706), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(G229));
  INV_X1    g287(.A(KEYINPUT100), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n481), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n485), .A2(G119), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n484), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n715), .B1(new_n724), .B2(G29), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT94), .B(G16), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(G290), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G24), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n729), .ZN(new_n732));
  INV_X1    g307(.A(G1986), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n730), .B(G1986), .C1(new_n731), .C2(new_n729), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n727), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n570), .B2(new_n573), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(G23), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT33), .B(G1976), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT95), .ZN(new_n741));
  OR3_X1    g316(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n738), .B2(new_n739), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n510), .B(new_n729), .C1(new_n519), .C2(new_n520), .ZN(new_n745));
  INV_X1    g320(.A(G1971), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n729), .A2(G22), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n746), .B1(new_n745), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n602), .A2(G16), .A3(new_n603), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G6), .B2(G16), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT32), .B(G1981), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n750), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n751), .B(new_n753), .C1(G6), .C2(G16), .ZN(new_n756));
  AND3_X1   g331(.A1(new_n755), .A2(KEYINPUT34), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(KEYINPUT34), .B1(new_n755), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n736), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT36), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT36), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n736), .B(new_n761), .C1(new_n757), .C2(new_n758), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n737), .A2(G4), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n639), .B2(new_n737), .ZN(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n714), .A2(G27), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT99), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n494), .A2(new_n495), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n499), .B1(new_n770), .B2(G2105), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n491), .A2(new_n492), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(new_n484), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n769), .B1(new_n774), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2078), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n737), .A2(G5), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G301), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n767), .B(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n481), .A2(G141), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n485), .A2(G129), .ZN(new_n782));
  NAND3_X1  g357(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT26), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n484), .A2(G105), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n785), .A2(new_n786), .B1(new_n469), .B2(new_n787), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n781), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G29), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G29), .B2(G32), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT24), .ZN(new_n796));
  INV_X1    g371(.A(G34), .ZN(new_n797));
  AOI21_X1  g372(.A(G29), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G160), .B2(new_n714), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G2084), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n481), .A2(G139), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT25), .Z(new_n804));
  AOI22_X1  g379(.A1(new_n653), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n802), .B(new_n804), .C1(new_n484), .C2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G33), .B(new_n806), .S(G29), .Z(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G2072), .Z(new_n808));
  AND3_X1   g383(.A1(new_n795), .A2(new_n801), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n780), .B1(new_n809), .B2(KEYINPUT97), .ZN(new_n810));
  INV_X1    g385(.A(new_n794), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n792), .B(new_n811), .C1(G29), .C2(G32), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n800), .A2(G2084), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n778), .A2(new_n779), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT98), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n728), .A2(G20), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT23), .Z(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G299), .B2(G16), .ZN(new_n819));
  INV_X1    g394(.A(G1956), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n795), .A2(new_n801), .A3(new_n808), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n714), .A2(G35), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G162), .B2(new_n714), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT29), .ZN(new_n827));
  INV_X1    g402(.A(G2090), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(KEYINPUT29), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n729), .A2(G19), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n549), .B2(new_n729), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(G1341), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n737), .A2(G21), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G168), .B2(new_n737), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(G1966), .ZN(new_n837));
  INV_X1    g412(.A(G28), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT30), .ZN(new_n839));
  AOI21_X1  g414(.A(G29), .B1(new_n838), .B2(KEYINPUT30), .ZN(new_n840));
  OR2_X1    g415(.A1(KEYINPUT31), .A2(G11), .ZN(new_n841));
  NAND2_X1  g416(.A1(KEYINPUT31), .A2(G11), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n839), .A2(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n651), .B2(new_n714), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n836), .B2(G1966), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n481), .A2(G140), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n485), .A2(G128), .ZN(new_n847));
  OR2_X1    g422(.A1(G104), .A2(G2105), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(G2104), .C1(G116), .C2(new_n484), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(G29), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n714), .A2(G26), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT28), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G2067), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n834), .A2(new_n837), .A3(new_n845), .A4(new_n856), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n830), .A2(new_n831), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n810), .A2(new_n816), .A3(new_n824), .A4(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n713), .B1(new_n763), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g436(.A(KEYINPUT100), .B(new_n859), .C1(new_n760), .C2(new_n762), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(G311));
  NAND2_X1  g438(.A1(new_n763), .A2(new_n860), .ZN(G150));
  NAND2_X1  g439(.A1(new_n639), .A2(G559), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(new_n598), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n516), .A2(G55), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n513), .A2(G93), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT102), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT102), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n548), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n549), .B(new_n869), .C1(new_n872), .C2(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n867), .B(new_n877), .Z(new_n878));
  AND2_X1   g453(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n879), .A2(new_n880), .A3(G860), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n874), .A2(G860), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT37), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n881), .A2(new_n883), .ZN(G145));
  XNOR2_X1  g459(.A(new_n774), .B(new_n850), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n806), .ZN(new_n886));
  INV_X1    g461(.A(new_n656), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n722), .A2(new_n723), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n485), .A2(G130), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n481), .A2(G142), .ZN(new_n892));
  NOR2_X1   g467(.A1(G106), .A2(G2105), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(new_n484), .B2(G118), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n891), .A2(new_n895), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n724), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n789), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n888), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n888), .A2(new_n901), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n651), .B(G160), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(G162), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g487(.A1(new_n874), .A2(new_n635), .ZN(new_n913));
  INV_X1    g488(.A(G288), .ZN(new_n914));
  NAND2_X1  g489(.A1(G290), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n619), .A2(G288), .A3(new_n621), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n603), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n601), .A2(KEYINPUT81), .ZN(new_n919));
  OAI21_X1  g494(.A(G166), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n602), .A2(G303), .A3(new_n603), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n915), .A2(new_n920), .A3(new_n916), .A4(new_n921), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n877), .B(new_n642), .ZN(new_n928));
  INV_X1    g503(.A(new_n565), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n559), .A2(new_n555), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n930), .B2(KEYINPUT75), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n561), .A3(new_n632), .ZN(new_n932));
  AND3_X1   g507(.A1(G299), .A2(KEYINPUT104), .A3(new_n639), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT104), .B1(G299), .B2(new_n639), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G299), .A2(new_n639), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT41), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n632), .B1(new_n931), .B2(new_n561), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT104), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(G299), .A2(new_n639), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT41), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n938), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n936), .B1(new_n947), .B2(new_n928), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n926), .A2(new_n927), .B1(KEYINPUT105), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(KEYINPUT105), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n926), .A2(new_n927), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n913), .B1(new_n952), .B2(new_n635), .ZN(G295));
  OAI21_X1  g528(.A(new_n913), .B1(new_n952), .B2(new_n635), .ZN(G331));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n944), .B1(new_n940), .B2(new_n942), .ZN(new_n956));
  OAI21_X1  g531(.A(G168), .B1(new_n538), .B2(new_n539), .ZN(new_n957));
  INV_X1    g532(.A(new_n539), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(G286), .A3(new_n537), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n877), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n875), .A2(new_n957), .A3(new_n959), .A4(new_n876), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(new_n965), .A3(new_n962), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n877), .A2(new_n960), .A3(KEYINPUT106), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n943), .A2(new_n946), .ZN(new_n969));
  INV_X1    g544(.A(new_n938), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n964), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G37), .B1(new_n972), .B2(new_n925), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n935), .A2(new_n945), .B1(new_n937), .B2(new_n946), .ZN(new_n974));
  INV_X1    g549(.A(new_n963), .ZN(new_n975));
  OAI22_X1  g550(.A1(new_n968), .A2(new_n956), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n925), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n924), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n973), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n966), .A2(new_n967), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n947), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n978), .B(new_n979), .C1(new_n984), .C2(new_n964), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n981), .B1(new_n973), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n955), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n973), .A2(new_n985), .A3(new_n981), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n981), .B1(new_n973), .B2(new_n980), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT44), .B(new_n988), .C1(new_n989), .C2(KEYINPUT108), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n991), .B(new_n981), .C1(new_n973), .C2(new_n980), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(new_n990), .B2(new_n992), .ZN(G397));
  AOI21_X1  g568(.A(G1384), .B1(new_n771), .B2(new_n773), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(KEYINPUT45), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n996));
  INV_X1    g571(.A(G40), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n478), .B2(G2105), .ZN(new_n998));
  AND2_X1   g573(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n999));
  NOR2_X1   g574(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G101), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(G2104), .B1(KEYINPUT69), .B2(KEYINPUT3), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1001), .A2(KEYINPUT3), .B1(new_n1005), .B2(new_n466), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1006), .B2(G137), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n996), .B(new_n998), .C1(new_n1007), .C2(G2105), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n477), .A2(new_n472), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n653), .B2(G125), .ZN(new_n1010));
  OAI21_X1  g585(.A(G40), .B1(new_n1010), .B2(new_n484), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT109), .B1(new_n471), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n995), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n850), .B(new_n855), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT110), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n889), .A2(new_n726), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n789), .B(G1996), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n889), .A2(new_n726), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G290), .A2(G1986), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n619), .A2(new_n733), .A3(new_n621), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1015), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G1384), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n774), .A2(new_n1028), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(G164), .B2(G1384), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT56), .B(G2072), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI211_X1 g607(.A(KEYINPUT50), .B(G1384), .C1(new_n771), .C2(new_n773), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1013), .B1(new_n994), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n1035), .B2(KEYINPUT117), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1013), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1032), .B1(new_n1040), .B2(new_n820), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n558), .A2(new_n561), .A3(KEYINPUT57), .A4(new_n565), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1043), .B1(new_n930), .B2(new_n929), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1026), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1956), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1045), .ZN(new_n1048));
  NOR4_X1   g623(.A1(new_n1047), .A2(new_n1048), .A3(KEYINPUT119), .A4(new_n1032), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1047), .B2(new_n1032), .ZN(new_n1051));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n774), .A2(new_n1034), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1037), .A2(new_n1013), .A3(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1013), .A2(new_n994), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1054), .A2(new_n766), .B1(new_n1055), .B2(new_n855), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1056), .A2(new_n632), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1050), .A2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n1051), .A2(KEYINPUT121), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(new_n1048), .C1(new_n1047), .C2(new_n1032), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1060), .B1(new_n1050), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1056), .A2(KEYINPUT60), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n1056), .B2(KEYINPUT60), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1068), .B2(new_n632), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n766), .B1(new_n1035), .B2(new_n1033), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1055), .A2(new_n855), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(KEYINPUT60), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT122), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1056), .A2(new_n1067), .A3(KEYINPUT60), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n639), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1040), .A2(new_n820), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1032), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1045), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(new_n1051), .A3(KEYINPUT61), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT58), .B(G1341), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1081), .A2(G1996), .B1(new_n1055), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n549), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1084), .B(KEYINPUT59), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1076), .A2(new_n1080), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1059), .B1(new_n1065), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1081), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(G2078), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1089), .A2(new_n1091), .B1(new_n1054), .B2(new_n779), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n774), .A2(new_n1028), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1013), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT111), .B1(new_n1094), .B2(new_n995), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT111), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1029), .A2(new_n1096), .A3(new_n1030), .ZN(new_n1097));
  AOI21_X1  g672(.A(G2078), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1092), .B(G301), .C1(new_n1098), .C2(KEYINPUT53), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT126), .ZN(new_n1100));
  INV_X1    g675(.A(G2078), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1097), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1096), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1090), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(G301), .A4(new_n1092), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1088), .B1(new_n1100), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT125), .B(G2078), .ZN(new_n1109));
  NOR4_X1   g684(.A1(new_n471), .A2(new_n1011), .A3(new_n1090), .A4(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1030), .A2(new_n1093), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1098), .B2(KEYINPUT53), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1054), .A2(new_n1113), .A3(new_n779), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1054), .B2(new_n779), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT127), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1116), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1114), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1105), .A2(new_n1120), .A3(new_n1121), .A4(new_n1111), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(G171), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1108), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1013), .A2(new_n994), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n570), .A2(G1976), .A3(new_n573), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(G8), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1128), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1125), .A2(G8), .A3(new_n1126), .A4(new_n1130), .ZN(new_n1131));
  OR3_X1    g706(.A1(new_n914), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(G8), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1055), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT115), .B(G1981), .Z(new_n1136));
  OAI211_X1 g711(.A(new_n585), .B(new_n1136), .C1(new_n594), .C2(new_n600), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n592), .A2(new_n593), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n583), .B1(new_n512), .B2(new_n575), .ZN(new_n1139));
  OAI21_X1  g714(.A(G1981), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(KEYINPUT49), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT49), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1135), .B(new_n1141), .C1(new_n1142), .C2(KEYINPUT116), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1142), .A2(KEYINPUT116), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1133), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(G303), .A2(G8), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1095), .A2(new_n746), .A3(new_n1097), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1035), .A2(KEYINPUT117), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(new_n1039), .A3(new_n828), .A4(new_n1053), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(G8), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1145), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(G1966), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1081), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G2084), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1037), .A2(new_n1053), .A3(new_n1158), .A4(new_n1013), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1134), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(G286), .A2(G8), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT51), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1035), .A2(G2084), .A3(new_n1033), .ZN(new_n1165));
  AOI21_X1  g740(.A(G1966), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1166));
  OAI211_X1 g741(.A(G8), .B(G168), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1161), .B(KEYINPUT123), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1167), .B1(new_n1160), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1164), .B1(new_n1170), .B2(KEYINPUT51), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1150), .A2(KEYINPUT112), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT112), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1095), .A2(new_n1173), .A3(new_n746), .A4(new_n1097), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1054), .A2(G2090), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(G8), .B(new_n1148), .C1(new_n1172), .C2(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1155), .A2(new_n1171), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1092), .B1(new_n1098), .B2(KEYINPUT53), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(G171), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1105), .A2(new_n1120), .A3(new_n1111), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(G171), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1088), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1124), .A2(new_n1178), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1087), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1167), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1154), .A2(new_n1149), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1145), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1177), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(G8), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1149), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1145), .A2(new_n1190), .A3(new_n1167), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1193), .A2(new_n1177), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1177), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1180), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n1199));
  OAI21_X1  g774(.A(G8), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n1168), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1162), .B1(new_n1201), .B2(new_n1167), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1199), .B1(new_n1202), .B2(new_n1164), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1171), .A2(KEYINPUT62), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1197), .A2(new_n1198), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1177), .A2(new_n1145), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1207), .A2(G1976), .A3(G288), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1137), .ZN(new_n1209));
  OR2_X1    g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1206), .B1(new_n1210), .B2(new_n1135), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1196), .A2(new_n1205), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1025), .B1(new_n1185), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1214));
  OAI22_X1  g789(.A1(new_n1214), .A2(new_n1020), .B1(G2067), .B2(new_n850), .ZN(new_n1215));
  AND2_X1   g790(.A1(new_n1215), .A2(new_n1015), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1023), .A2(new_n1014), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n1217), .B(KEYINPUT48), .Z(new_n1218));
  NAND2_X1  g793(.A1(new_n1021), .A2(new_n1015), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT47), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT46), .ZN(new_n1222));
  OR3_X1    g797(.A1(new_n1014), .A2(new_n1222), .A3(G1996), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1222), .B1(new_n1014), .B2(G1996), .ZN(new_n1224));
  AND2_X1   g799(.A1(new_n1017), .A2(new_n789), .ZN(new_n1225));
  OAI211_X1 g800(.A(new_n1223), .B(new_n1224), .C1(new_n1225), .C2(new_n1014), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1220), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  AOI211_X1 g802(.A(new_n1216), .B(new_n1227), .C1(new_n1221), .C2(new_n1226), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1213), .A2(new_n1228), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g804(.A(G319), .ZN(new_n1231));
  OR3_X1    g805(.A1(G401), .A2(new_n1231), .A3(G227), .ZN(new_n1232));
  NOR2_X1   g806(.A1(G229), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g807(.A(new_n911), .B(new_n1233), .C1(new_n982), .C2(new_n986), .ZN(G225));
  INV_X1    g808(.A(G225), .ZN(G308));
endmodule


