//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  AOI21_X1  g000(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n202));
  OR2_X1    g001(.A1(G197gat), .A2(G204gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT29), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT3), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G141gat), .B(G148gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  OAI22_X1  g020(.A1(new_n219), .A2(KEYINPUT77), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n220), .B(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n213), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n211), .B1(new_n226), .B2(new_n212), .ZN(new_n227));
  INV_X1    g026(.A(G228gat), .ZN(new_n228));
  INV_X1    g027(.A(G233gat), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n224), .A2(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n227), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n228), .A2(new_n229), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n231), .B(new_n232), .C1(new_n223), .C2(new_n213), .ZN(new_n233));
  INV_X1    g032(.A(G22gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n234), .B1(new_n230), .B2(new_n233), .ZN(new_n237));
  XNOR2_X1  g036(.A(G78gat), .B(G106gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G50gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n236), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n237), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n230), .A2(new_n233), .A3(KEYINPUT81), .A4(new_n234), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n241), .B(KEYINPUT80), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT82), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(KEYINPUT82), .A3(new_n248), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n242), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G8gat), .B(G36gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(G64gat), .B(G92gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT76), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n258));
  INV_X1    g057(.A(G183gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G190gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT67), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n260), .A2(new_n262), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270));
  NAND3_X1  g069(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n266), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT68), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n266), .A2(new_n272), .A3(new_n276), .A4(new_n273), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(G169gat), .B2(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n278), .A2(G169gat), .A3(G176gat), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n275), .A2(new_n277), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT64), .B1(new_n281), .B2(new_n283), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n288), .A2(new_n289), .A3(new_n279), .A4(new_n280), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n270), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n291), .B(new_n273), .C1(G183gat), .C2(G190gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n286), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n282), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n287), .A2(KEYINPUT26), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n267), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(new_n287), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT27), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(KEYINPUT27), .B2(G183gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n262), .A2(new_n264), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT28), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT28), .ZN(new_n308));
  AND2_X1   g107(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n301), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n257), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n285), .A2(new_n319), .A3(new_n294), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n319), .B1(new_n285), .B2(new_n294), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT27), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(new_n260), .B2(new_n265), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n306), .B1(new_n324), .B2(new_n310), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n312), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n301), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT70), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n330), .B(new_n301), .C1(new_n307), .C2(new_n312), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT29), .B1(new_n322), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n318), .B1(new_n333), .B2(new_n316), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n285), .A2(new_n294), .A3(new_n319), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n212), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(KEYINPUT76), .A3(new_n315), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n211), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n211), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n335), .A2(new_n332), .A3(new_n336), .A4(new_n316), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n314), .A2(new_n212), .A3(new_n315), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n256), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n317), .B1(new_n338), .B2(new_n315), .ZN(new_n346));
  AOI211_X1 g145(.A(new_n257), .B(new_n316), .C1(new_n337), .C2(new_n212), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n341), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n344), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n255), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(KEYINPUT30), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n316), .B1(new_n337), .B2(new_n212), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n339), .B1(new_n352), .B2(new_n317), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n344), .B1(new_n353), .B2(new_n341), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT30), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n255), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n351), .A2(KEYINPUT83), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT83), .B1(new_n351), .B2(new_n356), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n252), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(G227gat), .A2(G233gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G127gat), .B(G134gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT71), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT1), .ZN(new_n364));
  INV_X1    g163(.A(G113gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G120gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n365), .A2(G120gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(KEYINPUT72), .B2(new_n366), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(KEYINPUT72), .B2(new_n366), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n361), .A2(new_n364), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n363), .A2(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n337), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n373), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n335), .A2(new_n332), .A3(new_n375), .A4(new_n336), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n360), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT74), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT34), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n374), .A2(new_n360), .A3(new_n376), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT32), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT33), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(G15gat), .B(G43gat), .Z(new_n387));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n389), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n383), .B(KEYINPUT32), .C1(new_n385), .C2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n382), .B1(new_n390), .B2(new_n392), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n223), .A2(new_n373), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n223), .A2(new_n373), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n223), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT3), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n226), .A3(new_n375), .ZN(new_n404));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n223), .B(new_n373), .ZN(new_n407));
  INV_X1    g206(.A(new_n405), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(KEYINPUT5), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n398), .A2(new_n411), .A3(new_n400), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n400), .A2(new_n411), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n408), .A2(KEYINPUT5), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n404), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(G57gat), .B(G85gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n410), .A2(new_n415), .A3(new_n420), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n421), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n396), .A2(KEYINPUT35), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n382), .A2(KEYINPUT73), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n394), .B2(new_n395), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n390), .A2(new_n392), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(KEYINPUT73), .A3(new_n382), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n427), .B1(new_n356), .B2(new_n351), .ZN(new_n434));
  INV_X1    g233(.A(new_n242), .ZN(new_n435));
  INV_X1    g234(.A(new_n251), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(new_n249), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n359), .A2(new_n428), .B1(new_n438), .B2(KEYINPUT35), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n434), .A2(new_n437), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n351), .A2(new_n356), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT83), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n351), .A2(KEYINPUT83), .A3(new_n356), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n412), .A2(new_n404), .A3(new_n413), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n408), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n446), .A2(new_n408), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT39), .B1(new_n407), .B2(new_n408), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n420), .B(new_n448), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT40), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n422), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n452), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n451), .A2(KEYINPUT84), .A3(new_n452), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n252), .B1(new_n445), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT87), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT38), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n348), .A2(new_n349), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(new_n256), .C1(new_n462), .C2(KEYINPUT37), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n342), .A2(new_n341), .A3(new_n343), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT85), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n342), .A2(new_n343), .A3(new_n467), .A4(new_n341), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n339), .B(new_n211), .C1(new_n352), .C2(new_n317), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n464), .B1(new_n471), .B2(KEYINPUT37), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  AOI211_X1 g272(.A(KEYINPUT86), .B(new_n473), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n463), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n425), .A2(new_n350), .A3(new_n426), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n460), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n466), .A2(new_n468), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n346), .A2(new_n347), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n211), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT86), .B1(new_n481), .B2(new_n473), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n255), .B1(new_n354), .B2(new_n473), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n471), .A2(new_n464), .A3(KEYINPUT37), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n461), .A4(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(KEYINPUT87), .A3(new_n476), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n462), .A2(KEYINPUT37), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n461), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n478), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n440), .B1(new_n459), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n382), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n431), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n493), .A2(new_n393), .B1(KEYINPUT73), .B2(new_n382), .ZN(new_n494));
  INV_X1    g293(.A(new_n432), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT36), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT36), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n439), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(G29gat), .A2(G36gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT14), .ZN(new_n502));
  AND2_X1   g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(G43gat), .B(G50gat), .Z(new_n505));
  INV_X1    g304(.A(KEYINPUT15), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT89), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n503), .A2(KEYINPUT90), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n503), .A2(KEYINPUT90), .ZN(new_n512));
  NOR4_X1   g311(.A1(new_n507), .A2(new_n502), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n514), .B1(new_n510), .B2(new_n513), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n508), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n508), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n510), .A2(new_n513), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n521), .B1(new_n523), .B2(new_n515), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT17), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G1gat), .B2(new_n526), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n524), .A2(new_n531), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n532), .A2(KEYINPUT18), .A3(new_n533), .A4(new_n535), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n533), .B(KEYINPUT13), .Z(new_n544));
  AND2_X1   g343(.A1(new_n524), .A2(new_n531), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(new_n534), .ZN(new_n546));
  XOR2_X1   g345(.A(G113gat), .B(G141gat), .Z(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G169gat), .B(G197gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT12), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n543), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n546), .A3(new_n543), .ZN(new_n555));
  INV_X1    g354(.A(new_n552), .ZN(new_n556));
  AOI22_X1  g355(.A1(new_n542), .A2(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G134gat), .B(G162gat), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT41), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT97), .ZN(new_n563));
  INV_X1    g362(.A(G99gat), .ZN(new_n564));
  INV_X1    g363(.A(G106gat), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT8), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT98), .ZN(new_n568));
  OAI221_X1 g367(.A(new_n566), .B1(G85gat), .B2(G92gat), .C1(new_n568), .C2(KEYINPUT7), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT7), .B1(new_n567), .B2(KEYINPUT98), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n570), .B1(KEYINPUT98), .B2(new_n567), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(new_n574), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n518), .A2(new_n575), .B1(KEYINPUT41), .B2(new_n560), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n572), .B(new_n573), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n524), .B2(KEYINPUT17), .ZN(new_n578));
  AOI211_X1 g377(.A(new_n519), .B(new_n521), .C1(new_n523), .C2(new_n515), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n578), .A2(KEYINPUT99), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n575), .B1(new_n518), .B2(new_n519), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(new_n525), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n576), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G190gat), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT99), .B1(new_n578), .B2(new_n579), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n581), .A3(new_n525), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n261), .A3(new_n576), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G218gat), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n563), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n585), .A2(G218gat), .A3(new_n589), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n562), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n261), .B1(new_n588), .B2(new_n576), .ZN(new_n595));
  INV_X1    g394(.A(new_n576), .ZN(new_n596));
  AOI211_X1 g395(.A(G190gat), .B(new_n596), .C1(new_n586), .C2(new_n587), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n591), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  AND4_X1   g397(.A1(KEYINPUT97), .A2(new_n598), .A3(new_n593), .A4(new_n562), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n559), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G71gat), .B(G78gat), .Z(new_n604));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G71gat), .B(G78gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT95), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G64gat), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n610), .A2(G57gat), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT94), .B(G57gat), .Z(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(G64gat), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n610), .A2(G57gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n603), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n604), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G127gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n531), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n622), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT96), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G155gat), .ZN(new_n628));
  XOR2_X1   g427(.A(G183gat), .B(G211gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n592), .A2(new_n562), .A3(new_n593), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n598), .A2(new_n593), .A3(KEYINPUT97), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n561), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n636), .A3(new_n558), .ZN(new_n637));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n572), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n618), .A2(new_n577), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n614), .A2(new_n640), .A3(new_n617), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n575), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT10), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n618), .A2(new_n575), .A3(KEYINPUT10), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n638), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n643), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n638), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G120gat), .B(G148gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n600), .A2(new_n633), .A3(new_n637), .A4(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n500), .A2(new_n557), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n427), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT101), .B(G1gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1324gat));
  INV_X1    g460(.A(new_n445), .ZN(new_n662));
  NOR4_X1   g461(.A1(new_n500), .A2(new_n662), .A3(new_n557), .A4(new_n657), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n530), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT102), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT42), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(new_n658), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT36), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n430), .B2(new_n432), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT103), .B1(new_n672), .B2(new_n497), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n496), .A2(new_n674), .A3(new_n498), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n396), .A2(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n670), .B2(new_n678), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n658), .A2(new_n252), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  INV_X1    g481(.A(new_n637), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n558), .B1(new_n634), .B2(new_n636), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(new_n633), .A3(new_n655), .ZN(new_n686));
  INV_X1    g485(.A(new_n440), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n485), .A2(KEYINPUT87), .A3(new_n476), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT87), .B1(new_n485), .B2(new_n476), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n688), .A2(new_n689), .A3(new_n488), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n458), .B1(new_n357), .B2(new_n358), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n437), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n499), .B(new_n687), .C1(new_n690), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n359), .A2(new_n428), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n438), .A2(KEYINPUT35), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n557), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n686), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n427), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n699), .A2(G29gat), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n500), .B2(new_n685), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n687), .B1(new_n690), .B2(new_n692), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n673), .A2(new_n675), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n696), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n685), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n633), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n655), .B(KEYINPUT105), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n698), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(KEYINPUT106), .Z(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n700), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n703), .A2(new_n717), .ZN(G1328gat));
  NOR3_X1   g517(.A1(new_n699), .A2(G36gat), .A3(new_n662), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT46), .ZN(new_n720));
  OAI21_X1  g519(.A(G36gat), .B1(new_n716), .B2(new_n662), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1329gat));
  NOR2_X1   g521(.A1(new_n396), .A2(G43gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI22_X1  g523(.A1(new_n699), .A2(new_n724), .B1(KEYINPUT108), .B2(KEYINPUT47), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n711), .A2(new_n706), .A3(new_n715), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(G43gat), .ZN(new_n727));
  AND2_X1   g526(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1330gat));
  NAND2_X1  g528(.A1(new_n252), .A2(G50gat), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n699), .A2(new_n437), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n716), .A2(new_n730), .B1(new_n731), .B2(G50gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g532(.A(new_n439), .B1(new_n491), .B2(new_n676), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n685), .A2(new_n633), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n734), .A2(new_n735), .A3(new_n698), .A4(new_n713), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n427), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(new_n612), .Z(G1332gat));
  AOI21_X1  g537(.A(new_n662), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT109), .Z(new_n740));
  NAND2_X1  g539(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT110), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1333gat));
  NAND2_X1  g543(.A1(new_n736), .A2(new_n706), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n396), .A2(G71gat), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n745), .A2(G71gat), .B1(new_n736), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n736), .A2(new_n252), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n633), .A2(new_n698), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n655), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT111), .ZN(new_n753));
  INV_X1    g552(.A(new_n709), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n734), .A2(new_n685), .A3(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n697), .B2(new_n708), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n753), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n711), .A2(KEYINPUT112), .A3(new_n753), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762), .B2(new_n700), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n707), .A2(new_n708), .A3(new_n751), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n491), .A2(new_n676), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n685), .B1(new_n767), .B2(new_n696), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(KEYINPUT51), .A3(new_n751), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n700), .A2(new_n656), .A3(G85gat), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT113), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n763), .B1(new_n771), .B2(new_n773), .ZN(G1336gat));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n764), .A2(new_n775), .A3(KEYINPUT51), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT51), .B1(new_n764), .B2(new_n775), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n662), .A2(G92gat), .A3(new_n713), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n760), .A2(new_n445), .A3(new_n761), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(G92gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT51), .B1(new_n768), .B2(new_n751), .ZN(new_n784));
  INV_X1    g583(.A(new_n751), .ZN(new_n785));
  NOR4_X1   g584(.A1(new_n734), .A2(new_n765), .A3(new_n685), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n778), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n783), .ZN(new_n788));
  INV_X1    g587(.A(G92gat), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n752), .B(KEYINPUT111), .Z(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n704), .B2(new_n710), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n789), .B1(new_n791), .B2(new_n445), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n788), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(new_n770), .B2(new_n778), .ZN(new_n795));
  OAI21_X1  g594(.A(G92gat), .B1(new_n758), .B2(new_n662), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT115), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n782), .A2(new_n783), .B1(new_n794), .B2(new_n797), .ZN(G1337gat));
  OAI21_X1  g597(.A(G99gat), .B1(new_n762), .B2(new_n676), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n396), .A2(new_n656), .A3(G99gat), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT116), .Z(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n771), .B2(new_n801), .ZN(G1338gat));
  NOR3_X1   g601(.A1(new_n713), .A2(G106gat), .A3(new_n437), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n776), .A2(new_n777), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n760), .A2(new_n252), .A3(new_n761), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n805), .B1(new_n806), .B2(G106gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n784), .B2(new_n786), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n808), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n565), .B1(new_n791), .B2(new_n252), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT53), .B1(new_n770), .B2(new_n803), .ZN(new_n814));
  OAI21_X1  g613(.A(G106gat), .B1(new_n758), .B2(new_n437), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT117), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n807), .A2(new_n808), .B1(new_n813), .B2(new_n816), .ZN(G1339gat));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n644), .A2(new_n638), .A3(new_n645), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n646), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n652), .B1(new_n646), .B2(KEYINPUT54), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n818), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n821), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n646), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n653), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n533), .B1(new_n532), .B2(new_n535), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n545), .A2(new_n534), .A3(new_n544), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n551), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(KEYINPUT118), .B(new_n551), .C1(new_n828), .C2(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n541), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n553), .A3(new_n539), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n827), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n683), .B2(new_n684), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n834), .A2(new_n836), .A3(new_n655), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n557), .B2(new_n826), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n841), .B(KEYINPUT119), .C1(new_n557), .C2(new_n826), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n600), .A2(new_n844), .A3(new_n637), .A4(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n633), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n657), .A2(new_n698), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n359), .A2(new_n433), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n427), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT121), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n365), .A3(new_n698), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n437), .B1(new_n847), .B2(new_n848), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n396), .B1(new_n854), .B2(KEYINPUT120), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n856), .B(new_n437), .C1(new_n847), .C2(new_n848), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n445), .A2(new_n700), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n858), .A2(new_n557), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n853), .B1(new_n365), .B2(new_n861), .ZN(G1340gat));
  INV_X1    g661(.A(G120gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n852), .A2(new_n863), .A3(new_n655), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n858), .A2(new_n713), .A3(new_n860), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(G1341gat));
  NAND4_X1  g665(.A1(new_n855), .A2(new_n633), .A3(new_n859), .A4(new_n857), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G127gat), .ZN(new_n868));
  OR3_X1    g667(.A1(new_n851), .A2(G127gat), .A3(new_n712), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT122), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n868), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1342gat));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT123), .ZN(new_n876));
  INV_X1    g675(.A(G134gat), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n708), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n876), .B1(new_n851), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n875), .A2(KEYINPUT123), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n858), .A2(new_n685), .A3(new_n860), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n877), .B2(new_n882), .ZN(G1343gat));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n706), .A2(new_n437), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n427), .B(new_n885), .C1(new_n847), .C2(new_n848), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n557), .A2(G141gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n888), .A2(new_n662), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n252), .B1(new_n847), .B2(new_n848), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n600), .A2(new_n637), .A3(new_n842), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n838), .B1(new_n600), .B2(new_n637), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n712), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n698), .B2(new_n657), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n252), .A2(KEYINPUT57), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n892), .A2(new_n893), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n706), .A2(new_n860), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n900), .A2(new_n557), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(G141gat), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n884), .B(new_n891), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NOR4_X1   g704(.A1(new_n886), .A2(G141gat), .A3(new_n445), .A4(new_n557), .ZN(new_n906));
  INV_X1    g705(.A(new_n900), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n698), .A3(new_n901), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n908), .B2(G141gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n909), .B2(new_n884), .ZN(G1344gat));
  AOI21_X1  g709(.A(KEYINPUT57), .B1(new_n897), .B2(new_n252), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n847), .A2(new_n848), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n898), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n655), .B(new_n901), .C1(new_n911), .C2(new_n913), .ZN(new_n914));
  AND2_X1   g713(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n902), .A2(KEYINPUT59), .A3(new_n656), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n914), .A2(new_n915), .B1(new_n907), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n888), .A2(new_n662), .A3(new_n890), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n655), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n920), .B2(G148gat), .ZN(G1345gat));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n214), .A3(new_n633), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n900), .A2(new_n712), .A3(new_n902), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n214), .B2(new_n923), .ZN(G1346gat));
  NAND2_X1  g723(.A1(new_n919), .A2(new_n708), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n900), .A2(new_n902), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n685), .A2(new_n215), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n925), .A2(new_n215), .B1(new_n926), .B2(new_n927), .ZN(G1347gat));
  NAND2_X1  g727(.A1(new_n445), .A2(new_n700), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n698), .A2(G169gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n858), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n929), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(new_n433), .A3(new_n437), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n849), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n698), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n931), .A2(new_n935), .ZN(G1348gat));
  INV_X1    g735(.A(G176gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n937), .A3(new_n655), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n858), .A2(new_n713), .A3(new_n929), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n937), .ZN(G1349gat));
  NAND4_X1  g739(.A1(new_n855), .A2(new_n633), .A3(new_n857), .A4(new_n932), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n260), .A2(new_n265), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g742(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n712), .A2(new_n311), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n933), .B(new_n945), .C1(new_n847), .C2(new_n848), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  AOI22_X1  g748(.A1(new_n948), .A2(new_n949), .B1(KEYINPUT126), .B2(KEYINPUT60), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n943), .A2(new_n944), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n944), .B1(new_n943), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n934), .A2(new_n306), .A3(new_n708), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n855), .A2(new_n708), .A3(new_n857), .A4(new_n932), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n955), .A2(new_n956), .A3(G190gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n955), .B2(G190gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  INV_X1    g758(.A(new_n893), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n706), .A2(new_n929), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n698), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n911), .A2(new_n913), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n961), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n698), .A2(G197gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1352gat));
  OAI21_X1  g768(.A(G204gat), .B1(new_n966), .B2(new_n713), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n656), .A2(G204gat), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT62), .B1(new_n962), .B2(new_n972), .ZN(new_n973));
  OR3_X1    g772(.A1(new_n962), .A2(KEYINPUT62), .A3(new_n972), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(G1353gat));
  INV_X1    g774(.A(G211gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n963), .A2(new_n976), .A3(new_n633), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n633), .B(new_n961), .C1(new_n911), .C2(new_n913), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT63), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n976), .B1(KEYINPUT127), .B2(new_n979), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n980), .B1(new_n978), .B2(new_n981), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n977), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  OAI21_X1  g783(.A(G218gat), .B1(new_n966), .B2(new_n685), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n963), .A2(new_n591), .A3(new_n708), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


