//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT81), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  INV_X1    g007(.A(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n191), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT2), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G116), .B(G119), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT66), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n196), .A2(new_n197), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT4), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G107), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT3), .A3(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G107), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n209), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n217), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n213), .A2(KEYINPUT3), .A3(G104), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n213), .B2(G104), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n209), .B(new_n216), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT4), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n222), .A2(KEYINPUT73), .A3(new_n217), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT73), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n213), .A2(G104), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(new_n212), .B2(new_n214), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n208), .B1(new_n226), .B2(new_n209), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G101), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n224), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n218), .B(KEYINPUT79), .C1(new_n223), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n199), .B1(new_n204), .B2(KEYINPUT5), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT80), .B1(new_n193), .B2(KEYINPUT5), .ZN(new_n233));
  OR3_X1    g047(.A1(new_n193), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n206), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT74), .B1(new_n213), .B2(G104), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n211), .A3(G107), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n213), .A2(G104), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G101), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n221), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n236), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n231), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT73), .B1(new_n222), .B2(new_n217), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n227), .A2(new_n229), .A3(new_n224), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT79), .B1(new_n248), .B2(new_n218), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n190), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n218), .B1(new_n223), .B2(new_n230), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT79), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n190), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n244), .A4(new_n231), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n250), .A2(KEYINPUT82), .A3(new_n255), .A4(KEYINPUT6), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n250), .A2(KEYINPUT6), .A3(new_n255), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n258), .B(new_n190), .C1(new_n245), .C2(new_n249), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n256), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G143), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(KEYINPUT1), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(G128), .ZN(new_n269));
  INV_X1    g083(.A(G128), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n264), .B(new_n266), .C1(KEYINPUT1), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G125), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n275));
  XNOR2_X1  g089(.A(G143), .B(G146), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT0), .B(G128), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  NOR2_X1   g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n267), .A2(new_n281), .A3(KEYINPUT64), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n264), .A2(new_n266), .A3(new_n279), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n276), .A2(KEYINPUT65), .A3(new_n279), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n278), .A2(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n274), .B1(new_n287), .B2(new_n273), .ZN(new_n288));
  INV_X1    g102(.A(G953), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n289), .A2(G224), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n288), .B(new_n290), .Z(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n262), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G210), .B1(G237), .B2(G902), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n236), .B(new_n243), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n190), .B(KEYINPUT8), .Z(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT7), .ZN(new_n298));
  OR3_X1    g112(.A1(new_n288), .A2(new_n298), .A3(new_n290), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n288), .B1(new_n298), .B2(new_n290), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n301), .B2(new_n255), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n293), .A2(new_n294), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n294), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n250), .A2(KEYINPUT6), .A3(new_n255), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n260), .A3(new_n259), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n291), .B1(new_n306), .B2(new_n256), .ZN(new_n307));
  INV_X1    g121(.A(new_n302), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n188), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT78), .B(G469), .ZN(new_n312));
  XNOR2_X1  g126(.A(G110), .B(G140), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n289), .A2(G227), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n278), .A2(new_n282), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n285), .A2(new_n286), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n228), .A2(new_n208), .A3(G101), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n223), .B2(new_n230), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT11), .ZN(new_n321));
  INV_X1    g135(.A(G134), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(G137), .ZN(new_n323));
  INV_X1    g137(.A(G137), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT11), .A3(G134), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(G137), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G131), .ZN(new_n328));
  INV_X1    g142(.A(G131), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n323), .A2(new_n325), .A3(new_n329), .A4(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n328), .A2(KEYINPUT67), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n269), .A2(new_n271), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT10), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n221), .A4(new_n242), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n242), .A2(new_n221), .A3(new_n269), .A4(new_n271), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT10), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n320), .A2(new_n336), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n320), .A2(KEYINPUT75), .A3(new_n336), .A4(new_n342), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n315), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n243), .A2(new_n272), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n340), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT12), .A3(new_n331), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n351));
  AOI211_X1 g165(.A(new_n351), .B(KEYINPUT12), .C1(new_n349), .C2(new_n335), .ZN(new_n352));
  INV_X1    g166(.A(new_n340), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n242), .A2(new_n221), .B1(new_n269), .B2(new_n271), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n328), .A2(KEYINPUT67), .A3(new_n330), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT67), .B1(new_n328), .B2(new_n330), .ZN(new_n356));
  OAI22_X1  g170(.A1(new_n353), .A2(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT12), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT76), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n350), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n347), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n315), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n345), .A2(new_n346), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n320), .A2(new_n342), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n335), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n311), .B(new_n312), .C1(new_n361), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n363), .A2(new_n368), .A3(new_n360), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n363), .B2(new_n360), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n315), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n347), .A2(new_n365), .ZN(new_n372));
  AOI21_X1  g186(.A(G902), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G469), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n367), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G221), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT9), .B(G234), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n378), .B2(new_n311), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G952), .ZN(new_n381));
  AOI211_X1 g195(.A(G953), .B(new_n381), .C1(G234), .C2(G237), .ZN(new_n382));
  AOI211_X1 g196(.A(new_n311), .B(new_n289), .C1(G234), .C2(G237), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT21), .B(G898), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G475), .ZN(new_n387));
  NOR2_X1   g201(.A1(G237), .A2(G953), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G214), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT83), .A3(new_n265), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n265), .A2(KEYINPUT83), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(G214), .A3(new_n388), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n329), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G125), .B(G140), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT16), .ZN(new_n398));
  INV_X1    g212(.A(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G125), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(KEYINPUT16), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n263), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n398), .B(G146), .C1(KEYINPUT16), .C2(new_n400), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n393), .A2(KEYINPUT17), .A3(G131), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT72), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n273), .A2(G140), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n399), .A2(G125), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n273), .A2(G140), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n410), .A3(KEYINPUT72), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n263), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n263), .B2(new_n397), .ZN(new_n413));
  NAND2_X1  g227(.A1(KEYINPUT18), .A2(G131), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n393), .B(new_n414), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n396), .A2(new_n405), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G113), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT86), .B(G104), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n416), .B(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n387), .B1(new_n421), .B2(new_n311), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT87), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n416), .B2(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n415), .A2(new_n413), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT19), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n409), .A2(new_n427), .A3(new_n411), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT19), .B1(new_n407), .B2(new_n408), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n263), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n428), .A2(KEYINPUT84), .A3(new_n263), .A4(new_n429), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n403), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n394), .B1(new_n434), .B2(KEYINPUT85), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT85), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n432), .A2(new_n436), .A3(new_n403), .A4(new_n433), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n426), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n424), .B1(new_n438), .B2(new_n420), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n430), .A2(new_n431), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n403), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT85), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n394), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n437), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n425), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n423), .A3(new_n419), .ZN(new_n446));
  NOR2_X1   g260(.A1(G475), .A2(G902), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n439), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n422), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT88), .B(G122), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(new_n194), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n194), .A2(G122), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT14), .ZN(new_n456));
  OR3_X1    g270(.A1(new_n455), .A2(KEYINPUT90), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT90), .B1(new_n455), .B2(new_n456), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n454), .A2(KEYINPUT14), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT91), .ZN(new_n461));
  OAI21_X1  g275(.A(G107), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n453), .A2(new_n213), .A3(new_n454), .ZN(new_n463));
  XNOR2_X1  g277(.A(G128), .B(G143), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n322), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G107), .B1(new_n452), .B2(new_n455), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT13), .B1(new_n270), .B2(G143), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(new_n322), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n464), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n468), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n469), .B1(new_n468), .B2(new_n472), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G217), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n377), .A2(new_n476), .A3(G953), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n466), .B(new_n477), .C1(new_n473), .C2(new_n474), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  AOI211_X1 g299(.A(G902), .B(new_n483), .C1(new_n479), .C2(new_n480), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n439), .A2(new_n446), .A3(KEYINPUT20), .A4(new_n447), .ZN(new_n488));
  AND4_X1   g302(.A1(new_n386), .A2(new_n450), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n310), .A2(new_n375), .A3(new_n380), .A4(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT70), .ZN(new_n491));
  NOR2_X1   g305(.A1(G472), .A2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n287), .B1(new_n355), .B2(new_n356), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n322), .A2(G137), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n324), .A2(G134), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n330), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n271), .A3(new_n269), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(KEYINPUT30), .A3(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n276), .A2(new_n277), .A3(new_n275), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT64), .B1(new_n267), .B2(new_n281), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT65), .B1(new_n276), .B2(new_n279), .ZN(new_n503));
  AND4_X1   g317(.A1(KEYINPUT65), .A2(new_n264), .A3(new_n266), .A4(new_n279), .ZN(new_n504));
  OAI22_X1  g318(.A1(new_n501), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n328), .A2(new_n330), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n206), .A2(new_n207), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n500), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n388), .A2(G210), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT27), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT26), .B(G101), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n510), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n494), .A2(new_n516), .A3(new_n499), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT31), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n511), .A2(new_n520), .A3(new_n515), .A4(new_n517), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n515), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT68), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n287), .A2(new_n331), .B1(new_n337), .B2(new_n498), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n516), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n507), .A2(KEYINPUT68), .A3(new_n510), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n517), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n528), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n517), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n528), .A2(KEYINPUT28), .B1(new_n531), .B2(KEYINPUT69), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n523), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n493), .B1(new_n522), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n491), .B1(new_n534), .B2(KEYINPUT32), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n528), .A2(KEYINPUT28), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(KEYINPUT69), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n528), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n515), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n519), .A2(new_n521), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n492), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT32), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(KEYINPUT70), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n534), .A2(KEYINPUT32), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n511), .A2(new_n517), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n523), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n529), .A2(new_n532), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n515), .ZN(new_n551));
  INV_X1    g365(.A(new_n517), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n516), .B1(new_n494), .B2(new_n499), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT28), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n523), .A2(new_n548), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n531), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n311), .ZN(new_n557));
  OAI21_X1  g371(.A(G472), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n535), .A2(new_n544), .A3(new_n545), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n476), .B1(G234), .B2(new_n311), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n402), .A2(new_n403), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n192), .A2(G128), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n563), .A2(KEYINPUT23), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n270), .A2(G119), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(KEYINPUT71), .A2(KEYINPUT23), .ZN(new_n568));
  OAI22_X1  g382(.A1(new_n564), .A2(new_n567), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G110), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n563), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT24), .B(G110), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n562), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n574), .B1(new_n569), .B2(G110), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n412), .A3(new_n403), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n289), .A2(G221), .A3(G234), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n578), .B(new_n579), .Z(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n573), .A2(new_n576), .A3(new_n580), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(KEYINPUT25), .A3(new_n311), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n311), .A3(new_n583), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT25), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n561), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n560), .A2(G902), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n559), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n490), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT92), .B(G101), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G3));
  OAI21_X1  g410(.A(new_n311), .B1(new_n540), .B2(new_n541), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n534), .B1(G472), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n375), .A2(new_n592), .A3(new_n380), .A4(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT94), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n448), .A2(new_n449), .ZN(new_n601));
  INV_X1    g415(.A(new_n422), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n488), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n479), .A2(new_n480), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT33), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n479), .A2(new_n607), .A3(new_n480), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(G478), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n482), .A2(new_n311), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n481), .B2(new_n482), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n603), .A2(new_n604), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n604), .B1(new_n603), .B2(new_n612), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n294), .B1(new_n293), .B2(new_n302), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n307), .A2(new_n304), .A3(new_n308), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n187), .B(new_n386), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n600), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n603), .A2(new_n612), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT93), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n603), .A2(new_n604), .A3(new_n612), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI211_X1 g437(.A(new_n188), .B(new_n385), .C1(new_n303), .C2(new_n309), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT94), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n599), .B1(new_n619), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT34), .B(G104), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NAND2_X1  g442(.A1(new_n303), .A2(new_n309), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n603), .A2(new_n487), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n187), .A4(new_n386), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT95), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n310), .A2(KEYINPUT95), .A3(new_n386), .A4(new_n630), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n599), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT35), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n585), .A2(new_n588), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n560), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n577), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n590), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n638), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n643), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n589), .A2(KEYINPUT96), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n598), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n490), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT37), .B(G110), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  AND3_X1   g465(.A1(new_n310), .A2(new_n380), .A3(new_n375), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n559), .A2(new_n647), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n481), .B(new_n484), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n383), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n382), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n450), .A2(new_n655), .A3(new_n488), .A4(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XNOR2_X1  g477(.A(new_n629), .B(KEYINPUT38), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n187), .B1(new_n485), .B2(new_n486), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n450), .B2(new_n488), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n640), .A2(new_n643), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT97), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n546), .A2(new_n515), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n552), .A2(new_n553), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n671), .B(new_n311), .C1(new_n515), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n535), .A2(new_n544), .A3(new_n545), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n668), .A2(KEYINPUT97), .A3(new_n669), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n665), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n375), .A2(new_n380), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n659), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n678), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  NAND3_X1  g499(.A1(new_n603), .A2(new_n612), .A3(new_n659), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n654), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NAND2_X1  g503(.A1(new_n363), .A2(new_n365), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n690), .A2(new_n315), .B1(new_n347), .B2(new_n360), .ZN(new_n691));
  OAI21_X1  g505(.A(G469), .B1(new_n691), .B2(G902), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n380), .A3(new_n367), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n559), .A2(new_n592), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n615), .A2(new_n600), .A3(new_n618), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT94), .B1(new_n623), .B2(new_n624), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT98), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n619), .A2(new_n625), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT98), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n702), .A3(new_n696), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT99), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n704), .B(new_n706), .ZN(G15));
  AOI21_X1  g521(.A(new_n695), .B1(new_n633), .B2(new_n634), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n194), .ZN(G18));
  NAND2_X1  g523(.A1(new_n559), .A2(new_n647), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n310), .A2(new_n694), .ZN(new_n711));
  INV_X1    g525(.A(new_n489), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n192), .ZN(G21));
  NOR2_X1   g528(.A1(new_n693), .A2(new_n385), .ZN(new_n715));
  AOI21_X1  g529(.A(G902), .B1(new_n522), .B2(new_n533), .ZN(new_n716));
  INV_X1    g530(.A(G472), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT100), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT100), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n597), .A2(new_n719), .A3(G472), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n554), .A2(new_n531), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n515), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n492), .B1(new_n723), .B2(new_n541), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n715), .A2(new_n721), .A3(new_n592), .A4(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n629), .A2(new_n726), .A3(new_n667), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n667), .B1(new_n616), .B2(new_n617), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT101), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n725), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n730), .B(G122), .Z(G24));
  NAND3_X1  g545(.A1(new_n721), .A2(new_n669), .A3(new_n724), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n686), .ZN(new_n733));
  INV_X1    g547(.A(new_n711), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n303), .A2(new_n309), .A3(new_n187), .ZN(new_n738));
  NAND2_X1  g552(.A1(G469), .A2(G902), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT102), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n690), .A2(new_n315), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n347), .A2(new_n360), .ZN(new_n742));
  AOI21_X1  g556(.A(G902), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n740), .B1(new_n743), .B2(new_n312), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n371), .A2(G469), .A3(new_n372), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n379), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n738), .A2(new_n559), .A3(new_n592), .A4(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n737), .B1(new_n747), .B2(new_n686), .ZN(new_n748));
  AND4_X1   g562(.A1(KEYINPUT42), .A2(new_n603), .A3(new_n612), .A4(new_n659), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n738), .A2(new_n749), .A3(new_n746), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n534), .B2(KEYINPUT32), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n542), .A2(KEYINPUT103), .A3(new_n543), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n545), .A4(new_n558), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n592), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT104), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n592), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n538), .A2(new_n515), .A3(new_n539), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT29), .B1(new_n546), .B2(new_n523), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n557), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI22_X1  g574(.A1(new_n542), .A2(new_n543), .B1(new_n760), .B2(new_n717), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT103), .B1(new_n542), .B2(new_n543), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n757), .B1(new_n763), .B2(new_n753), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n363), .A2(new_n360), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT77), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n363), .A2(new_n360), .A3(new_n368), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n362), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n372), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n768), .A2(new_n374), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n740), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n367), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n380), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n303), .A2(new_n309), .A3(new_n187), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT104), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n764), .A2(new_n775), .A3(new_n776), .A4(new_n749), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n748), .A2(new_n756), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  INV_X1    g593(.A(KEYINPUT105), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n660), .B(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT106), .B1(new_n747), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n559), .A2(new_n592), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n660), .B(KEYINPUT105), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n775), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  INV_X1    g602(.A(new_n598), .ZN(new_n789));
  INV_X1    g603(.A(new_n603), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n612), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT43), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n793), .A3(new_n612), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n789), .B(new_n669), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n768), .B2(new_n769), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n371), .A2(KEYINPUT45), .A3(new_n372), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(G469), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT107), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n805), .A3(KEYINPUT46), .A4(new_n771), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n804), .A2(new_n771), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n367), .B(new_n806), .C1(new_n807), .C2(KEYINPUT46), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(KEYINPUT46), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n380), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n680), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n798), .A2(new_n799), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n800), .A2(new_n738), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  XNOR2_X1  g629(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n380), .B(new_n816), .C1(new_n808), .C2(new_n809), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n559), .A2(new_n774), .A3(new_n592), .A4(new_n686), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  NAND2_X1  g637(.A1(new_n738), .A2(new_n694), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n824), .A2(new_n675), .A3(new_n757), .A4(new_n658), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n381), .B(G953), .C1(new_n825), .C2(new_n623), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT114), .B1(new_n795), .B2(new_n658), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n792), .A2(new_n828), .A3(new_n382), .A4(new_n794), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n824), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(KEYINPUT119), .A3(KEYINPUT48), .A4(new_n764), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n830), .A2(new_n764), .ZN(new_n832));
  XNOR2_X1  g646(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n826), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n721), .A2(new_n592), .A3(new_n724), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n827), .B2(new_n829), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n734), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(KEYINPUT118), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n834), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n732), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n603), .A2(new_n612), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n830), .A2(new_n841), .B1(new_n825), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n664), .A2(new_n187), .A3(new_n693), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n836), .A2(KEYINPUT50), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT50), .B1(new_n836), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n827), .A2(new_n829), .ZN(new_n848));
  INV_X1    g662(.A(new_n835), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n738), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n692), .A2(new_n367), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT111), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(new_n380), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n818), .A2(new_n819), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n847), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n840), .B1(new_n857), .B2(KEYINPUT51), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(KEYINPUT116), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n818), .A2(new_n860), .A3(new_n819), .A4(new_n855), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n852), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(KEYINPUT51), .B(new_n843), .C1(new_n845), .C2(new_n846), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n862), .A2(KEYINPUT117), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT117), .B1(new_n862), .B2(new_n864), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n858), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n708), .A2(new_n730), .A3(new_n713), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n702), .B1(new_n701), .B2(new_n696), .ZN(new_n869));
  AOI211_X1 g683(.A(KEYINPUT98), .B(new_n695), .C1(new_n619), .C2(new_n625), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n490), .B1(new_n593), .B2(new_n648), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n620), .B1(new_n487), .B2(new_n603), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(new_n310), .A3(new_n386), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n599), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n603), .A2(new_n655), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n375), .A2(new_n380), .A3(new_n877), .A4(new_n659), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n774), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n879), .A2(new_n653), .B1(new_n733), .B2(new_n775), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n778), .A2(new_n876), .A3(new_n787), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT112), .B1(new_n871), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n715), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n835), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n729), .A2(new_n727), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n559), .A2(new_n489), .A3(new_n647), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n884), .A2(new_n885), .B1(new_n886), .B2(new_n734), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n633), .A2(new_n634), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n696), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n700), .B2(new_n703), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n778), .A2(new_n876), .A3(new_n787), .A4(new_n880), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT112), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n882), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n652), .B(new_n653), .C1(new_n661), .C2(new_n687), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n640), .A2(new_n643), .A3(new_n659), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n773), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n727), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n726), .B1(new_n629), .B2(new_n667), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n675), .B(new_n899), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n897), .A2(new_n735), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT113), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n897), .A2(new_n902), .A3(new_n735), .A4(KEYINPUT113), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT52), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n903), .A2(KEYINPUT52), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n895), .A2(new_n896), .A3(new_n909), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n905), .A2(KEYINPUT52), .A3(new_n906), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n907), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n893), .B1(new_n891), .B2(new_n892), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n871), .A2(KEYINPUT112), .A3(new_n881), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  OAI211_X1 g730(.A(KEYINPUT54), .B(new_n910), .C1(new_n916), .C2(new_n896), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n896), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n871), .A2(new_n881), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n909), .A2(KEYINPUT53), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n867), .A2(new_n924), .B1(G952), .B2(G953), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n854), .B(KEYINPUT49), .Z(new_n926));
  NAND3_X1  g740(.A1(new_n592), .A2(new_n187), .A3(new_n380), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT110), .Z(new_n928));
  NOR3_X1   g742(.A1(new_n928), .A2(new_n675), .A3(new_n791), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n926), .A2(new_n665), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(G75));
  XNOR2_X1  g745(.A(new_n262), .B(new_n292), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT53), .B1(new_n895), .B2(new_n912), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n920), .ZN(new_n938));
  NAND2_X1  g752(.A1(G210), .A2(G902), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n289), .A2(G952), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT123), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n918), .A2(new_n921), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(KEYINPUT121), .A3(G210), .A4(G902), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n938), .B2(new_n939), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT56), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n943), .B1(new_n949), .B2(new_n934), .ZN(G51));
  XNOR2_X1  g764(.A(new_n740), .B(KEYINPUT57), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n922), .B1(new_n918), .B2(new_n921), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n937), .A2(new_n920), .A3(KEYINPUT54), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n691), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n804), .ZN(new_n957));
  OAI211_X1 g771(.A(G902), .B(new_n957), .C1(new_n937), .C2(new_n920), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n941), .B1(new_n956), .B2(new_n960), .ZN(G54));
  NAND4_X1  g775(.A1(new_n944), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n439), .A2(new_n446), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n941), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n938), .A2(new_n311), .ZN(new_n965));
  INV_X1    g779(.A(new_n963), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(KEYINPUT58), .A3(G475), .A4(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n964), .A2(new_n967), .ZN(G60));
  NAND2_X1  g782(.A1(new_n606), .A2(new_n608), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n610), .B(KEYINPUT59), .Z(new_n970));
  OAI211_X1 g784(.A(new_n969), .B(new_n970), .C1(new_n952), .C2(new_n953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n942), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n924), .B2(new_n970), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G63));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n642), .B(new_n977), .C1(new_n937), .C2(new_n920), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n918), .B2(new_n921), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n942), .B(new_n978), .C1(new_n979), .C2(new_n584), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n584), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n938), .B2(new_n976), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n984), .A2(KEYINPUT61), .A3(new_n942), .A4(new_n978), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(new_n985), .ZN(G66));
  INV_X1    g800(.A(new_n384), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n289), .B1(new_n987), .B2(G224), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n891), .A2(new_n876), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(new_n289), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n306), .B(new_n256), .C1(G898), .C2(new_n289), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT125), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n990), .B(new_n992), .ZN(G69));
  NAND2_X1  g807(.A1(new_n814), .A2(new_n822), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n812), .A2(new_n885), .A3(new_n764), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n897), .A2(new_n735), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n995), .A2(new_n778), .A3(new_n787), .A4(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n289), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n500), .A2(new_n509), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT126), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n428), .A2(new_n429), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n999), .B(new_n1003), .C1(new_n656), .C2(new_n289), .ZN(new_n1004));
  INV_X1    g818(.A(new_n994), .ZN(new_n1005));
  INV_X1    g819(.A(new_n681), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1006), .A2(new_n783), .A3(new_n738), .A4(new_n873), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n684), .A2(new_n996), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n684), .A2(KEYINPUT62), .A3(new_n996), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1005), .A2(KEYINPUT127), .A3(new_n1007), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1007), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1014), .B1(new_n1015), .B2(new_n994), .ZN(new_n1016));
  AOI21_X1  g830(.A(G953), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1004), .B1(new_n1017), .B2(new_n1003), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n289), .B1(G227), .B2(G900), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1019), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n1004), .B(new_n1021), .C1(new_n1017), .C2(new_n1003), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1020), .A2(new_n1022), .ZN(G72));
  INV_X1    g837(.A(new_n989), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1013), .A2(new_n1024), .A3(new_n1016), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  AOI21_X1  g841(.A(new_n671), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n910), .B1(new_n916), .B2(new_n896), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n511), .A2(new_n523), .A3(new_n517), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n671), .A2(new_n1030), .A3(new_n1027), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n998), .A2(new_n1024), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1030), .B1(new_n1033), .B2(new_n1027), .ZN(new_n1034));
  NOR4_X1   g848(.A1(new_n1028), .A2(new_n1032), .A3(new_n1034), .A4(new_n941), .ZN(G57));
endmodule


