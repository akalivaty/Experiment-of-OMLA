//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n578, new_n579, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G137), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n462), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G113), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n464), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n460), .A2(new_n461), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n460), .B2(new_n461), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n496), .B(new_n499), .C1(new_n461), .C2(new_n460), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(KEYINPUT67), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(KEYINPUT67), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n508), .A2(G88), .B1(new_n509), .B2(G50), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  AND3_X1   g086(.A1(KEYINPUT67), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(G543), .B1(KEYINPUT67), .B2(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(G62), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(new_n515), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n504), .B2(new_n505), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT68), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n511), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n510), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n523), .B1(new_n518), .B2(KEYINPUT68), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n514), .A2(new_n515), .ZN(new_n525));
  OAI21_X1  g100(.A(G651), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(KEYINPUT69), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(G166));
  NAND2_X1  g103(.A1(new_n509), .A2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n504), .A2(new_n505), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n508), .A2(G89), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n536));
  OR3_X1    g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n534), .B2(new_n535), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n511), .ZN(new_n541));
  INV_X1    g116(.A(new_n507), .ZN(new_n542));
  NOR2_X1   g117(.A1(KEYINPUT6), .A2(G651), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n512), .A2(new_n513), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI21_X1  g120(.A(G543), .B1(new_n542), .B2(new_n543), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n541), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n530), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n511), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n544), .A2(new_n552), .B1(new_n546), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT73), .ZN(new_n560));
  XOR2_X1   g135(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n561));
  XNOR2_X1  g136(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n509), .A2(G53), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n511), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n508), .A2(G91), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT74), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n565), .A2(new_n572), .A3(new_n567), .A4(new_n568), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  AND2_X1   g151(.A1(new_n537), .A2(new_n538), .ZN(G286));
  NAND2_X1  g152(.A1(new_n520), .A2(new_n521), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n526), .A2(KEYINPUT69), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(new_n579), .A3(new_n510), .ZN(G303));
  AOI22_X1  g155(.A1(new_n508), .A2(G87), .B1(new_n509), .B2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n508), .A2(G86), .B1(new_n509), .B2(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT75), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n504), .B2(new_n505), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n584), .A2(new_n589), .ZN(G305));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n544), .A2(new_n591), .B1(new_n546), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI221_X1 g170(.A(KEYINPUT76), .B1(new_n546), .B2(new_n592), .C1(new_n544), .C2(new_n591), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n530), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n597), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n508), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT10), .Z(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n599), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n509), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n604), .B1(new_n611), .B2(G868), .ZN(G321));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(G286), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n614), .ZN(G297));
  AOI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(new_n614), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n611), .B1(new_n619), .B2(G860), .ZN(G148));
  INV_X1    g195(.A(new_n555), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n614), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n611), .A2(new_n619), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n624), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n480), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n483), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n482), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT77), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2096), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT3), .B(G2104), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(new_n465), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n633), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT79), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(KEYINPUT80), .B(KEYINPUT18), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n660), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n663), .B2(new_n659), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT81), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT81), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n673), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n674), .A2(new_n675), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(new_n677), .ZN(new_n683));
  MUX2_X1   g258(.A(new_n683), .B(new_n682), .S(new_n673), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G229));
  MUX2_X1   g266(.A(G6), .B(G305), .S(G16), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT32), .ZN(new_n693));
  INV_X1    g268(.A(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(G166), .A2(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G16), .B2(G22), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n695), .A2(new_n699), .A3(new_n700), .A4(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G24), .ZN(new_n710));
  INV_X1    g285(.A(G290), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT83), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT82), .B(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n480), .A2(G131), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n483), .A2(G119), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n482), .A2(G107), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n708), .A2(new_n709), .A3(new_n715), .A4(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT36), .Z(new_n725));
  XOR2_X1   g300(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(G29), .B1(new_n727), .B2(G34), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G34), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(G160), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2084), .ZN(new_n732));
  NOR2_X1   g307(.A1(G29), .A2(G33), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT86), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G139), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT87), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n634), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n737));
  NAND2_X1  g312(.A1(G103), .A2(G2104), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G2105), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(KEYINPUT25), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT25), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n738), .A2(new_n741), .A3(G2105), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n736), .B1(new_n482), .B2(new_n737), .C1(new_n740), .C2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n734), .B1(new_n743), .B2(new_n730), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G2072), .Z(new_n745));
  INV_X1    g320(.A(G1348), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n611), .A2(new_n701), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G4), .B2(new_n701), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n732), .B(new_n745), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n730), .A2(G32), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n483), .A2(G129), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n480), .A2(G141), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n465), .A2(G105), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n750), .B1(new_n758), .B2(new_n730), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT27), .B(G1996), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT89), .Z(new_n762));
  XOR2_X1   g337(.A(KEYINPUT31), .B(G11), .Z(new_n763));
  INV_X1    g338(.A(G28), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(KEYINPUT30), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT91), .ZN(new_n766));
  AOI21_X1  g341(.A(G29), .B1(new_n764), .B2(KEYINPUT30), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n631), .B2(new_n730), .ZN(new_n769));
  NOR2_X1   g344(.A1(G27), .A2(G29), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G164), .B2(G29), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n769), .B1(G2078), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(G2078), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n759), .B2(new_n760), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n762), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n701), .A2(G5), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G171), .B2(new_n701), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1961), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n748), .A2(new_n746), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n775), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n749), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT93), .B(KEYINPUT23), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n701), .A2(G20), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n616), .B2(new_n701), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1956), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n730), .A2(G26), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT85), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n480), .A2(G140), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n483), .A2(G128), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n482), .A2(G116), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT84), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(G29), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2067), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n730), .A2(G35), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT92), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G162), .B2(new_n730), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT29), .B(G2090), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n701), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n555), .B2(new_n701), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n802), .B1(G1341), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n797), .B(new_n805), .C1(G1341), .C2(new_n804), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G21), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G168), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT90), .B(G1966), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n781), .A2(new_n786), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n725), .A2(new_n812), .ZN(G311));
  INV_X1    g388(.A(G311), .ZN(G150));
  NAND2_X1  g389(.A1(new_n611), .A2(G559), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT38), .Z(new_n816));
  AOI22_X1  g391(.A1(new_n508), .A2(G93), .B1(new_n509), .B2(G55), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n530), .A2(G67), .ZN(new_n818));
  NAND2_X1  g393(.A1(G80), .A2(G543), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n511), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT94), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g397(.A(KEYINPUT94), .B(new_n511), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n621), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT95), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n621), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n816), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n832));
  AOI21_X1  g407(.A(G860), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  OAI21_X1  g409(.A(G860), .B1(new_n822), .B2(new_n823), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  NAND2_X1  g412(.A1(new_n483), .A2(G130), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n482), .A2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G142), .B2(new_n480), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n636), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n720), .ZN(new_n844));
  INV_X1    g419(.A(new_n795), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n743), .B(new_n758), .ZN(new_n847));
  INV_X1    g422(.A(new_n500), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n499), .B1(new_n634), .B2(new_n496), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n489), .B(new_n493), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT97), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n498), .A2(new_n500), .ZN(new_n852));
  INV_X1    g427(.A(new_n494), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n847), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n846), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n477), .B(new_n631), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n487), .ZN(new_n860));
  AOI21_X1  g435(.A(G37), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(new_n860), .B2(new_n858), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n711), .B(G303), .ZN(new_n865));
  XNOR2_X1  g440(.A(G305), .B(G288), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G303), .B(G290), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n871), .B1(KEYINPUT100), .B2(KEYINPUT42), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n623), .B1(new_n826), .B2(new_n829), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n611), .A2(new_n570), .A3(new_n573), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n611), .B1(new_n573), .B2(new_n570), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n611), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n571), .B2(new_n574), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n879), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n826), .A2(new_n623), .A3(new_n829), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n877), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n879), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n826), .A2(new_n623), .A3(new_n829), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(new_n876), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT99), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n877), .A2(new_n888), .A3(new_n895), .A4(new_n889), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n875), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n894), .A2(new_n896), .B1(new_n874), .B2(new_n873), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n875), .A2(new_n894), .A3(KEYINPUT101), .A4(new_n896), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(G868), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n824), .A2(G868), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n864), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n614), .B1(new_n900), .B2(new_n901), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n907), .A2(KEYINPUT102), .A3(new_n904), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(G295));
  OR3_X1    g484(.A1(new_n907), .A2(KEYINPUT103), .A3(new_n904), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT103), .B1(new_n907), .B2(new_n904), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(G331));
  NAND2_X1  g487(.A1(G286), .A2(KEYINPUT105), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n914));
  NAND2_X1  g489(.A1(G168), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G171), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(G301), .A3(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n919), .A2(new_n830), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n830), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT106), .B1(new_n891), .B2(new_n878), .ZN(new_n922));
  OR3_X1    g497(.A1(new_n891), .A2(KEYINPUT106), .A3(new_n878), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n921), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n919), .A2(new_n830), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n891), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n891), .A2(new_n885), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n870), .A3(new_n868), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n920), .A2(new_n888), .A3(new_n921), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n932), .A3(new_n871), .ZN(new_n933));
  XOR2_X1   g508(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n934));
  NAND4_X1  g509(.A1(new_n930), .A2(new_n931), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  INV_X1    g511(.A(new_n934), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n931), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n871), .B1(new_n927), .B2(new_n932), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n935), .A2(new_n936), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n920), .A2(new_n921), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n891), .B1(new_n942), .B2(new_n885), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n871), .B1(new_n943), .B2(new_n924), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n944), .B2(new_n938), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(KEYINPUT43), .C1(new_n944), .C2(new_n938), .ZN(new_n948));
  OR3_X1    g523(.A1(new_n938), .A2(new_n939), .A3(new_n937), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n941), .B1(new_n950), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n851), .A2(new_n952), .A3(new_n855), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G40), .ZN(new_n956));
  OAI22_X1  g531(.A1(new_n479), .A2(new_n470), .B1(new_n474), .B2(new_n464), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(G2105), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n482), .A2(G137), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n471), .B2(new_n472), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n482), .A2(G101), .A3(G2104), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT66), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n958), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G2067), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n795), .B(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT109), .ZN(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n758), .B(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n722), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n720), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n845), .A2(new_n967), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n966), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT127), .ZN(new_n978));
  INV_X1    g553(.A(new_n758), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n965), .B1(new_n969), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n966), .B2(G1996), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n965), .A2(KEYINPUT46), .A3(new_n970), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  XOR2_X1   g559(.A(new_n984), .B(KEYINPUT47), .Z(new_n985));
  NOR2_X1   g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n965), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT48), .Z(new_n988));
  XNOR2_X1  g563(.A(new_n720), .B(new_n722), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n972), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n990), .B2(new_n965), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n978), .A2(new_n985), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT126), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n965), .ZN(new_n994));
  INV_X1    g569(.A(new_n986), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n996));
  NAND2_X1  g571(.A1(G290), .A2(G1986), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n998), .B(new_n965), .C1(new_n996), .C2(new_n997), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT55), .B(G8), .C1(new_n522), .C2(new_n527), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT111), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(G166), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n1006));
  NAND4_X1  g581(.A1(G303), .A2(new_n1006), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1002), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n954), .A2(G1384), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n851), .A2(new_n855), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n850), .A2(new_n952), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n954), .ZN(new_n1012));
  AND4_X1   g587(.A1(G40), .A2(new_n962), .A3(new_n476), .A4(new_n963), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n698), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n852), .B2(new_n853), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n1013), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1016), .B1(new_n1021), .B2(G2090), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n964), .B1(KEYINPUT50), .B2(new_n1011), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(KEYINPUT110), .A3(new_n1024), .A4(new_n1019), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1015), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1008), .A2(new_n1026), .A3(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n584), .A2(new_n589), .A3(new_n694), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n694), .B1(new_n584), .B2(new_n589), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G305), .A2(G1981), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(KEYINPUT49), .A3(new_n1029), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1004), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1037), .B(new_n1038), .C1(new_n703), .C2(G1976), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1976), .B1(new_n581), .B2(new_n582), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT114), .B1(new_n1040), .B2(KEYINPUT52), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(G288), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n581), .A2(KEYINPUT112), .A3(G1976), .A4(new_n582), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1043), .A2(new_n1046), .A3(G8), .A4(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1036), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1027), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1966), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1009), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n469), .B(new_n958), .C1(G164), .C2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT45), .B1(new_n850), .B2(new_n952), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT117), .ZN(new_n1061));
  INV_X1    g636(.A(G2084), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1019), .A2(new_n1020), .A3(new_n1062), .A4(new_n1013), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(new_n1056), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(G8), .A3(G168), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT63), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1026), .A2(G8), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1055), .B(new_n1069), .C1(new_n1008), .C2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT115), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n1073));
  NOR4_X1   g648(.A1(G164), .A2(new_n1073), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1023), .B(new_n1024), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1015), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1004), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1015), .A2(new_n1075), .A3(KEYINPUT116), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1008), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1027), .A2(new_n1054), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n1067), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1071), .B1(new_n1082), .B2(KEYINPUT63), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1027), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1036), .A2(new_n1045), .A3(new_n703), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1029), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1084), .A2(new_n1054), .B1(new_n1035), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n1090));
  INV_X1    g665(.A(G2078), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1010), .A2(new_n1012), .A3(new_n1091), .A4(new_n1013), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(G2078), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n955), .A2(new_n1013), .A3(new_n1095), .A4(new_n1010), .ZN(new_n1096));
  INV_X1    g671(.A(G1961), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1021), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1092), .A2(new_n1093), .B1(new_n1097), .B2(new_n1021), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n850), .A2(new_n1009), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1012), .A2(new_n1013), .A3(new_n1102), .A4(new_n1095), .ZN(new_n1103));
  AOI21_X1  g678(.A(G301), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1090), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1090), .B1(new_n1099), .B2(G171), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1101), .A2(G301), .A3(new_n1103), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT125), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1099), .A2(G171), .ZN(new_n1109));
  AND4_X1   g684(.A1(KEYINPUT125), .A2(new_n1109), .A3(KEYINPUT54), .A4(new_n1107), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1089), .B(new_n1105), .C1(new_n1108), .C2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1020), .A2(new_n1013), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1019), .A2(new_n1073), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1017), .A2(KEYINPUT115), .A3(new_n1018), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1113), .B1(new_n1117), .B2(G1956), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n565), .A2(new_n567), .A3(new_n568), .A4(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1122), .B(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1118), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1021), .A2(new_n746), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1043), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n967), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1021), .A2(new_n746), .B1(new_n1129), .B2(new_n967), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT119), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1127), .B1(new_n1136), .B2(new_n883), .ZN(new_n1137));
  INV_X1    g712(.A(G1956), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(new_n1114), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n1125), .A3(new_n1113), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n883), .B1(new_n1136), .B2(KEYINPUT60), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1134), .A2(KEYINPUT119), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1128), .A2(new_n1130), .A3(KEYINPUT119), .ZN(new_n1145));
  OR3_X1    g720(.A1(new_n1144), .A2(new_n1145), .A3(KEYINPUT60), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1010), .A2(new_n1012), .A3(new_n970), .A4(new_n1013), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT58), .B(G1341), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n1043), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n621), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1150), .B2(KEYINPUT120), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1143), .A2(new_n1146), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1127), .A2(KEYINPUT61), .A3(new_n1141), .ZN(new_n1157));
  OAI211_X1 g732(.A(KEYINPUT60), .B(new_n883), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1141), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1125), .B1(new_n1140), .B2(new_n1113), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(KEYINPUT121), .B(new_n1161), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1156), .A2(new_n1160), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1111), .B1(new_n1142), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1065), .A2(new_n1063), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1102), .B(new_n1013), .C1(KEYINPUT45), .C2(new_n1017), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1064), .B1(new_n1172), .B2(new_n1056), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1170), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(G168), .A2(new_n1004), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1061), .A2(KEYINPUT122), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1066), .A2(G8), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT51), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1178), .B(new_n1179), .C1(new_n1004), .C2(G168), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1174), .A2(G8), .A3(new_n1176), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1175), .B(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1179), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1180), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g761(.A(KEYINPUT124), .B(new_n1179), .C1(new_n1181), .C2(new_n1183), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1177), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1088), .B1(new_n1169), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(KEYINPUT62), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1191), .B(new_n1177), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1089), .A2(new_n1104), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n993), .B(new_n1000), .C1(new_n1189), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1168), .A2(new_n1142), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1111), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1196), .A2(new_n1188), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1088), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1194), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1000), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT126), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n992), .B1(new_n1195), .B2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g778(.A(G319), .ZN(new_n1205));
  NOR3_X1   g779(.A1(G229), .A2(new_n1205), .A3(G227), .ZN(new_n1206));
  AND3_X1   g780(.A1(new_n862), .A2(new_n657), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n935), .A2(new_n940), .ZN(new_n1208));
  AND2_X1   g782(.A1(new_n1207), .A2(new_n1208), .ZN(G308));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(G225));
endmodule


