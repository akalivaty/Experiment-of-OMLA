//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941;
  NOR2_X1   g000(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT79), .B(KEYINPUT22), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT71), .A2(G125), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT71), .A2(G125), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n197));
  INV_X1    g011(.A(G140), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT71), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT71), .A2(G125), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(G140), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n198), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n200), .B1(new_n207), .B2(KEYINPUT16), .ZN(new_n208));
  AOI211_X1 g022(.A(KEYINPUT72), .B(new_n197), .C1(new_n205), .C2(new_n206), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n199), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(G146), .B(new_n199), .C1(new_n208), .C2(new_n209), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(KEYINPUT73), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n206), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(new_n196), .B2(G140), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT72), .B1(new_n216), .B2(new_n197), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n207), .A2(new_n200), .A3(KEYINPUT16), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT73), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G146), .A4(new_n199), .ZN(new_n221));
  INV_X1    g035(.A(G119), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G128), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G119), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT24), .B(G110), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n231), .B2(new_n223), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n228), .B1(G110), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n214), .A2(new_n221), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT74), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n214), .A2(KEYINPUT74), .A3(new_n221), .A4(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT77), .ZN(new_n239));
  NAND2_X1  g053(.A1(G125), .A2(G140), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n206), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT76), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n206), .A2(KEYINPUT76), .A3(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n239), .B1(new_n245), .B2(new_n211), .ZN(new_n246));
  AOI211_X1 g060(.A(KEYINPUT77), .B(G146), .C1(new_n243), .C2(new_n244), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n232), .ZN(new_n249));
  INV_X1    g063(.A(G110), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n249), .A2(new_n250), .B1(new_n226), .B2(new_n227), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT75), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n213), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n219), .A2(KEYINPUT75), .A3(G146), .A4(new_n199), .ZN(new_n254));
  AOI211_X1 g068(.A(new_n248), .B(new_n251), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n193), .B1(new_n238), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT78), .B1(new_n238), .B2(new_n256), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT78), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n259), .B(new_n255), .C1(new_n236), .C2(new_n237), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n257), .B1(new_n261), .B2(new_n193), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n187), .B1(new_n262), .B2(G902), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  INV_X1    g079(.A(new_n187), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n258), .A2(new_n260), .A3(new_n192), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n265), .B(new_n266), .C1(new_n267), .C2(new_n257), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n263), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G217), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(G234), .B2(new_n265), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(G902), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n262), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n278));
  INV_X1    g092(.A(G137), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(G134), .ZN(new_n280));
  INV_X1    g094(.A(G134), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G137), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT65), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n281), .A2(G137), .ZN(new_n284));
  OAI211_X1 g098(.A(G131), .B(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT11), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n281), .B2(G137), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(KEYINPUT11), .A3(G134), .ZN(new_n288));
  INV_X1    g102(.A(G131), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .A4(new_n282), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n292));
  XNOR2_X1  g106(.A(G143), .B(G146), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(G128), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n224), .A2(new_n211), .A3(G143), .ZN(new_n296));
  INV_X1    g110(.A(G143), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(G146), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n285), .A2(new_n290), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n292), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n287), .A2(new_n288), .A3(new_n282), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G131), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n290), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT0), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n293), .B1(new_n307), .B2(new_n224), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT0), .B(G128), .Z(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n293), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(G116), .B(G119), .Z(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT2), .B(G113), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT70), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(KEYINPUT70), .A3(new_n317), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT69), .B1(new_n312), .B2(new_n315), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n316), .B(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n320), .B(new_n321), .C1(new_n323), .C2(new_n317), .ZN(new_n324));
  INV_X1    g138(.A(G237), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n188), .A3(G210), .ZN(new_n326));
  INV_X1    g140(.A(G101), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n328), .B(new_n329), .Z(new_n330));
  INV_X1    g144(.A(KEYINPUT64), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n310), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n308), .B(KEYINPUT64), .C1(new_n293), .C2(new_n309), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n306), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT66), .ZN(new_n335));
  INV_X1    g149(.A(new_n299), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(new_n300), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n291), .A2(KEYINPUT66), .A3(new_n299), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n315), .ZN(new_n340));
  OR3_X1    g154(.A1(new_n312), .A2(new_n317), .A3(new_n315), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n318), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n330), .B1(new_n342), .B2(KEYINPUT29), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n265), .B1(new_n324), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n303), .A2(KEYINPUT30), .A3(new_n311), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n315), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n316), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n330), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G472), .B1(new_n344), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT31), .B1(new_n349), .B2(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n342), .A2(new_n351), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT31), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n348), .A2(new_n316), .A3(new_n357), .A4(new_n330), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT68), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n358), .A2(new_n359), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n355), .B(new_n356), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(G472), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT32), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(KEYINPUT32), .A3(new_n363), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n354), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n277), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n253), .A2(new_n254), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n216), .A2(KEYINPUT19), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n243), .A2(new_n244), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n211), .B(new_n372), .C1(new_n373), .C2(KEYINPUT19), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n325), .A2(new_n188), .A3(G214), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(new_n297), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G131), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n375), .B(G143), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n289), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n371), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n246), .A2(new_n247), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n216), .A2(G146), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(KEYINPUT18), .A2(G131), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n376), .B(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n383), .A2(KEYINPUT90), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G113), .B(G122), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT90), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n381), .B1(new_n253), .B2(new_n254), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n388), .B1(new_n384), .B2(new_n385), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n391), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT91), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n214), .A2(new_n221), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n376), .A2(KEYINPUT17), .A3(G131), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n403), .B(new_n404), .C1(KEYINPUT17), .C2(new_n380), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n394), .A3(new_n390), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n391), .A2(new_n399), .A3(KEYINPUT91), .A4(new_n395), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(G475), .A2(G902), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT92), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n410), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n410), .A2(KEYINPUT20), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n406), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n394), .B1(new_n405), .B2(new_n390), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n265), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G475), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n224), .A2(G143), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n224), .A2(G143), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n281), .ZN(new_n426));
  INV_X1    g240(.A(G116), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n427), .A2(G122), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT93), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(G122), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G107), .ZN(new_n432));
  INV_X1    g246(.A(G107), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n422), .B1(new_n436), .B2(new_n424), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT95), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n424), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n426), .B(new_n435), .C1(new_n440), .C2(new_n281), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n430), .A2(KEYINPUT14), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT96), .Z(new_n443));
  OAI21_X1  g257(.A(new_n429), .B1(KEYINPUT14), .B2(new_n430), .ZN(new_n444));
  OAI21_X1  g258(.A(G107), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n425), .B(new_n281), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n434), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT9), .B(G234), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(new_n270), .A3(G953), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n448), .B(new_n451), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n452), .A2(G902), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT97), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT15), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n454), .A2(KEYINPUT15), .ZN(new_n457));
  OAI21_X1  g271(.A(G478), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n453), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n417), .A2(new_n421), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G469), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n188), .A2(G227), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(G104), .A3(new_n433), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n393), .A2(G107), .B1(KEYINPUT81), .B2(KEYINPUT3), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n393), .A2(G107), .B1(KEYINPUT81), .B2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n327), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(KEYINPUT4), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT82), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n471), .A2(KEYINPUT4), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT82), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n471), .A2(new_n477), .A3(KEYINPUT4), .A4(new_n472), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n474), .A2(new_n476), .A3(new_n310), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT83), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n475), .B1(KEYINPUT82), .B2(new_n473), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n310), .A4(new_n478), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n433), .A2(G104), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n393), .A2(G107), .ZN(new_n486));
  OAI21_X1  g300(.A(G101), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n472), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n336), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT10), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n306), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n484), .A2(new_n305), .A3(new_n290), .A4(new_n491), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n465), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n299), .B1(new_n472), .B2(new_n487), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n306), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n497), .B(KEYINPUT12), .Z(new_n498));
  AND3_X1   g312(.A1(new_n494), .A2(new_n465), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n462), .B(new_n265), .C1(new_n495), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(G469), .A2(G902), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n493), .A2(new_n494), .A3(new_n465), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n494), .A2(new_n498), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n465), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n500), .B(new_n501), .C1(new_n504), .C2(new_n462), .ZN(new_n505));
  OAI21_X1  g319(.A(G221), .B1(new_n450), .B2(G902), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G952), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n508), .A2(KEYINPUT98), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(KEYINPUT98), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n188), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(G234), .A2(G237), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT21), .B(G898), .Z(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(G902), .A3(G953), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G214), .B1(G237), .B2(G902), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT84), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n474), .A2(new_n476), .A3(new_n315), .A4(new_n478), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT5), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n222), .A3(G116), .ZN(new_n522));
  OAI211_X1 g336(.A(G113), .B(new_n522), .C1(new_n313), .C2(new_n521), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n314), .B2(new_n313), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(new_n488), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT85), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(G110), .B(G122), .Z(new_n529));
  NAND3_X1  g343(.A1(new_n520), .A2(KEYINPUT85), .A3(new_n525), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n526), .A2(new_n529), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n528), .A2(KEYINPUT6), .A3(new_n529), .A4(new_n530), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n310), .A2(new_n196), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n336), .B2(new_n196), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n188), .A2(G224), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n524), .B(new_n488), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT86), .B(KEYINPUT8), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n529), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n538), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n546), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n538), .A2(new_n546), .A3(new_n547), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n534), .A2(new_n545), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n265), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT88), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(KEYINPUT88), .A3(new_n265), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n541), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G210), .B1(G237), .B2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n541), .A2(new_n555), .A3(new_n558), .A4(new_n556), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n519), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n507), .A2(new_n517), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n370), .A2(new_n461), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(G101), .ZN(G3));
  INV_X1    g380(.A(new_n362), .ZN(new_n567));
  OAI21_X1  g381(.A(G472), .B1(new_n567), .B2(G902), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n364), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n275), .B1(new_n269), .B2(new_n271), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT33), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT99), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n452), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n573), .A2(KEYINPUT99), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n452), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n575), .A2(G478), .A3(new_n265), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT100), .B(G478), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n453), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n417), .B2(new_n421), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n572), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT34), .B(G104), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT101), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n585), .B(new_n587), .ZN(G6));
  INV_X1    g402(.A(new_n411), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n408), .A2(new_n409), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n413), .A2(new_n415), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n459), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n591), .A2(new_n421), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n570), .A2(new_n571), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G107), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT102), .B(KEYINPUT35), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G9));
  NOR3_X1   g411(.A1(new_n460), .A2(new_n563), .A3(new_n569), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n261), .B1(KEYINPUT36), .B2(new_n193), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n193), .A2(KEYINPUT36), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n258), .B2(new_n260), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n274), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT103), .B1(new_n272), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT103), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n605), .B(new_n602), .C1(new_n269), .C2(new_n271), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n598), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT37), .B(G110), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G12));
  OAI21_X1  g423(.A(new_n514), .B1(G900), .B2(new_n516), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT104), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n591), .A2(new_n421), .A3(new_n592), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n368), .A2(new_n507), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n562), .B(new_n615), .C1(new_n604), .C2(new_n606), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G128), .ZN(G30));
  NAND2_X1  g431(.A1(new_n560), .A2(new_n561), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT38), .Z(new_n619));
  NAND2_X1  g433(.A1(new_n417), .A2(new_n421), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n592), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n619), .A2(new_n621), .A3(new_n519), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n611), .B(KEYINPUT39), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n507), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n625), .B(KEYINPUT40), .Z(new_n626));
  AOI21_X1  g440(.A(new_n602), .B1(new_n269), .B2(new_n271), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n366), .A2(new_n367), .ZN(new_n628));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  AOI21_X1  g443(.A(G902), .B1(new_n323), .B2(new_n351), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n350), .A2(new_n351), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n622), .A2(new_n626), .A3(new_n627), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G143), .ZN(G45));
  AOI21_X1  g450(.A(new_n414), .B1(new_n410), .B2(new_n411), .ZN(new_n637));
  AOI211_X1 g451(.A(KEYINPUT92), .B(new_n589), .C1(new_n408), .C2(new_n409), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n410), .A2(KEYINPUT20), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n421), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n581), .B(new_n612), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n614), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n643), .B(new_n562), .C1(new_n604), .C2(new_n606), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G146), .ZN(G48));
  OR2_X1    g459(.A1(new_n495), .A2(new_n499), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n265), .ZN(new_n647));
  NAND2_X1  g461(.A1(KEYINPUT105), .A2(G469), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n506), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n562), .A2(new_n517), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n652), .A2(new_n277), .A3(new_n369), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n583), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT41), .B(G113), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G15));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n593), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G116), .ZN(G18));
  NOR2_X1   g472(.A1(new_n652), .A2(new_n369), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n659), .B(new_n461), .C1(new_n604), .C2(new_n606), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G119), .ZN(G21));
  INV_X1    g475(.A(new_n621), .ZN(new_n662));
  INV_X1    g476(.A(new_n652), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n272), .B2(new_n276), .ZN(new_n665));
  AOI211_X1 g479(.A(KEYINPUT107), .B(new_n275), .C1(new_n269), .C2(new_n271), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n324), .A2(new_n351), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n668), .B(new_n355), .C1(new_n360), .C2(new_n361), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n363), .B(KEYINPUT106), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n568), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT108), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n665), .A2(new_n666), .A3(new_n675), .A4(new_n672), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n662), .B(new_n663), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G122), .ZN(G24));
  INV_X1    g492(.A(new_n562), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n650), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n627), .A2(new_n672), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n642), .A2(KEYINPUT109), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n583), .B2(new_n612), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n680), .B(new_n681), .C1(new_n682), .C2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G125), .ZN(G27));
  NAND2_X1  g500(.A1(new_n642), .A2(KEYINPUT109), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n583), .A2(new_n683), .A3(new_n612), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n618), .A2(new_n519), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n507), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n667), .A2(new_n689), .A3(new_n368), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n370), .A2(new_n693), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n697), .A3(new_n689), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n289), .ZN(G33));
  INV_X1    g514(.A(new_n613), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT110), .B(G134), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G36));
  NAND3_X1  g518(.A1(new_n417), .A2(new_n421), .A3(new_n581), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT112), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n709), .A3(new_n706), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n708), .B(new_n710), .C1(new_n711), .C2(new_n705), .ZN(new_n712));
  INV_X1    g526(.A(new_n627), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n569), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT44), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n690), .B(KEYINPUT113), .Z(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n504), .B(KEYINPUT45), .ZN(new_n719));
  OAI21_X1  g533(.A(G469), .B1(new_n719), .B2(G902), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n720), .A2(KEYINPUT46), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(KEYINPUT46), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n500), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n506), .A3(new_n624), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G137), .ZN(G39));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n506), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(KEYINPUT114), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(KEYINPUT114), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n730), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n731), .A2(new_n733), .A3(new_n642), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n369), .A3(new_n277), .A4(new_n690), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G140), .ZN(G42));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n620), .A2(new_n459), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n570), .A3(new_n571), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n607), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n607), .A2(new_n739), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n585), .B1(new_n742), .B2(KEYINPUT115), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n677), .A2(new_n565), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n660), .A2(new_n654), .A3(new_n657), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n681), .B1(new_n682), .B2(new_n684), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n368), .A2(new_n591), .A3(new_n421), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n592), .A2(new_n611), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n749), .B(new_n750), .C1(new_n604), .C2(new_n606), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n693), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n695), .A2(new_n753), .A3(new_n698), .A4(new_n702), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n685), .A2(new_n616), .A3(new_n644), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n621), .A2(new_n679), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n692), .A2(new_n611), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n627), .A3(new_n634), .A4(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT52), .A4(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n685), .A2(new_n644), .A3(new_n759), .A4(new_n616), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT116), .B1(new_n761), .B2(new_n762), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n747), .A2(KEYINPUT53), .A3(new_n754), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n737), .B1(new_n607), .B2(new_n739), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n740), .A2(new_n768), .A3(new_n585), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n565), .A3(new_n677), .A4(new_n745), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n761), .B(KEYINPUT52), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n753), .A2(new_n695), .A3(new_n698), .A4(new_n702), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n766), .B(new_n767), .C1(KEYINPUT53), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT118), .ZN(new_n775));
  INV_X1    g589(.A(new_n744), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n761), .B(new_n762), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n754), .A3(new_n745), .A4(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n767), .A4(new_n766), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n650), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n690), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT120), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(KEYINPUT120), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n786), .A2(new_n787), .A3(new_n514), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(new_n712), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n368), .A3(new_n667), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT48), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(KEYINPUT121), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n277), .A2(KEYINPUT107), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n571), .A2(new_n664), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n673), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n675), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n667), .A2(KEYINPUT108), .A3(new_n673), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n514), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n680), .A3(new_n712), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n791), .A2(KEYINPUT121), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n790), .A2(new_n792), .A3(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n793), .A2(new_n512), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n717), .A3(new_n712), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n649), .ZN(new_n807));
  OAI22_X1  g621(.A1(new_n731), .A2(new_n733), .B1(new_n506), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n799), .A2(KEYINPUT119), .A3(new_n717), .A4(new_n712), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n789), .A2(new_n681), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  INV_X1    g627(.A(new_n634), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n788), .A2(new_n571), .A3(new_n814), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n815), .A2(new_n620), .A3(new_n581), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n619), .A2(new_n519), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n799), .A2(new_n784), .A3(new_n712), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n812), .A2(new_n813), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n810), .A3(new_n816), .A4(new_n811), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT51), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n803), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n677), .A2(new_n741), .A3(new_n743), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n754), .A3(new_n565), .A4(new_n745), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n779), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT117), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n778), .A2(new_n779), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n765), .A2(new_n776), .A3(new_n754), .A4(new_n745), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n779), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n829), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT54), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n815), .A2(new_n584), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n783), .A2(new_n824), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n508), .A2(new_n188), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT49), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n519), .B1(new_n649), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n619), .A2(new_n842), .A3(new_n506), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n705), .B1(KEYINPUT49), .B2(new_n807), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n667), .A3(new_n814), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n840), .A2(new_n846), .ZN(G75));
  AOI21_X1  g661(.A(new_n265), .B1(new_n780), .B2(new_n766), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(G210), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n536), .B(new_n540), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT55), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n853), .B2(KEYINPUT56), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(new_n849), .B2(new_n850), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n188), .A2(G952), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G51));
  XOR2_X1   g672(.A(new_n501), .B(KEYINPUT57), .Z(new_n859));
  AND3_X1   g673(.A1(new_n780), .A2(new_n767), .A3(new_n766), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n767), .B1(new_n780), .B2(new_n766), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(KEYINPUT123), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n646), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n848), .A2(G469), .A3(new_n719), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n857), .B1(new_n866), .B2(new_n867), .ZN(G54));
  NAND3_X1  g682(.A1(new_n848), .A2(KEYINPUT58), .A3(G475), .ZN(new_n869));
  INV_X1    g683(.A(new_n408), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n871), .A2(new_n872), .A3(new_n857), .ZN(G60));
  AND2_X1   g687(.A1(new_n575), .A2(new_n577), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n744), .A2(new_n772), .A3(new_n746), .ZN(new_n875));
  AOI211_X1 g689(.A(KEYINPUT117), .B(KEYINPUT53), .C1(new_n875), .C2(new_n765), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n833), .B1(new_n832), .B2(new_n779), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n876), .A2(new_n877), .A3(new_n830), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n775), .B(new_n782), .C1(new_n878), .C2(new_n767), .ZN(new_n879));
  NAND2_X1  g693(.A1(G478), .A2(G902), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT59), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n874), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n874), .A2(new_n881), .ZN(new_n884));
  INV_X1    g698(.A(new_n766), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n875), .B2(new_n777), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT54), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n887), .B2(new_n774), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n883), .B1(new_n888), .B2(new_n857), .ZN(new_n889));
  INV_X1    g703(.A(new_n884), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n860), .B2(new_n861), .ZN(new_n891));
  INV_X1    g705(.A(new_n857), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(KEYINPUT124), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n882), .A2(new_n894), .ZN(G63));
  NAND2_X1  g709(.A1(new_n780), .A2(new_n766), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n599), .A2(new_n601), .ZN(new_n897));
  NAND2_X1  g711(.A1(G217), .A2(G902), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT60), .Z(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n892), .ZN(new_n901));
  INV_X1    g715(.A(new_n262), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n896), .B2(new_n899), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT61), .ZN(G66));
  NAND2_X1  g719(.A1(new_n515), .A2(G224), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(G953), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n747), .B2(G953), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT125), .Z(new_n909));
  INV_X1    g723(.A(G898), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n536), .B1(new_n910), .B2(G953), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n909), .B(new_n911), .ZN(G69));
  AOI21_X1  g726(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n346), .A2(new_n347), .ZN(new_n914));
  MUX2_X1   g728(.A(new_n373), .B(new_n207), .S(KEYINPUT19), .Z(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT127), .B(G900), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n696), .B(new_n624), .C1(new_n583), .C2(new_n738), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n755), .A2(new_n635), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT62), .Z(new_n921));
  NAND4_X1  g735(.A1(new_n726), .A2(new_n735), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n188), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n913), .B1(new_n923), .B2(new_n916), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n667), .A2(new_n368), .A3(new_n757), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n725), .B1(new_n718), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n699), .B1(new_n701), .B2(new_n696), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n926), .A2(new_n735), .A3(new_n927), .A4(new_n755), .ZN(new_n928));
  INV_X1    g742(.A(new_n916), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n188), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n924), .A2(KEYINPUT126), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT126), .B1(new_n924), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n918), .B1(new_n931), .B2(new_n932), .ZN(G72));
  NAND2_X1  g747(.A1(G472), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT63), .Z(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n928), .B2(new_n770), .ZN(new_n936));
  INV_X1    g750(.A(new_n352), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n857), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n835), .A2(new_n352), .A3(new_n632), .A4(new_n935), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n935), .B1(new_n922), .B2(new_n770), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n631), .B2(new_n941), .ZN(G57));
endmodule


