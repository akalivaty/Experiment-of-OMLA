//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383;
  NOR4_X1   g0000(.A1(KEYINPUT64), .A2(G50), .A3(G58), .A4(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(G50), .ZN(new_n204));
  AOI21_X1  g0004(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NOR3_X1   g0005(.A1(new_n201), .A2(new_n205), .A3(G77), .ZN(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n210), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n203), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n225), .B1(new_n229), .B2(new_n231), .C1(KEYINPUT1), .C2(new_n220), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n222), .A2(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G226), .B(G232), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT67), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n204), .A2(G68), .ZN(new_n247));
  INV_X1    g0047(.A(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n246), .B(new_n252), .ZN(G351));
  AOI21_X1  g0053(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(G1698), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g0060(.A(KEYINPUT69), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  OAI211_X1 g0063(.A(G222), .B(new_n263), .C1(new_n256), .C2(new_n257), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n264), .B1(new_n212), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n254), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G274), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT68), .B(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n276), .B1(G226), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n271), .A2(G190), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT79), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G200), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n271), .B2(new_n281), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT9), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G150), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT72), .B1(new_n266), .B2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT72), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(new_n227), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n290), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n297));
  OAI21_X1  g0097(.A(G20), .B1(new_n201), .B2(new_n205), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT74), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT74), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n300), .B(G20), .C1(new_n201), .C2(new_n205), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT73), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n302), .B(new_n290), .C1(new_n294), .C2(new_n295), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n297), .A2(new_n299), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n306), .A2(KEYINPUT70), .A3(new_n226), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT70), .B1(new_n306), .B2(new_n226), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n226), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT70), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n306), .A2(KEYINPUT70), .A3(new_n226), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(KEYINPUT71), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n304), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n272), .A2(G20), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n315), .A2(G50), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n318), .A2(G50), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AND4_X1   g0122(.A1(new_n288), .A2(new_n317), .A3(new_n320), .A4(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n321), .B1(new_n304), .B2(new_n316), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n288), .B1(new_n324), .B2(new_n320), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n287), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT10), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT10), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n287), .B(new_n328), .C1(new_n323), .C2(new_n325), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n248), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n294), .B2(new_n212), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n309), .A2(new_n332), .A3(new_n314), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT11), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n309), .A2(new_n332), .A3(new_n314), .A4(KEYINPUT11), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT80), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(KEYINPUT80), .A3(new_n336), .ZN(new_n340));
  INV_X1    g0140(.A(G13), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(G1), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT78), .A3(G20), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n318), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n307), .A2(new_n308), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n248), .B1(new_n272), .B2(G20), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT12), .B1(new_n346), .B2(G68), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT12), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n342), .A2(new_n352), .A3(G20), .A4(new_n248), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n349), .A2(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n339), .A2(new_n340), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT14), .ZN(new_n356));
  OAI211_X1 g0156(.A(G226), .B(new_n263), .C1(new_n256), .C2(new_n257), .ZN(new_n357));
  OAI211_X1 g0157(.A(G232), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n254), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  INV_X1    g0162(.A(G41), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT68), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT68), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G41), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n366), .A3(new_n275), .ZN(new_n367));
  INV_X1    g0167(.A(new_n273), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n280), .A2(G238), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n361), .A2(new_n362), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n362), .B1(new_n361), .B2(new_n369), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n356), .B(G169), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n361), .A2(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT13), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n361), .A2(new_n362), .A3(new_n369), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(G179), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n375), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n356), .B1(new_n378), .B2(G169), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n355), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n340), .A2(new_n354), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(G200), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n374), .A2(G190), .A3(new_n375), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(new_n339), .A4(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n330), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G179), .ZN(new_n386));
  OAI211_X1 g0186(.A(G232), .B(new_n263), .C1(new_n256), .C2(new_n257), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n269), .A2(new_n389), .A3(G232), .A4(new_n263), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n256), .A2(new_n257), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G107), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n388), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G238), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n260), .B2(new_n261), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n254), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT77), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n276), .B1(G244), .B2(new_n280), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n397), .B1(new_n396), .B2(new_n398), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n386), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT77), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  XOR2_X1   g0206(.A(KEYINPUT15), .B(G87), .Z(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n293), .A3(new_n291), .ZN(new_n408));
  INV_X1    g0208(.A(new_n289), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n408), .B1(new_n227), .B2(new_n212), .C1(new_n409), .C2(new_n295), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n348), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n349), .A2(G77), .A3(new_n319), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n347), .A2(new_n212), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n401), .A2(new_n406), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(G190), .B1(new_n399), .B2(new_n400), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n403), .A2(G200), .A3(new_n405), .ZN(new_n417));
  INV_X1    g0217(.A(new_n414), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT75), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n271), .A2(new_n281), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(G179), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n271), .A2(KEYINPUT75), .A3(new_n386), .A4(new_n281), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n324), .A2(new_n320), .B1(new_n404), .B2(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n415), .A2(new_n419), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n278), .A2(G232), .A3(new_n279), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT82), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT82), .A4(G232), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n276), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT84), .ZN(new_n433));
  OAI211_X1 g0233(.A(G223), .B(new_n263), .C1(new_n256), .C2(new_n257), .ZN(new_n434));
  OAI211_X1 g0234(.A(G226), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G87), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n254), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n432), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n433), .B1(new_n432), .B2(new_n438), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n285), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G190), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n432), .A2(new_n442), .A3(new_n438), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n315), .A2(new_n318), .ZN(new_n445));
  INV_X1    g0245(.A(new_n295), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n319), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n445), .A2(new_n447), .B1(new_n318), .B2(new_n446), .ZN(new_n448));
  INV_X1    g0248(.A(G58), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n248), .ZN(new_n450));
  OAI21_X1  g0250(.A(G20), .B1(new_n450), .B2(new_n203), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n289), .A2(G159), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n267), .A2(new_n227), .A3(new_n268), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT7), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n268), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n248), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(KEYINPUT81), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT81), .ZN(new_n461));
  AOI211_X1 g0261(.A(new_n461), .B(new_n248), .C1(new_n457), .C2(new_n458), .ZN(new_n462));
  OAI211_X1 g0262(.A(KEYINPUT16), .B(new_n454), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n348), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT7), .B1(new_n391), .B2(new_n227), .ZN(new_n465));
  INV_X1    g0265(.A(new_n458), .ZN(new_n466));
  OAI21_X1  g0266(.A(G68), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n454), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT16), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n448), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n444), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT17), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n404), .B1(new_n439), .B2(new_n440), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n432), .A2(new_n386), .A3(new_n438), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT83), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT83), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n432), .A2(new_n438), .A3(new_n478), .A4(new_n386), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT18), .B1(new_n481), .B2(new_n471), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n432), .A2(new_n438), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT84), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n432), .A2(new_n433), .A3(new_n438), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n486), .A2(new_n404), .B1(new_n477), .B2(new_n479), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n463), .A2(new_n470), .ZN(new_n488));
  INV_X1    g0288(.A(new_n448), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT18), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n444), .A2(KEYINPUT17), .A3(new_n471), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n474), .A2(new_n482), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n385), .A2(new_n427), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(G250), .B1(new_n275), .B2(G1), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT87), .B1(new_n254), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n272), .A2(G45), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n278), .A2(new_n498), .A3(G250), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G274), .ZN(new_n501));
  AND2_X1   g0301(.A1(G1), .A2(G13), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(new_n277), .ZN(new_n503));
  INV_X1    g0303(.A(new_n499), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n497), .A2(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n506));
  OAI211_X1 g0306(.A(G238), .B(new_n263), .C1(new_n256), .C2(new_n257), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G116), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n254), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n505), .A2(new_n510), .A3(new_n442), .ZN(new_n511));
  AOI21_X1  g0311(.A(G200), .B1(new_n505), .B2(new_n510), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n272), .A2(G33), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n315), .A2(G87), .A3(new_n318), .A4(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n346), .A2(new_n407), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n291), .A2(new_n293), .A3(G97), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n269), .A2(new_n227), .A3(G68), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n227), .B1(new_n359), .B2(new_n518), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(G87), .B2(new_n208), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n516), .B1(new_n523), .B2(new_n348), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n505), .A2(new_n510), .A3(new_n386), .ZN(new_n526));
  AOI21_X1  g0326(.A(G169), .B1(new_n505), .B2(new_n510), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n315), .A2(new_n318), .A3(new_n407), .A4(new_n514), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n524), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n513), .A2(new_n525), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n533));
  OAI211_X1 g0333(.A(G244), .B(new_n263), .C1(new_n256), .C2(new_n257), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT85), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n213), .B1(new_n267), .B2(new_n268), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT85), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT4), .A4(new_n263), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n535), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n533), .A2(new_n536), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n254), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT5), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(G41), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(new_n499), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n503), .C1(KEYINPUT5), .C2(new_n274), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT86), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n272), .B(G45), .C1(new_n543), .C2(G41), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n364), .A2(new_n366), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(new_n543), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT86), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n551), .A3(new_n503), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n543), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n254), .B1(new_n553), .B2(new_n545), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n547), .A2(new_n552), .B1(new_n554), .B2(G257), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n542), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G200), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n315), .A2(G97), .A3(new_n318), .A4(new_n514), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n318), .A2(G97), .ZN(new_n559));
  OAI21_X1  g0359(.A(G107), .B1(new_n465), .B2(new_n466), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  AND2_X1   g0361(.A1(G97), .A2(G107), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n207), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n214), .A2(KEYINPUT6), .A3(G97), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n565), .A2(G20), .B1(G77), .B2(new_n289), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n559), .B1(new_n567), .B2(new_n348), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n542), .A2(new_n555), .A3(G190), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n557), .A2(new_n558), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n556), .A2(new_n404), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n542), .A2(new_n555), .A3(new_n386), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n558), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G257), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n575));
  OAI211_X1 g0375(.A(G250), .B(new_n263), .C1(new_n256), .C2(new_n257), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G294), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n554), .A2(G264), .B1(new_n578), .B2(new_n254), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n547), .A2(new_n552), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n315), .A2(G107), .A3(new_n318), .A4(new_n514), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n318), .A2(G107), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT90), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(KEYINPUT25), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(KEYINPUT25), .ZN(new_n587));
  MUX2_X1   g0387(.A(new_n584), .B(new_n586), .S(new_n587), .Z(new_n588));
  AND2_X1   g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n227), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT22), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n269), .A2(new_n592), .A3(new_n227), .A4(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n214), .A3(G20), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT89), .ZN(new_n597));
  NAND2_X1  g0397(.A1(KEYINPUT23), .A2(G107), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n596), .A2(KEYINPUT89), .B1(new_n600), .B2(G20), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT24), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n594), .A2(new_n602), .A3(KEYINPUT24), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n348), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n579), .A2(new_n580), .A3(G190), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n582), .A2(new_n589), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n531), .A2(new_n570), .A3(new_n574), .A4(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT91), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n579), .A2(new_n580), .A3(G179), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n404), .B1(new_n579), .B2(new_n580), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n581), .A2(G169), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n579), .A2(new_n580), .A3(G179), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(KEYINPUT91), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n589), .A2(new_n607), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(G303), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n258), .A2(new_n215), .B1(new_n269), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(G257), .B(new_n263), .C1(new_n256), .C2(new_n257), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n254), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n553), .A2(new_n545), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(G270), .A3(new_n278), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n546), .A2(KEYINPUT86), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n551), .B1(new_n550), .B2(new_n503), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n625), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n580), .A2(KEYINPUT88), .A3(new_n625), .A4(new_n627), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G190), .ZN(new_n635));
  AOI21_X1  g0435(.A(G20), .B1(G33), .B2(G283), .ZN(new_n636));
  INV_X1    g0436(.A(G97), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n636), .B1(G33), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(G116), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G20), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n310), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT20), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n638), .A2(new_n310), .A3(KEYINPUT20), .A4(new_n640), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n643), .A2(new_n644), .B1(new_n347), .B2(new_n639), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n464), .A2(new_n346), .A3(G116), .A4(new_n514), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n632), .A2(G200), .A3(new_n633), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n635), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n404), .B1(new_n645), .B2(new_n646), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n632), .A2(new_n633), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT21), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n580), .A2(G179), .A3(new_n625), .A4(new_n627), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n647), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n632), .A2(KEYINPUT21), .A3(new_n633), .A4(new_n651), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n495), .A2(new_n620), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT92), .Z(G372));
  NAND2_X1  g0462(.A1(new_n615), .A2(new_n616), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT93), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n663), .A2(new_n618), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n664), .B1(new_n663), .B2(new_n618), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n610), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n505), .A2(new_n510), .A3(new_n386), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n505), .A2(new_n510), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n404), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n530), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT26), .B1(new_n674), .B2(new_n531), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n524), .B(new_n515), .C1(new_n511), .C2(new_n512), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n574), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n673), .B1(new_n675), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n495), .B1(new_n669), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n426), .ZN(new_n682));
  INV_X1    g0482(.A(new_n384), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n380), .B1(new_n683), .B2(new_n415), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n444), .A2(KEYINPUT17), .A3(new_n471), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT17), .B1(new_n444), .B2(new_n471), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n492), .A2(new_n482), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n682), .B1(new_n690), .B2(new_n330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n681), .A2(new_n691), .ZN(G369));
  NAND2_X1  g0492(.A1(new_n342), .A2(new_n227), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n648), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n659), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n635), .A2(new_n648), .A3(new_n649), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n668), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n703), .B2(new_n700), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n618), .A2(new_n698), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT94), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n614), .A2(new_n617), .A3(new_n618), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(new_n609), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n619), .A2(new_n698), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n659), .A2(new_n699), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n663), .A2(new_n618), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT93), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n663), .A2(new_n618), .A3(new_n664), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n715), .B1(new_n719), .B2(new_n699), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n713), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n223), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n549), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n231), .B2(new_n724), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n285), .B1(new_n542), .B2(new_n555), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n573), .A2(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n556), .A2(new_n404), .B1(new_n568), .B2(new_n558), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n731), .A2(new_n569), .B1(new_n732), .B2(new_n572), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n609), .A2(new_n673), .A3(new_n676), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n733), .B(new_n734), .C1(new_n659), .C2(new_n619), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT96), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n674), .A2(KEYINPUT26), .A3(new_n531), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n678), .B1(new_n574), .B2(new_n677), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n574), .A2(new_n677), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT96), .B1(new_n740), .B2(KEYINPUT26), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n735), .B(new_n673), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n729), .B1(new_n742), .B2(new_n699), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n733), .B(new_n734), .C1(new_n719), .C2(new_n659), .ZN(new_n744));
  INV_X1    g0544(.A(new_n673), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n737), .B2(new_n738), .ZN(new_n746));
  AOI211_X1 g0546(.A(KEYINPUT29), .B(new_n698), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n556), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n579), .A2(new_n510), .A3(new_n505), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n749), .A2(new_n656), .A3(KEYINPUT30), .A4(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT30), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n505), .A2(new_n510), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n542), .A2(new_n753), .A3(new_n555), .A4(new_n579), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n752), .B1(new_n754), .B2(new_n655), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(KEYINPUT95), .ZN(new_n756));
  AOI21_X1  g0556(.A(G179), .B1(new_n579), .B2(new_n580), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT95), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n671), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n556), .A2(new_n756), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n751), .B(new_n755), .C1(new_n634), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n698), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT31), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n733), .A2(new_n734), .A3(new_n708), .A4(new_n699), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n764), .B(new_n765), .C1(new_n703), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G330), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n748), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n728), .B1(new_n770), .B2(G1), .ZN(G364));
  INV_X1    g0571(.A(new_n705), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n341), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n272), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n723), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n704), .ZN(new_n778));
  INV_X1    g0578(.A(new_n776), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n722), .A2(new_n391), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n780), .A2(G355), .B1(new_n639), .B2(new_n722), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n252), .A2(new_n275), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n722), .A2(new_n269), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G45), .B2(new_n231), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n781), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n226), .B1(G20), .B2(new_n404), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n779), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT97), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G179), .A2(G200), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G20), .A3(new_n442), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT100), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT100), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n227), .A2(new_n285), .A3(G179), .A4(G190), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT99), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n799), .A2(G329), .B1(G283), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT101), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n227), .A2(new_n386), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(new_n442), .A3(new_n285), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n227), .A2(new_n442), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(G179), .A3(new_n285), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G311), .A2(new_n806), .B1(new_n809), .B2(G322), .ZN(new_n810));
  INV_X1    g0610(.A(new_n807), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n811), .A2(new_n285), .A3(G179), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n810), .B(new_n391), .C1(new_n621), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n804), .A2(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(G190), .ZN(new_n816));
  INV_X1    g0616(.A(G317), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G294), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n227), .B1(new_n793), .B2(G190), .ZN(new_n822));
  INV_X1    g0622(.A(G326), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n815), .A2(new_n442), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n820), .B1(new_n821), .B2(new_n822), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  OR3_X1    g0626(.A1(new_n803), .A2(new_n814), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n822), .A2(new_n637), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n825), .A2(new_n204), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT32), .ZN(new_n830));
  INV_X1    g0630(.A(G159), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n794), .A2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n816), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n834), .A2(new_n248), .B1(new_n830), .B2(new_n832), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n812), .A2(G87), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n269), .B1(new_n805), .B2(new_n212), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n808), .B(KEYINPUT98), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G58), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n801), .A2(G107), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n833), .A2(new_n838), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n827), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n789), .ZN(new_n845));
  INV_X1    g0645(.A(new_n788), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n792), .B1(new_n844), .B2(new_n845), .C1(new_n704), .C2(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n778), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  NOR2_X1   g0649(.A1(new_n789), .A2(new_n786), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n779), .B1(new_n212), .B2(new_n850), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n391), .B1(new_n821), .B2(new_n808), .C1(new_n813), .C2(new_n214), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n828), .B(new_n852), .C1(G303), .C2(new_n824), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n801), .A2(G87), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n799), .A2(G311), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G283), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n834), .A2(new_n857), .B1(new_n805), .B2(new_n639), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT102), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n269), .B1(new_n813), .B2(new_n204), .ZN(new_n860));
  INV_X1    g0660(.A(new_n822), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n860), .B1(G58), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n801), .A2(G68), .ZN(new_n863));
  INV_X1    g0663(.A(G132), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n798), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G137), .A2(new_n824), .B1(new_n806), .B2(G159), .ZN(new_n866));
  INV_X1    g0666(.A(G150), .ZN(new_n867));
  INV_X1    g0667(.A(G143), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n866), .B1(new_n867), .B2(new_n834), .C1(new_n839), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT34), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n856), .A2(new_n859), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND4_X1   g0673(.A1(new_n406), .A2(new_n401), .A3(new_n414), .A4(new_n699), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n414), .A2(new_n698), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n419), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n876), .B2(new_n415), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n851), .B1(new_n873), .B2(new_n845), .C1(new_n877), .C2(new_n787), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n699), .B1(new_n669), .B2(new_n680), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n415), .ZN(new_n880));
  INV_X1    g0680(.A(new_n874), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n699), .B(new_n877), .C1(new_n669), .C2(new_n680), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(KEYINPUT103), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT103), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n879), .A2(new_n886), .A3(new_n882), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n768), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n779), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n768), .B1(new_n885), .B2(new_n887), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n878), .B1(new_n889), .B2(new_n890), .ZN(G384));
  NOR2_X1   g0691(.A1(new_n773), .A2(new_n272), .ZN(new_n892));
  INV_X1    g0692(.A(G330), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  INV_X1    g0696(.A(new_n696), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n469), .B1(new_n459), .B2(new_n453), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n348), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n467), .A2(new_n461), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n459), .A2(KEYINPUT81), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n453), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n902), .B2(KEYINPUT16), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n897), .B1(new_n903), .B2(new_n448), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT104), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n896), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n487), .A2(new_n490), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(new_n472), .A4(new_n904), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n472), .A3(new_n904), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n471), .A2(new_n696), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n910), .B2(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n904), .B1(new_n689), .B2(new_n687), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n895), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n315), .B1(new_n902), .B2(KEYINPUT16), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n454), .B1(new_n460), .B2(new_n462), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n469), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n448), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n472), .B1(new_n919), .B2(new_n696), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n481), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n907), .A2(new_n472), .A3(new_n896), .A4(new_n904), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n463), .A2(new_n316), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n900), .A2(new_n901), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT16), .B1(new_n926), .B2(new_n454), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n489), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n494), .A2(new_n897), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(new_n929), .A3(KEYINPUT38), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n894), .B1(new_n915), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n355), .A2(new_n698), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n380), .A2(new_n384), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n355), .B(new_n698), .C1(new_n377), .C2(new_n379), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n881), .A3(new_n880), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n620), .A2(new_n660), .A3(new_n699), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT31), .B1(new_n761), .B2(new_n698), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n936), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT105), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n936), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n767), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT105), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n931), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n928), .A2(new_n897), .B1(new_n471), .B2(new_n444), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n928), .A2(new_n487), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n896), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n923), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n928), .A2(new_n897), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n689), .B2(new_n687), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n952), .A2(new_n954), .A3(new_n895), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT38), .B1(new_n924), .B2(new_n929), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n941), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n947), .B1(new_n894), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n495), .A2(new_n767), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT106), .Z(new_n960));
  AOI21_X1  g0760(.A(new_n893), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT39), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n955), .A2(new_n956), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT39), .B1(new_n915), .B2(new_n930), .ZN(new_n965));
  INV_X1    g0765(.A(new_n380), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n699), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n933), .A2(new_n934), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n884), .B2(new_n881), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n895), .B1(new_n952), .B2(new_n954), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n930), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n689), .B2(new_n897), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n495), .B1(new_n743), .B2(new_n747), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(new_n691), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n975), .B(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n892), .B1(new_n962), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n978), .B2(new_n962), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n639), .B(new_n229), .C1(new_n565), .C2(KEYINPUT35), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(KEYINPUT35), .B2(new_n565), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT36), .ZN(new_n983));
  OAI21_X1  g0783(.A(G77), .B1(new_n449), .B2(new_n248), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n247), .B1(new_n231), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n985), .A2(G1), .A3(new_n341), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(new_n983), .A3(new_n986), .ZN(G367));
  NAND2_X1  g0787(.A1(new_n242), .A2(new_n783), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n789), .B(new_n788), .C1(new_n722), .C2(new_n407), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n779), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n525), .A2(new_n699), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n745), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n677), .B2(new_n991), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n822), .A2(new_n248), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G150), .B2(new_n809), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n996), .A2(KEYINPUT113), .B1(new_n868), .B2(new_n825), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(KEYINPUT113), .B2(new_n996), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT114), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT114), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n800), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n813), .A2(new_n449), .B1(new_n212), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(G137), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n269), .B1(new_n794), .B2(new_n1003), .C1(new_n834), .C2(new_n831), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1002), .B(new_n1004), .C1(G50), .C2(new_n806), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n999), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT115), .Z(new_n1007));
  INV_X1    g0807(.A(KEYINPUT46), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n813), .B2(new_n639), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n812), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(new_n821), .C2(new_n834), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT111), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n805), .A2(new_n857), .B1(new_n822), .B2(new_n214), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G311), .B2(new_n824), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n621), .B2(new_n839), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n391), .B1(new_n794), .B2(new_n817), .C1(new_n1001), .C2(new_n637), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT112), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1007), .A2(new_n1018), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1019), .A2(KEYINPUT47), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n789), .B1(new_n1019), .B2(KEYINPUT47), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n990), .B1(new_n846), .B2(new_n993), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n719), .A2(new_n699), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n573), .A2(new_n698), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n733), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n674), .A2(new_n698), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1023), .B(new_n1027), .C1(new_n709), .C2(new_n714), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT110), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT110), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT44), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n720), .B2(new_n1027), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n715), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n1023), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1027), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(KEYINPUT44), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1029), .A2(KEYINPUT45), .A3(new_n1030), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1033), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n712), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n711), .A2(new_n714), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n1036), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(new_n772), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1033), .A2(new_n1040), .A3(new_n713), .A4(new_n1041), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n770), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n770), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n723), .B(KEYINPUT41), .Z(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n775), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n712), .A2(new_n1027), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT109), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OR3_X1    g0855(.A1(new_n1036), .A2(KEYINPUT42), .A3(new_n1038), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n574), .B1(new_n1025), .B2(new_n708), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT107), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1059), .A2(new_n699), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(KEYINPUT42), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1056), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT108), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT108), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1056), .A2(new_n1065), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n993), .B(KEYINPUT43), .Z(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1055), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1072), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1074), .A2(new_n1054), .A3(new_n1069), .A4(new_n1053), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1022), .B1(new_n1052), .B2(new_n1076), .ZN(G387));
  NAND2_X1  g0877(.A1(new_n1046), .A2(new_n770), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1045), .B(new_n705), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n769), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1080), .A3(new_n723), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n725), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1082), .A2(new_n780), .B1(new_n214), .B2(new_n722), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n239), .A2(new_n275), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n295), .A2(G50), .ZN(new_n1085));
  XOR2_X1   g0885(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1086));
  XNOR2_X1  g0886(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n725), .B(new_n275), .C1(new_n248), .C2(new_n212), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n783), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1083), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n779), .B1(new_n1090), .B2(new_n790), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n812), .A2(G77), .B1(new_n809), .B2(G50), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n801), .A2(G97), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(new_n248), .C2(new_n805), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n269), .B1(new_n794), .B2(new_n867), .C1(new_n834), .C2(new_n295), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n861), .A2(new_n407), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n825), .B2(new_n831), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G311), .A2(new_n816), .B1(new_n806), .B2(G303), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n824), .A2(G322), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n839), .C2(new_n817), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT48), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n812), .A2(G294), .B1(G283), .B2(new_n861), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1107), .A2(KEYINPUT49), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n391), .B1(new_n794), .B2(new_n823), .C1(new_n1001), .C2(new_n639), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n1107), .B2(KEYINPUT49), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1098), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1091), .B1(new_n1111), .B2(new_n845), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n711), .B2(new_n788), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1046), .B2(new_n775), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1081), .A2(new_n1114), .ZN(G393));
  NAND2_X1  g0915(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT117), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n774), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1117), .B2(new_n1116), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n783), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n790), .B1(new_n637), .B2(new_n223), .C1(new_n246), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n776), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n269), .B1(new_n795), .B2(G322), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n842), .B(new_n1123), .C1(new_n857), .C2(new_n813), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT118), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n834), .A2(new_n621), .B1(new_n822), .B2(new_n639), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1127), .A2(KEYINPUT119), .B1(new_n821), .B2(new_n805), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(KEYINPUT119), .B2(new_n1127), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G317), .A2(new_n824), .B1(new_n809), .B2(G311), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT52), .Z(new_n1131));
  NAND2_X1  g0931(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1126), .A2(new_n1129), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G150), .A2(new_n824), .B1(new_n809), .B2(G159), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT51), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n391), .B1(new_n806), .B2(new_n446), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n812), .A2(G68), .B1(G143), .B2(new_n795), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n816), .A2(G50), .B1(G77), .B2(new_n861), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n854), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1133), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1122), .B1(new_n1140), .B2(new_n789), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1027), .B2(new_n846), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1116), .A2(new_n1078), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n723), .A3(new_n1048), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1119), .A2(new_n1142), .A3(new_n1144), .ZN(G390));
  NAND2_X1  g0945(.A1(new_n915), .A2(new_n930), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n963), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n971), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n884), .A2(new_n881), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n935), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1147), .A2(new_n1148), .B1(new_n1150), .B2(new_n967), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1146), .A2(new_n967), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT120), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n935), .B(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n742), .A2(new_n699), .A3(new_n880), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n881), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n768), .A2(new_n882), .A3(new_n969), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1151), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n893), .B1(new_n940), .B2(new_n937), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n877), .A3(new_n935), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n967), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n964), .A2(new_n965), .B1(new_n1162), .B2(new_n970), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n915), .B2(new_n930), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1155), .A2(new_n881), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n1154), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1161), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1154), .B1(new_n768), .B2(new_n882), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1165), .A2(new_n1168), .A3(new_n1161), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n969), .B1(new_n768), .B2(new_n882), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1170), .A2(new_n1161), .B1(new_n881), .B2(new_n884), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1160), .A2(new_n495), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n976), .A2(new_n691), .A3(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1159), .A2(new_n1167), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1158), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n935), .B1(new_n1160), .B2(new_n877), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1149), .B1(new_n1158), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1165), .A2(new_n1168), .A3(new_n1161), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1174), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1163), .A2(new_n1166), .A3(new_n1161), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1176), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1175), .A2(new_n723), .A3(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n269), .B(new_n836), .C1(G97), .C2(new_n806), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G107), .A2(new_n816), .B1(new_n824), .B2(G283), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n799), .A2(G294), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1184), .A2(new_n863), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n808), .A2(new_n639), .B1(new_n822), .B2(new_n212), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT121), .Z(new_n1189));
  INV_X1    g0989(.A(G128), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n834), .A2(new_n1003), .B1(new_n825), .B2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n269), .B1(new_n805), .B2(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1001), .A2(new_n204), .B1(new_n808), .B2(new_n864), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(G125), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n798), .ZN(new_n1197));
  OR3_X1    g0997(.A1(new_n813), .A2(KEYINPUT53), .A3(new_n867), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT53), .B1(new_n813), .B2(new_n867), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n831), .C2(new_n822), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n1187), .A2(new_n1189), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n789), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n850), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1202), .B(new_n776), .C1(new_n446), .C2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1205), .B2(new_n786), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1159), .A2(new_n1167), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1206), .B1(new_n1207), .B2(new_n775), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1183), .A2(new_n1208), .ZN(G378));
  OAI221_X1 g1009(.A(new_n973), .B1(new_n689), .B2(new_n897), .C1(new_n1205), .C2(new_n967), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n893), .B1(new_n957), .B2(new_n894), .ZN(new_n1211));
  XOR2_X1   g1011(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n696), .B1(new_n324), .B2(new_n320), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n330), .B2(new_n426), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n682), .C1(new_n327), .C2(new_n329), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1216), .A2(new_n1217), .A3(KEYINPUT123), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT123), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n324), .A2(new_n320), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT9), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n324), .A2(new_n288), .A3(new_n320), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n328), .B1(new_n1223), .B2(new_n287), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n329), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n426), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1214), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n330), .A2(new_n426), .A3(new_n1215), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1219), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1213), .B1(new_n1218), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT123), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1227), .A2(new_n1219), .A3(new_n1228), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1212), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n931), .A2(new_n943), .A3(new_n946), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1211), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1234), .B1(new_n1211), .B2(new_n1235), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1210), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1234), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n945), .B1(new_n930), .B2(new_n971), .ZN(new_n1240));
  OAI21_X1  g1040(.A(G330), .B1(new_n1240), .B2(KEYINPUT40), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1239), .B1(new_n1241), .B2(new_n947), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1211), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n975), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1238), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n775), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1239), .A2(new_n786), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n776), .B1(G50), .B2(new_n1203), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n799), .A2(G283), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n391), .A2(new_n274), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1250), .B(new_n994), .C1(new_n812), .C2(G77), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G97), .A2(new_n816), .B1(new_n824), .B2(G116), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1001), .A2(new_n449), .B1(new_n808), .B2(new_n214), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n407), .B2(new_n806), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT58), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G50), .B1(new_n266), .B2(new_n363), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1255), .A2(new_n1256), .B1(new_n1250), .B2(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n824), .A2(G125), .B1(G150), .B2(new_n861), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT122), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n834), .A2(new_n864), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n808), .A2(new_n1190), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n813), .A2(new_n1192), .B1(new_n805), .B2(new_n1003), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT59), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n266), .B(new_n363), .C1(new_n1001), .C2(new_n831), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G124), .B2(new_n795), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n1258), .B1(new_n1256), .B2(new_n1255), .C1(new_n1266), .C2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1248), .B1(new_n1270), .B2(new_n789), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1247), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1246), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1174), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1182), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1245), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT57), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n724), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1244), .A2(new_n1238), .B1(new_n1182), .B2(new_n1274), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT57), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1273), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(G375));
  OAI22_X1  g1082(.A1(new_n813), .A2(new_n831), .B1(new_n805), .B2(new_n867), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n391), .B(new_n1283), .C1(G58), .C2(new_n800), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n864), .A2(new_n825), .B1(new_n834), .B2(new_n1192), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(G50), .B2(new_n861), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n840), .A2(G137), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n799), .A2(G128), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1284), .A2(new_n1286), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n813), .A2(new_n637), .B1(new_n805), .B2(new_n214), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n269), .B(new_n1290), .C1(G283), .C2(new_n809), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n801), .A2(G77), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1291), .B(new_n1292), .C1(new_n621), .C2(new_n798), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n1096), .B1(new_n834), .B2(new_n639), .C1(new_n821), .C2(new_n825), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1289), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n789), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1296), .B(new_n776), .C1(G68), .C2(new_n1203), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1154), .B2(new_n786), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1172), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1299), .B2(new_n775), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1051), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1300), .B1(new_n1301), .B2(new_n1303), .ZN(G381));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G378), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1183), .A2(new_n1208), .A3(KEYINPUT124), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1281), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1081), .A2(new_n848), .A3(new_n1114), .ZN(new_n1309));
  OR3_X1    g1109(.A1(G381), .A2(G384), .A3(new_n1309), .ZN(new_n1310));
  OR4_X1    g1110(.A1(G387), .A2(new_n1308), .A3(G390), .A4(new_n1310), .ZN(G407));
  OAI211_X1 g1111(.A(G407), .B(G213), .C1(G343), .C2(new_n1308), .ZN(G409));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1245), .A2(new_n775), .B1(new_n1247), .B2(new_n1271), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n723), .B1(new_n1279), .B2(KEYINPUT57), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1245), .A2(new_n1275), .A3(KEYINPUT57), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G378), .B(new_n1314), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1245), .A2(new_n1275), .A3(new_n1051), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1314), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n697), .A2(G213), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT125), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G384), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  OR2_X1    g1126(.A1(G384), .A2(new_n1324), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1300), .A2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1178), .A2(new_n1174), .A3(new_n1179), .A4(KEYINPUT60), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n723), .ZN(new_n1330));
  OAI21_X1  g1130(.A(KEYINPUT60), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1330), .B1(new_n1331), .B2(new_n1302), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1326), .B1(new_n1328), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1328), .A2(new_n1332), .A3(new_n1326), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1313), .B1(new_n1323), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(G2897), .ZN(new_n1338));
  OAI22_X1  g1138(.A1(new_n1334), .A2(new_n1335), .B1(new_n1338), .B2(new_n1322), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1335), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1322), .A2(new_n1338), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1333), .A3(new_n1341), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(KEYINPUT61), .B1(new_n1323), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1309), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n848), .B1(new_n1081), .B2(new_n1114), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1022), .B(new_n1347), .C1(new_n1052), .C2(new_n1076), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT126), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1350), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1050), .B1(new_n1048), .B2(new_n770), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1073), .B(new_n1075), .C1(new_n1352), .C2(new_n775), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1351), .B1(new_n1353), .B2(new_n1022), .ZN(new_n1354));
  INV_X1    g1154(.A(G390), .ZN(new_n1355));
  NOR3_X1   g1155(.A1(new_n1349), .A2(new_n1354), .A3(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1351), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(G387), .A2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(G390), .B1(new_n1358), .B2(new_n1348), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1356), .A2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1322), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1361), .B1(new_n1317), .B2(new_n1320), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1336), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1362), .A2(KEYINPUT63), .A3(new_n1363), .ZN(new_n1364));
  NAND4_X1  g1164(.A1(new_n1337), .A2(new_n1344), .A3(new_n1360), .A4(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT62), .ZN(new_n1366));
  AND3_X1   g1166(.A1(new_n1362), .A2(new_n1366), .A3(new_n1363), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT61), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1369));
  OAI21_X1  g1169(.A(new_n1368), .B1(new_n1362), .B2(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1366), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1371));
  NOR3_X1   g1171(.A1(new_n1367), .A2(new_n1370), .A3(new_n1371), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1365), .B1(new_n1372), .B2(new_n1360), .ZN(G405));
  NAND2_X1  g1173(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1317), .B1(new_n1281), .B2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1375), .A2(KEYINPUT127), .ZN(new_n1376));
  INV_X1    g1176(.A(KEYINPUT127), .ZN(new_n1377));
  OAI211_X1 g1177(.A(new_n1317), .B(new_n1377), .C1(new_n1281), .C2(new_n1374), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1376), .A2(new_n1336), .A3(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1375), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1380), .A2(new_n1377), .A3(new_n1363), .ZN(new_n1381));
  AND3_X1   g1181(.A1(new_n1379), .A2(new_n1360), .A3(new_n1381), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1360), .B1(new_n1379), .B2(new_n1381), .ZN(new_n1383));
  NOR2_X1   g1183(.A1(new_n1382), .A2(new_n1383), .ZN(G402));
endmodule


