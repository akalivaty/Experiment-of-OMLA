//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n213), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n216), .B(new_n221), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  INV_X1    g0051(.A(G45), .ZN(new_n252));
  AOI21_X1  g0052(.A(G1), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G33), .A3(G41), .ZN(new_n257));
  INV_X1    g0057(.A(new_n219), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n219), .B1(KEYINPUT67), .B2(new_n254), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(new_n257), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n253), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G226), .ZN(new_n265));
  INV_X1    g0065(.A(new_n253), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n262), .B1(new_n261), .B2(new_n257), .ZN(new_n269));
  AND4_X1   g0069(.A1(new_n262), .A2(new_n255), .A3(new_n257), .A4(new_n258), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  OR2_X1    g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n275), .A2(G223), .B1(new_n278), .B2(G77), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1698), .B1(new_n273), .B2(new_n274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G222), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n258), .A2(new_n254), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n265), .B(new_n271), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  OR2_X1    g0084(.A1(new_n284), .A2(G179), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(KEYINPUT69), .ZN(new_n287));
  INV_X1    g0087(.A(G58), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n288), .A2(KEYINPUT8), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(KEYINPUT8), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT69), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n211), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n219), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G50), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n300), .B(new_n219), .C1(G1), .C2(new_n211), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n284), .A2(new_n311), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n285), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n275), .A2(G238), .B1(new_n278), .B2(G107), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n280), .A2(G232), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n271), .B1(new_n316), .B2(new_n283), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n264), .A2(G244), .ZN(new_n318));
  OAI21_X1  g0118(.A(G200), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n301), .ZN(new_n320));
  XOR2_X1   g0120(.A(KEYINPUT8), .B(G58), .Z(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n297), .B1(G20), .B2(G77), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT15), .B(G87), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n295), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n320), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G77), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n304), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n327), .B2(new_n307), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n317), .A2(new_n318), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n319), .B(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n311), .B1(new_n317), .B2(new_n318), .ZN(new_n334));
  INV_X1    g0134(.A(new_n330), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n334), .B(new_n335), .C1(new_n331), .C2(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT9), .B1(new_n302), .B2(new_n309), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n284), .A2(new_n332), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n284), .A2(G200), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n302), .A2(KEYINPUT9), .A3(new_n309), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n339), .A2(new_n340), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT10), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n302), .A2(KEYINPUT9), .A3(new_n309), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n338), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n340), .A4(new_n341), .ZN(new_n348));
  AOI211_X1 g0148(.A(new_n313), .B(new_n337), .C1(new_n344), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G97), .ZN(new_n350));
  INV_X1    g0150(.A(G226), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n272), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n235), .A2(G1698), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n350), .B1(new_n354), .B2(new_n278), .ZN(new_n355));
  INV_X1    g0155(.A(new_n283), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n271), .A2(new_n357), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n224), .B(new_n253), .C1(new_n260), .C2(new_n263), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT13), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(G238), .B(new_n266), .C1(new_n269), .C2(new_n270), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n361), .A2(new_n271), .A3(new_n362), .A4(new_n357), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(G179), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT70), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n360), .A2(new_n366), .A3(new_n363), .ZN(new_n367));
  INV_X1    g0167(.A(new_n358), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n368), .A2(KEYINPUT70), .A3(new_n362), .A4(new_n361), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(G169), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n367), .A2(KEYINPUT14), .A3(G169), .A4(new_n369), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n365), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n294), .A2(new_n327), .B1(new_n211), .B2(G68), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n305), .A2(G20), .A3(G33), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n301), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT11), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT12), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n304), .A2(new_n380), .A3(new_n381), .A4(new_n223), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n223), .B1(new_n380), .B2(new_n381), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n383), .A2(new_n303), .B1(KEYINPUT71), .B2(KEYINPUT12), .ZN(new_n384));
  INV_X1    g0184(.A(new_n307), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n382), .A2(new_n384), .B1(new_n385), .B2(G68), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n375), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n367), .A2(G200), .A3(new_n369), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n363), .A2(G190), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n390), .B2(new_n360), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT72), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT72), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n349), .A2(new_n388), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n351), .A2(G1698), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(G223), .B2(G1698), .ZN(new_n399));
  INV_X1    g0199(.A(G33), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n399), .A2(new_n278), .B1(new_n400), .B2(new_n225), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n356), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n271), .A2(new_n402), .ZN(new_n403));
  AOI211_X1 g0203(.A(new_n235), .B(new_n253), .C1(new_n260), .C2(new_n263), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT74), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n260), .A2(new_n263), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n268), .B1(new_n401), .B2(new_n356), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n264), .A2(G232), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n311), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n303), .B1(new_n287), .B2(new_n292), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n321), .A2(new_n291), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n286), .A2(KEYINPUT69), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n307), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n415), .A3(KEYINPUT73), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT73), .B1(new_n412), .B2(new_n415), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT7), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n273), .A2(new_n274), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(G20), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n223), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n288), .A2(new_n223), .ZN(new_n426));
  OAI21_X1  g0226(.A(G20), .B1(new_n426), .B2(new_n202), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n297), .A2(G159), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n420), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n422), .A2(new_n421), .A3(G20), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT7), .B1(new_n278), .B2(new_n211), .ZN(new_n432));
  OAI21_X1  g0232(.A(G68), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n429), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(KEYINPUT16), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n430), .A2(new_n435), .A3(new_n301), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n419), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n408), .A2(new_n409), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G179), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n411), .A2(KEYINPUT18), .A3(new_n437), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT75), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n411), .A2(new_n437), .A3(new_n441), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n443), .A3(new_n446), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT73), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n287), .A2(new_n292), .A3(new_n385), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n304), .B1(new_n413), .B2(new_n414), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n416), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n433), .A2(new_n434), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n320), .B1(new_n456), .B2(new_n420), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n435), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT74), .B1(new_n403), .B2(new_n404), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n408), .A2(new_n409), .A3(new_n406), .ZN(new_n460));
  AOI21_X1  g0260(.A(G200), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n438), .A2(G190), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT17), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n458), .B(KEYINPUT17), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n450), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n397), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n252), .A2(G1), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n260), .B2(new_n263), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G270), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT79), .A2(G303), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT79), .A2(G303), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n273), .B(new_n274), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(G264), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n481));
  OAI211_X1 g0281(.A(G257), .B(new_n272), .C1(new_n276), .C2(new_n277), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n356), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT76), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n471), .B(G274), .C1(new_n473), .C2(new_n472), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n407), .B2(new_n487), .ZN(new_n488));
  AOI211_X1 g0288(.A(KEYINPUT76), .B(new_n486), .C1(new_n260), .C2(new_n263), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n477), .B(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G200), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n269), .B2(new_n270), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT76), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n407), .A2(new_n485), .A3(new_n487), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n495), .A2(G190), .A3(new_n477), .A4(new_n484), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n303), .A2(G116), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n210), .A2(G33), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n303), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(new_n301), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n500), .B2(G116), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT80), .ZN(new_n502));
  INV_X1    g0302(.A(G116), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n300), .A2(new_n219), .B1(G20), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  INV_X1    g0305(.A(G97), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(new_n211), .C1(G33), .C2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT20), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n504), .A2(KEYINPUT20), .A3(new_n507), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n501), .B(new_n502), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n508), .ZN(new_n511));
  INV_X1    g0311(.A(new_n497), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n320), .A2(new_n303), .A3(new_n498), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n503), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT80), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n491), .A2(new_n496), .A3(new_n510), .A4(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n493), .A2(new_n494), .B1(G270), .B2(new_n476), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n510), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(G179), .A4(new_n484), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n311), .B1(new_n515), .B2(new_n510), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n520), .A2(new_n521), .A3(new_n490), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n520), .B2(new_n490), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n516), .B(new_n519), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT25), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n303), .B2(G107), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n303), .A2(new_n526), .A3(G107), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n527), .A2(new_n529), .B1(new_n500), .B2(G107), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT81), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n211), .B2(G107), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT23), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n532), .B(new_n535), .C1(new_n211), .C2(G107), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n534), .A2(new_n536), .B1(G116), .B2(new_n295), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  AOI21_X1  g0338(.A(G20), .B1(new_n273), .B2(new_n274), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(G87), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n211), .B(G87), .C1(new_n276), .C2(new_n277), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(KEYINPUT22), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n537), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT24), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n541), .A2(KEYINPUT22), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n422), .A2(new_n538), .A3(new_n211), .A4(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n548), .A3(new_n537), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n531), .B1(new_n550), .B2(new_n301), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n488), .A2(new_n489), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n476), .A2(G264), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n280), .A2(G250), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n422), .A2(G257), .A3(G1698), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G294), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n356), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(G200), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n476), .A2(G264), .B1(new_n557), .B2(new_n356), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n495), .A2(G190), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n551), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT83), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n552), .A2(new_n559), .A3(new_n440), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n311), .B1(new_n495), .B2(new_n561), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n495), .A2(new_n561), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G169), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n495), .A2(G179), .A3(new_n561), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(KEYINPUT83), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT82), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n320), .B1(new_n544), .B2(new_n549), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n531), .ZN(new_n576));
  INV_X1    g0376(.A(new_n549), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n548), .B1(new_n547), .B2(new_n537), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n301), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(KEYINPUT82), .A3(new_n530), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n564), .B1(new_n573), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n476), .A2(G257), .ZN(new_n584));
  OAI211_X1 g0384(.A(G250), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n585));
  OAI211_X1 g0385(.A(G244), .B(new_n272), .C1(new_n276), .C2(new_n277), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n505), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT4), .B1(new_n280), .B2(G244), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n356), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n311), .B1(new_n552), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n304), .A2(new_n506), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n513), .B2(new_n506), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT6), .ZN(new_n595));
  INV_X1    g0395(.A(G107), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n506), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n597), .B2(new_n205), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(KEYINPUT6), .A3(G97), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(G20), .B1(G77), .B2(new_n297), .ZN(new_n601));
  OAI21_X1  g0401(.A(G107), .B1(new_n431), .B2(new_n432), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n594), .B1(new_n603), .B2(new_n301), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n586), .A2(new_n587), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n422), .A2(KEYINPUT4), .A3(G244), .A4(new_n272), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n505), .A4(new_n585), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n356), .A2(new_n608), .B1(new_n476), .B2(G257), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n495), .A2(new_n609), .A3(new_n440), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n592), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(G200), .B1(new_n552), .B2(new_n591), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n495), .A2(new_n609), .A3(G190), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n604), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT78), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT19), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n211), .B1(new_n350), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(G87), .B2(new_n206), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n211), .B(G68), .C1(new_n276), .C2(new_n277), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n294), .B2(new_n506), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n301), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n324), .A2(new_n303), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n622), .B(new_n624), .C1(new_n225), .C2(new_n513), .ZN(new_n625));
  INV_X1    g0425(.A(G200), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n210), .A2(G45), .ZN(new_n627));
  NAND2_X1  g0427(.A1(KEYINPUT77), .A2(G250), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n226), .A2(KEYINPUT77), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n210), .A2(new_n267), .A3(G45), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n269), .B2(new_n270), .ZN(new_n634));
  OAI211_X1 g0434(.A(G238), .B(new_n272), .C1(new_n276), .C2(new_n277), .ZN(new_n635));
  OAI211_X1 g0435(.A(G244), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n635), .B(new_n636), .C1(new_n400), .C2(new_n503), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n356), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n626), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n615), .B1(new_n625), .B2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n275), .A2(G244), .B1(G33), .B2(G116), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n283), .B1(new_n641), .B2(new_n635), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n632), .B1(new_n260), .B2(new_n263), .ZN(new_n643));
  OAI21_X1  g0443(.A(G200), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n499), .A2(new_n225), .A3(new_n301), .ZN(new_n645));
  AOI211_X1 g0445(.A(new_n645), .B(new_n623), .C1(new_n621), .C2(new_n301), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(KEYINPUT78), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n634), .A2(new_n638), .A3(G190), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n640), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n634), .A2(new_n638), .A3(new_n440), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n500), .A2(new_n324), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n622), .A2(new_n624), .A3(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n407), .A2(new_n633), .B1(new_n637), .B2(new_n356), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n650), .B(new_n652), .C1(G169), .C2(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n611), .A2(new_n614), .A3(new_n649), .A4(new_n654), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n470), .A2(new_n525), .A3(new_n583), .A4(new_n655), .ZN(G372));
  INV_X1    g0456(.A(new_n654), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n495), .A2(new_n609), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n604), .B1(new_n658), .B2(new_n311), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n649), .A2(new_n659), .A3(new_n610), .A4(new_n654), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n657), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n611), .A2(KEYINPUT84), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT84), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n592), .A2(new_n605), .A3(new_n664), .A4(new_n610), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n644), .A2(new_n646), .A3(new_n648), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(new_n654), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n662), .A2(new_n663), .A3(new_n665), .A4(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n551), .B1(new_n570), .B2(new_n571), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n563), .A2(new_n611), .A3(new_n614), .A4(new_n667), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n661), .B(new_n668), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n470), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n313), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n447), .A2(new_n442), .ZN(new_n676));
  INV_X1    g0476(.A(new_n396), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n388), .B1(new_n677), .B2(new_n336), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n678), .B2(new_n468), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n344), .A2(new_n348), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n675), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n674), .A2(new_n682), .ZN(G369));
  NAND3_X1  g0483(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  INV_X1    g0486(.A(G213), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n684), .B2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G343), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n518), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n525), .B2(KEYINPUT86), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT86), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n524), .A2(new_n695), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n694), .A2(new_n696), .B1(new_n669), .B2(new_n693), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT87), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n697), .B(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n583), .B1(new_n581), .B2(new_n691), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n581), .B1(new_n568), .B2(new_n572), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n703), .B2(new_n691), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n669), .A2(new_n691), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n583), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n670), .B2(new_n691), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT88), .ZN(G399));
  INV_X1    g0512(.A(new_n214), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n217), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  INV_X1    g0519(.A(G330), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n440), .B1(new_n483), .B2(new_n356), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n722), .A2(new_n638), .A3(new_n634), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n495), .A3(new_n609), .A4(new_n561), .ZN(new_n724));
  INV_X1    g0524(.A(new_n517), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n552), .A2(new_n591), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n634), .A3(new_n638), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n559), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n727), .A2(KEYINPUT30), .A3(new_n729), .A4(new_n517), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n653), .A2(G179), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n658), .A2(new_n569), .A3(new_n490), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n726), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n733), .B2(new_n692), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n583), .A2(new_n525), .A3(new_n655), .A4(new_n691), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n720), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n563), .A2(new_n611), .A3(new_n614), .A4(new_n667), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n702), .B2(new_n669), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n662), .A2(KEYINPUT26), .A3(new_n665), .A4(new_n667), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n660), .A2(new_n663), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(new_n743), .A3(new_n654), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n744), .A2(KEYINPUT89), .A3(new_n691), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT89), .B1(new_n744), .B2(new_n691), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT29), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n673), .A2(new_n691), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n738), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n719), .B1(new_n751), .B2(G1), .ZN(G364));
  AND2_X1   g0552(.A1(new_n211), .A2(G13), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n210), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n714), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT90), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n219), .B1(G20), .B2(new_n311), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n214), .A2(new_n422), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n208), .A2(new_n763), .B1(G116), .B2(new_n214), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n713), .A2(new_n422), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n252), .B2(new_n218), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n249), .A2(G45), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n211), .A2(G190), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G179), .A2(G200), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n211), .B1(new_n772), .B2(G190), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n771), .A2(new_n223), .B1(new_n773), .B2(new_n506), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n770), .A2(new_n772), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n211), .A2(new_n440), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G190), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n626), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n780), .A2(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n778), .B1(new_n305), .B2(new_n782), .C1(new_n288), .C2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n779), .A2(new_n332), .A3(new_n626), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(KEYINPUT91), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(KEYINPUT91), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n774), .B(new_n785), .C1(G77), .C2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT92), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n626), .B2(G179), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n440), .A2(KEYINPUT92), .A3(G200), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(new_n795), .A3(new_n770), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n211), .A2(new_n332), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n794), .A2(new_n797), .A3(new_n795), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n422), .B1(new_n796), .B2(new_n596), .C1(new_n225), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  INV_X1    g0601(.A(G326), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n784), .A2(new_n801), .B1(new_n782), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n773), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G294), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n796), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n422), .B1(new_n787), .B2(G311), .ZN(new_n808));
  INV_X1    g0608(.A(new_n775), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G329), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT33), .B(G317), .Z(new_n811));
  OAI211_X1 g0611(.A(new_n808), .B(new_n810), .C1(new_n771), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n798), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n807), .B(new_n812), .C1(G303), .C2(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n792), .A2(new_n800), .B1(new_n805), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n760), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n756), .B1(new_n762), .B2(new_n769), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n697), .B2(new_n759), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n700), .A2(new_n756), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n699), .A2(G330), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  OAI21_X1  g0622(.A(new_n333), .B1(new_n330), .B2(new_n691), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n336), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n336), .A2(new_n692), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n748), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n736), .A2(new_n737), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G330), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n756), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n830), .B2(new_n828), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n827), .A2(new_n758), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n278), .B1(new_n775), .B2(new_n834), .C1(new_n806), .C2(new_n771), .ZN(new_n835));
  INV_X1    g0635(.A(new_n796), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n791), .A2(G116), .B1(G87), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n596), .B2(new_n798), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n835), .B(new_n838), .C1(G303), .C2(new_n781), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n783), .A2(G294), .B1(G97), .B2(new_n804), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT95), .ZN(new_n841));
  INV_X1    g0641(.A(new_n771), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n781), .A2(G137), .B1(new_n842), .B2(G150), .ZN(new_n843));
  INV_X1    g0643(.A(G143), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n844), .B2(new_n784), .C1(new_n790), .C2(new_n776), .ZN(new_n845));
  XOR2_X1   g0645(.A(KEYINPUT96), .B(KEYINPUT34), .Z(new_n846));
  XNOR2_X1  g0646(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n422), .B1(new_n775), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G58), .B2(new_n804), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n836), .A2(G68), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n850), .B(new_n851), .C1(new_n305), .C2(new_n798), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT97), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n839), .A2(new_n841), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n760), .A2(new_n757), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT94), .Z(new_n856));
  OAI22_X1  g0656(.A1(new_n854), .A2(new_n816), .B1(G77), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n756), .B1(new_n833), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n832), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT98), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  OR2_X1    g0661(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n862), .A2(G116), .A3(new_n220), .A4(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT36), .Z(new_n865));
  NOR3_X1   g0665(.A1(new_n426), .A2(new_n217), .A3(new_n327), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n201), .A2(G68), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(KEYINPUT99), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n867), .A2(KEYINPUT99), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n210), .B(G13), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n412), .A2(new_n415), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n436), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n690), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n450), .B2(new_n468), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n459), .A2(new_n460), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n878), .A2(new_n311), .B1(new_n440), .B2(new_n439), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n874), .B1(new_n879), .B2(new_n690), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n877), .B1(new_n880), .B2(new_n463), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n437), .A2(new_n690), .ZN(new_n882));
  AND4_X1   g0682(.A1(new_n877), .A2(new_n463), .A3(new_n445), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n872), .B1(new_n876), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n411), .A2(new_n441), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n886), .A2(new_n689), .B1(new_n436), .B2(new_n873), .ZN(new_n887));
  INV_X1    g0687(.A(new_n463), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n463), .A2(new_n445), .A3(new_n877), .A4(new_n882), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n872), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n467), .B1(new_n448), .B2(new_n449), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n875), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n372), .A2(new_n373), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT72), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT72), .B1(new_n389), .B2(new_n391), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n895), .B(new_n364), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n387), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(new_n691), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(KEYINPUT100), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n900), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n396), .B(new_n902), .C1(new_n899), .C2(new_n374), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT100), .B1(new_n898), .B2(new_n900), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n827), .A2(new_n673), .A3(new_n691), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n825), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n894), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT101), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n676), .A2(new_n689), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n893), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n375), .A2(new_n387), .A3(new_n691), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT38), .B1(new_n881), .B2(new_n883), .ZN(new_n917));
  INV_X1    g0717(.A(new_n875), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n469), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n882), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n676), .B2(new_n467), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n463), .A2(new_n445), .A3(new_n882), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n890), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n914), .B(new_n916), .C1(new_n926), .C2(KEYINPUT39), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n913), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n744), .A2(new_n691), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT89), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n744), .A2(KEYINPUT89), .A3(new_n691), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n749), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n470), .A2(new_n750), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT102), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT102), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n747), .A2(new_n938), .A3(new_n470), .A4(new_n750), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n682), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n930), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n892), .A2(new_n875), .B1(new_n883), .B2(new_n881), .ZN(new_n943));
  INV_X1    g0743(.A(new_n876), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n943), .A2(new_n872), .B1(new_n944), .B2(new_n891), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n826), .B1(new_n736), .B2(new_n737), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n901), .A2(new_n903), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n946), .B1(new_n947), .B2(new_n905), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n942), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT40), .B1(new_n919), .B2(new_n925), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n470), .A2(new_n829), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(G330), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n941), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n210), .B2(new_n753), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n941), .A2(new_n955), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n871), .B1(new_n957), .B2(new_n958), .ZN(G367));
  OAI211_X1 g0759(.A(new_n611), .B(new_n614), .C1(new_n604), .C2(new_n691), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n611), .B2(new_n691), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n709), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n611), .B1(new_n703), .B2(new_n960), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n962), .A2(KEYINPUT42), .B1(new_n691), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(KEYINPUT42), .B2(new_n962), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n691), .A2(new_n646), .ZN(new_n966));
  MUX2_X1   g0766(.A(new_n667), .B(new_n657), .S(new_n966), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT103), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n970), .B(new_n971), .Z(new_n972));
  INV_X1    g0772(.A(new_n705), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n961), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n714), .B(KEYINPUT41), .Z(new_n976));
  AND2_X1   g0776(.A1(new_n710), .A2(new_n961), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT45), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n710), .A2(new_n961), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n973), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n708), .B1(new_n704), .B2(new_n707), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n700), .B(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n978), .A2(new_n705), .A3(new_n980), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n982), .A2(new_n751), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n976), .B1(new_n986), .B2(new_n751), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n975), .B1(new_n987), .B2(new_n755), .ZN(new_n988));
  INV_X1    g0788(.A(new_n756), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n762), .B1(new_n713), .B2(new_n324), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n765), .A2(new_n241), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n759), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n790), .A2(new_n201), .B1(new_n288), .B2(new_n798), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n796), .A2(new_n327), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n278), .B1(new_n842), .B2(G159), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT105), .B(G137), .Z(new_n998));
  OAI221_X1 g0798(.A(new_n997), .B1(new_n775), .B2(new_n998), .C1(new_n782), .C2(new_n844), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n804), .A2(G68), .ZN(new_n1000));
  INV_X1    g0800(.A(G150), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n784), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n999), .B1(KEYINPUT104), .B2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n996), .B(new_n1003), .C1(KEYINPUT104), .C2(new_n1002), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n796), .A2(new_n506), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n422), .B1(new_n809), .B2(G317), .ZN(new_n1006));
  INV_X1    g0806(.A(G294), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n771), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1005), .B(new_n1008), .C1(new_n791), .C2(G283), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n813), .A2(G116), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT46), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n782), .A2(new_n834), .B1(new_n773), .B2(new_n596), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n478), .A2(new_n479), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1012), .B1(new_n1014), .B2(new_n783), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1009), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1004), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT106), .Z(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n992), .B1(new_n993), .B2(new_n967), .C1(new_n1019), .C2(new_n816), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n988), .A2(new_n1020), .ZN(G387));
  OAI22_X1  g0821(.A1(new_n763), .A2(new_n716), .B1(G107), .B2(new_n214), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n238), .A2(new_n252), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n716), .ZN(new_n1024));
  AOI211_X1 g0824(.A(G45), .B(new_n1024), .C1(G68), .C2(G77), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n286), .A2(G50), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT50), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n766), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1022), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n756), .B1(new_n1029), .B2(new_n762), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n782), .A2(new_n801), .B1(new_n771), .B2(new_n834), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G317), .B2(new_n783), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1013), .B2(new_n790), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT48), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n813), .A2(G294), .B1(G283), .B2(new_n804), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT107), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT49), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n278), .B1(new_n775), .B2(new_n802), .C1(new_n796), .C2(new_n503), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT108), .Z(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n804), .A2(new_n324), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n782), .B2(new_n776), .C1(new_n305), .C2(new_n784), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n422), .B1(new_n786), .B2(new_n223), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1005), .B(new_n1047), .C1(G150), .C2(new_n809), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n293), .A2(new_n842), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n813), .A2(G77), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1041), .A2(new_n1044), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1030), .B1(new_n1052), .B2(new_n760), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n704), .B2(new_n993), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT109), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n755), .B2(new_n984), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n984), .A2(new_n751), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT110), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n984), .A2(new_n751), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n714), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1057), .A2(KEYINPUT110), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1056), .B1(new_n1060), .B2(new_n1061), .ZN(G393));
  NAND2_X1  g0862(.A1(new_n986), .A2(new_n714), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT111), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n982), .A2(new_n985), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n981), .A2(KEYINPUT111), .A3(new_n973), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n1059), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT113), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(KEYINPUT113), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1063), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n761), .B1(new_n506), .B2(new_n214), .C1(new_n246), .C2(new_n766), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n989), .B1(new_n1071), .B2(KEYINPUT112), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(KEYINPUT112), .B2(new_n1071), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G311), .A2(new_n783), .B1(new_n781), .B2(G317), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  NAND2_X1  g0875(.A1(new_n804), .A2(G116), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n771), .A2(new_n1013), .B1(new_n775), .B2(new_n801), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n422), .B(new_n1077), .C1(G294), .C2(new_n787), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G283), .A2(new_n813), .B1(new_n836), .B2(G107), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G150), .A2(new_n781), .B1(new_n783), .B2(G159), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT51), .Z(new_n1082));
  OAI221_X1 g0882(.A(new_n422), .B1(new_n775), .B2(new_n844), .C1(new_n201), .C2(new_n771), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G77), .B2(new_n804), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n791), .A2(new_n321), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G68), .A2(new_n813), .B1(new_n836), .B2(G87), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n816), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1073), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n961), .B2(new_n993), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1090), .B1(new_n1092), .B2(new_n754), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1070), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(G390));
  OAI21_X1  g0895(.A(new_n756), .B1(new_n856), .B2(new_n293), .ZN(new_n1096));
  INV_X1    g0896(.A(G125), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n422), .B1(new_n775), .B2(new_n1097), .C1(new_n998), .C2(new_n771), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT54), .B(G143), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n791), .B2(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n784), .A2(new_n848), .B1(new_n773), .B2(new_n776), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G128), .B2(new_n781), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(new_n201), .C2(new_n796), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n813), .A2(G150), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT53), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n783), .A2(G116), .B1(G77), .B2(new_n804), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n806), .B2(new_n782), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n278), .B1(new_n775), .B2(new_n1007), .C1(new_n596), .C2(new_n771), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G87), .B2(new_n813), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1110), .B(new_n851), .C1(new_n506), .C2(new_n790), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1104), .A2(new_n1106), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1096), .B1(new_n1112), .B2(new_n760), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT116), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n914), .B1(new_n926), .B2(KEYINPUT39), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n758), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n933), .A2(new_n934), .A3(new_n825), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1120), .A2(new_n824), .A3(new_n907), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n926), .A2(new_n916), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n908), .A2(new_n825), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n947), .A2(new_n905), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n915), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1116), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n946), .B(G330), .C1(new_n947), .C2(new_n905), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1123), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1119), .B1(new_n1133), .B2(new_n754), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(KEYINPUT117), .B(new_n1119), .C1(new_n1133), .C2(new_n754), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n830), .A2(new_n469), .A3(new_n397), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n682), .B(new_n1138), .C1(new_n937), .C2(new_n939), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT115), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n827), .B1(new_n830), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n738), .A2(KEYINPUT115), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1125), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1120), .A2(new_n824), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n1129), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n829), .A2(G330), .A3(new_n827), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n906), .A3(new_n904), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1129), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT114), .B1(new_n1148), .B2(new_n909), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT114), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1150), .B(new_n1124), .C1(new_n1147), .C2(new_n1129), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1145), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1139), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1133), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1131), .A2(new_n1139), .A3(new_n1152), .A4(new_n1132), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n714), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1136), .A2(new_n1137), .A3(new_n1156), .ZN(G378));
  NAND2_X1  g0957(.A1(new_n680), .A2(new_n675), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n310), .A2(new_n690), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1160), .B(new_n1161), .Z(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n948), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT40), .B1(new_n1164), .B2(new_n894), .ZN(new_n1165));
  OAI21_X1  g0965(.A(G330), .B1(new_n950), .B2(new_n948), .ZN(new_n1166));
  OAI21_X1  g0966(.A(KEYINPUT120), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n447), .A2(new_n442), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n882), .B1(new_n468), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n924), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n872), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n942), .B1(new_n1171), .B2(new_n893), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n720), .B1(new_n1164), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n949), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1163), .B1(new_n1167), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1174), .B1(new_n1173), .B2(new_n949), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(new_n1162), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1176), .A2(new_n1178), .B1(new_n929), .B2(new_n928), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1165), .A2(new_n1166), .A3(KEYINPUT120), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1162), .B1(new_n1180), .B2(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1167), .A2(new_n1163), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n930), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT121), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1179), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n1155), .B2(new_n1139), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1181), .A2(new_n930), .A3(new_n1182), .A4(KEYINPUT121), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1179), .A2(new_n1183), .B1(new_n1155), .B2(new_n1139), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1189), .B(new_n714), .C1(KEYINPUT57), .C2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n989), .B1(new_n201), .B2(new_n855), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n842), .A2(G97), .B1(new_n809), .B2(G283), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n278), .A2(new_n251), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n787), .B2(new_n324), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1195), .A3(new_n1050), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1000), .B1(new_n782), .B2(new_n503), .C1(new_n596), .C2(new_n784), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(G58), .C2(new_n836), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT58), .Z(new_n1199));
  AOI211_X1 g0999(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n776), .B2(new_n796), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT118), .Z(new_n1202));
  INV_X1    g1002(.A(G137), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n786), .A2(new_n1203), .B1(new_n771), .B2(new_n848), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G150), .B2(new_n804), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G125), .A2(new_n781), .B1(new_n783), .B2(G128), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(new_n798), .C2(new_n1099), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1202), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1194), .B(new_n305), .C1(G33), .C2(G41), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1199), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT119), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n760), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1192), .B1(new_n1214), .B2(new_n1216), .C1(new_n1163), .C2(new_n758), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1219), .B2(new_n755), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1191), .A2(new_n1220), .ZN(G375));
  AOI21_X1  g1021(.A(KEYINPUT122), .B1(new_n1152), .B2(new_n755), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n781), .A2(G132), .B1(new_n842), .B2(new_n1100), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n784), .B2(new_n998), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT123), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n278), .B1(new_n809), .B2(G128), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n305), .B2(new_n773), .C1(new_n1001), .C2(new_n786), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n798), .A2(new_n776), .B1(new_n796), .B2(new_n288), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n790), .A2(new_n596), .B1(new_n506), .B2(new_n798), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1045), .B1(new_n782), .B2(new_n1007), .C1(new_n806), .C2(new_n784), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n422), .B1(new_n809), .B2(G303), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n503), .B2(new_n771), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n995), .A4(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n760), .B1(new_n1231), .B2(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1237), .B(new_n756), .C1(G68), .C2(new_n856), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n1125), .B2(new_n757), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1222), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1152), .A2(KEYINPUT122), .A3(new_n755), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1139), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1152), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n976), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n1153), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1243), .A2(new_n1248), .ZN(G381));
  XOR2_X1   g1049(.A(G375), .B(KEYINPUT124), .Z(new_n1250));
  NOR4_X1   g1050(.A1(G387), .A2(G396), .A3(G393), .A4(G384), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1156), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(new_n1134), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(G381), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1094), .A3(new_n1251), .A4(new_n1254), .ZN(G407));
  INV_X1    g1055(.A(new_n1253), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n687), .A2(G343), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1250), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G407), .A2(new_n1258), .A3(G213), .ZN(G409));
  OAI211_X1 g1059(.A(new_n1020), .B(new_n988), .C1(new_n1070), .C2(new_n1093), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT127), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1094), .A2(G387), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(G396), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1261), .A2(new_n1260), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1261), .A2(new_n1263), .B1(new_n1262), .B2(new_n1260), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1139), .A2(new_n1152), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(KEYINPUT60), .B2(new_n1153), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1244), .A2(new_n1245), .A3(KEYINPUT60), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n714), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1243), .B(G384), .C1(new_n1270), .C2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n860), .B1(new_n1274), .B2(new_n1242), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1257), .A2(G2897), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1276), .B(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1218), .B1(new_n1190), .B2(new_n1247), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1185), .A2(new_n755), .A3(new_n1188), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1253), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n714), .B1(new_n1190), .B2(KEYINPUT57), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1185), .A2(new_n1188), .A3(new_n1187), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G378), .B(new_n1220), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT125), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1191), .A2(KEYINPUT125), .A3(G378), .A4(new_n1220), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1281), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1278), .B1(new_n1288), .B2(new_n1257), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1288), .A2(new_n1257), .A3(new_n1276), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1268), .B(new_n1289), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1281), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1257), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1276), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1267), .B1(new_n1292), .B2(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1289), .A2(new_n1268), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1266), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1264), .ZN(new_n1303));
  XOR2_X1   g1103(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1290), .A2(KEYINPUT63), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1301), .A2(new_n1303), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1300), .A2(new_n1307), .ZN(G405));
  NAND2_X1  g1108(.A1(G375), .A2(new_n1256), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1293), .A2(new_n1309), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(new_n1276), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(new_n1303), .ZN(G402));
endmodule


