//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT0), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n197), .B1(KEYINPUT0), .B2(G128), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n192), .A2(new_n193), .A3(new_n196), .A4(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G143), .B(G146), .ZN(new_n200));
  INV_X1    g014(.A(new_n193), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT65), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n199), .A2(new_n202), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n187), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n192), .B2(new_n193), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n198), .A2(new_n193), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n217), .A2(new_n192), .A3(new_n196), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n199), .A2(new_n202), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(KEYINPUT69), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n205), .A2(new_n215), .A3(new_n221), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n212), .A2(G131), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(G143), .B2(new_n188), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n192), .B1(new_n225), .B2(new_n195), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n200), .A2(new_n224), .A3(G128), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n209), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n207), .A2(G137), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n223), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n222), .A2(KEYINPUT30), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT30), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n214), .B1(new_n220), .B2(new_n219), .ZN(new_n235));
  INV_X1    g049(.A(new_n232), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n238));
  INV_X1    g052(.A(G113), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT66), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(KEYINPUT2), .B2(G113), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n240), .A2(new_n242), .B1(KEYINPUT2), .B2(G113), .ZN(new_n243));
  XNOR2_X1  g057(.A(G116), .B(G119), .ZN(new_n244));
  AOI211_X1 g058(.A(KEYINPUT67), .B(KEYINPUT68), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n242), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT2), .A2(G113), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(new_n244), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI22_X1  g065(.A1(new_n245), .A2(new_n251), .B1(new_n243), .B2(new_n244), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n243), .A2(new_n244), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n250), .A3(new_n246), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n233), .A2(new_n237), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n222), .A3(new_n232), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(G210), .ZN(new_n264));
  INV_X1    g078(.A(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n266), .B(new_n267), .Z(new_n268));
  NAND3_X1  g082(.A1(new_n260), .A2(new_n261), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n260), .A2(KEYINPUT31), .A3(new_n261), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n261), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n259), .B1(new_n236), .B2(new_n235), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n258), .A2(new_n222), .A3(KEYINPUT28), .A4(new_n232), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n268), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G472), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n281), .A2(KEYINPUT32), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(G902), .B1(new_n273), .B2(new_n280), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT32), .B1(new_n287), .B2(new_n282), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT32), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(KEYINPUT70), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n222), .A2(new_n232), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT72), .B1(new_n294), .B2(new_n259), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n275), .A3(new_n277), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n258), .A2(new_n222), .A3(KEYINPUT72), .A4(new_n232), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT29), .A3(new_n268), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT73), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n275), .A2(new_n277), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n301), .A2(KEYINPUT71), .A3(new_n268), .A4(new_n276), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n260), .A2(new_n261), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT29), .B1(new_n303), .B2(new_n279), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n305), .B1(new_n278), .B2(new_n279), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n298), .A2(new_n308), .A3(KEYINPUT29), .A4(new_n268), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n300), .A2(new_n283), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n310), .A2(KEYINPUT74), .A3(G472), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT74), .B1(new_n310), .B2(G472), .ZN(new_n312));
  OAI22_X1  g126(.A1(new_n289), .A2(new_n293), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT16), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(G125), .ZN(new_n316));
  XOR2_X1   g130(.A(G125), .B(G140), .Z(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(new_n314), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(G146), .ZN(new_n319));
  INV_X1    g133(.A(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n195), .A2(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT24), .B(G110), .Z(new_n325));
  AOI21_X1  g139(.A(new_n319), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n321), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G110), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(G146), .B(new_n316), .C1(new_n317), .C2(new_n314), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT76), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT75), .B(G110), .ZN(new_n335));
  OAI22_X1  g149(.A1(new_n330), .A2(new_n335), .B1(new_n324), .B2(new_n325), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n334), .B(new_n336), .C1(G146), .C2(new_n317), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(G137), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT77), .B(KEYINPUT22), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n338), .B(new_n342), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n343), .A2(KEYINPUT25), .A3(G902), .ZN(new_n344));
  INV_X1    g158(.A(G217), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(G234), .B2(new_n283), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT25), .B1(new_n343), .B2(G902), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OR3_X1    g162(.A1(new_n343), .A2(G902), .A3(new_n346), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n352));
  INV_X1    g166(.A(G104), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G107), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n353), .A2(G107), .ZN(new_n356));
  OAI21_X1  g170(.A(G101), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(new_n353), .B2(G107), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT3), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G104), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n358), .A2(new_n361), .A3(new_n265), .A4(new_n354), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n225), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n195), .B1(new_n225), .B2(new_n364), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n192), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n363), .B1(new_n368), .B2(new_n227), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n357), .A2(new_n362), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(new_n228), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n215), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT12), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n358), .A2(new_n361), .A3(new_n354), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G101), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n376), .A2(KEYINPUT4), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n376), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(new_n362), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n221), .A4(new_n205), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n205), .A2(new_n221), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT80), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n370), .B(KEYINPUT82), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n226), .B2(new_n227), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n200), .B1(new_n365), .B2(new_n366), .ZN(new_n391));
  INV_X1    g205(.A(new_n227), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n370), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n388), .A2(new_n390), .B1(new_n393), .B2(new_n389), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n384), .A2(new_n387), .A3(new_n394), .A4(new_n214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n374), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n263), .A2(G227), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(G140), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT78), .B(G110), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n384), .A2(new_n387), .A3(new_n394), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n215), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n395), .A3(new_n400), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n352), .B(G469), .C1(new_n407), .C2(G902), .ZN(new_n408));
  INV_X1    g222(.A(G469), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n395), .A2(new_n400), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n395), .A2(KEYINPUT84), .A3(new_n400), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n412), .A2(new_n374), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n400), .B1(new_n404), .B2(new_n395), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n409), .B(new_n283), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n409), .A2(new_n283), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(KEYINPUT83), .B(new_n418), .C1(new_n406), .C2(new_n409), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n408), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G214), .B1(G237), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n219), .A2(G125), .A3(new_n220), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n228), .A2(G125), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n263), .A2(G224), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n423), .A2(new_n424), .B1(KEYINPUT7), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n423), .B(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n428), .A2(KEYINPUT7), .A3(new_n425), .A4(new_n424), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n426), .B1(new_n429), .B2(KEYINPUT86), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n320), .A2(G116), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(KEYINPUT5), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n244), .B2(KEYINPUT5), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n433), .A2(G113), .B1(new_n243), .B2(new_n244), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n388), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g249(.A(G110), .B(G122), .Z(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n435), .B(new_n437), .C1(new_n258), .C2(new_n386), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n434), .A2(new_n363), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n436), .A2(KEYINPUT8), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n363), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(KEYINPUT8), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n439), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n430), .B(new_n444), .C1(KEYINPUT86), .C2(new_n429), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n428), .A2(new_n424), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(G224), .A3(new_n263), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n428), .A2(new_n425), .A3(new_n424), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n435), .B1(new_n258), .B2(new_n386), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n436), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT6), .A3(new_n438), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n453), .A3(new_n436), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n455), .A3(new_n283), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n445), .A2(new_n455), .A3(new_n283), .A4(new_n457), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n422), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT9), .B(G234), .Z(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G221), .B1(new_n463), .B2(G902), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n420), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n463), .A2(new_n345), .A3(G953), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n190), .A2(G128), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n195), .A2(G143), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(new_n207), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT92), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n472));
  INV_X1    g286(.A(G122), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(G116), .ZN(new_n474));
  INV_X1    g288(.A(G116), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT89), .A3(G122), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n474), .A2(new_n476), .B1(G116), .B2(new_n473), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n473), .A2(G116), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n360), .B1(new_n478), .B2(KEYINPUT14), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n477), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n477), .B(new_n360), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n469), .A2(new_n207), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(KEYINPUT91), .ZN(new_n484));
  INV_X1    g298(.A(new_n467), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n486));
  OR3_X1    g300(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT13), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n485), .B2(KEYINPUT13), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n468), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(KEYINPUT13), .B2(new_n485), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n482), .B(new_n484), .C1(new_n490), .C2(new_n207), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n466), .B1(new_n481), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n481), .A2(new_n491), .A3(new_n466), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n283), .ZN(new_n496));
  INV_X1    g310(.A(G478), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n496), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G475), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n262), .A2(new_n263), .A3(G214), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n501), .B(G143), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(new_n213), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT17), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n502), .B(new_n213), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n319), .B(new_n504), .C1(new_n505), .C2(KEYINPUT17), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n317), .B(G146), .ZN(new_n507));
  AND4_X1   g321(.A1(KEYINPUT87), .A2(new_n502), .A3(KEYINPUT18), .A4(G131), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n502), .A2(KEYINPUT87), .B1(KEYINPUT18), .B2(G131), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G113), .B(G122), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n353), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT88), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n506), .A2(new_n510), .A3(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n317), .B(KEYINPUT19), .Z(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n188), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n334), .A2(new_n516), .A3(new_n505), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n512), .B1(new_n517), .B2(new_n510), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n500), .B(new_n283), .C1(new_n514), .C2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT20), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n506), .A2(new_n510), .A3(new_n513), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n517), .A2(new_n510), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n521), .B1(new_n522), .B2(new_n512), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n500), .A4(new_n283), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n512), .B1(new_n506), .B2(new_n510), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n283), .B1(new_n514), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G475), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(G234), .A2(G237), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(G952), .A3(new_n263), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT21), .B(G898), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(G902), .A3(G953), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n499), .A2(new_n530), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n313), .A2(new_n351), .A3(new_n465), .A4(new_n539), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT93), .B(G101), .Z(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(G3));
  INV_X1    g356(.A(new_n538), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n461), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n281), .A2(new_n283), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G472), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n290), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n544), .A2(new_n547), .A3(new_n350), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n420), .A2(new_n464), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT33), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n493), .A2(new_n551), .A3(new_n494), .ZN(new_n552));
  INV_X1    g366(.A(new_n494), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT33), .B1(new_n553), .B2(new_n492), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n554), .A3(G478), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n497), .A2(new_n283), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n495), .A2(new_n497), .A3(new_n283), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n530), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n550), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT34), .B(G104), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(G6));
  XNOR2_X1  g378(.A(new_n526), .B(KEYINPUT94), .ZN(new_n565));
  INV_X1    g379(.A(new_n529), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n499), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n550), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT35), .B(G107), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(G9));
  INV_X1    g385(.A(new_n547), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n342), .A2(KEYINPUT36), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n338), .B(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n574), .B(new_n283), .C1(new_n345), .C2(G234), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n348), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n465), .A2(new_n539), .A3(new_n572), .A4(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT37), .B(G110), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G12));
  INV_X1    g393(.A(G900), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n533), .B1(new_n537), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n568), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n313), .A2(new_n465), .A3(new_n582), .A4(new_n576), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G128), .ZN(G30));
  INV_X1    g398(.A(new_n269), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n297), .A2(new_n279), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n261), .B2(new_n295), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n283), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G472), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n289), .B2(new_n293), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT96), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n290), .A2(new_n291), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(new_n285), .A3(new_n284), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n292), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n589), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n499), .A2(new_n530), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n576), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n459), .A2(new_n460), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(new_n422), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n597), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n597), .A2(KEYINPUT97), .A3(new_n599), .A4(new_n603), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n581), .B(KEYINPUT39), .Z(new_n608));
  NAND2_X1  g422(.A1(new_n549), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(new_n609), .B(KEYINPUT40), .Z(new_n610));
  NAND3_X1  g424(.A1(new_n606), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G143), .ZN(G45));
  NOR3_X1   g426(.A1(new_n561), .A2(KEYINPUT98), .A3(new_n581), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n614));
  INV_X1    g428(.A(new_n530), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n559), .ZN(new_n616));
  INV_X1    g430(.A(new_n581), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n313), .A2(new_n465), .A3(new_n619), .A4(new_n576), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G146), .ZN(G48));
  OAI21_X1  g435(.A(new_n283), .B1(new_n414), .B2(new_n415), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G469), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n623), .A2(new_n464), .A3(new_n416), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n313), .A2(new_n351), .A3(new_n616), .A4(new_n624), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n625), .A2(new_n544), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT41), .B(G113), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G15));
  NAND2_X1  g442(.A1(new_n310), .A2(G472), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT74), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n310), .A2(KEYINPUT74), .A3(G472), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n350), .B1(new_n633), .B2(new_n594), .ZN(new_n634));
  INV_X1    g448(.A(new_n544), .ZN(new_n635));
  INV_X1    g449(.A(new_n568), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n624), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G116), .ZN(G18));
  NAND4_X1  g452(.A1(new_n461), .A2(new_n623), .A3(new_n464), .A4(new_n416), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n313), .A2(new_n539), .A3(new_n576), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G119), .ZN(G21));
  OAI21_X1  g456(.A(new_n273), .B1(new_n268), .B2(new_n298), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n282), .A3(new_n283), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n546), .A2(new_n348), .A3(new_n349), .A4(new_n644), .ZN(new_n645));
  NOR4_X1   g459(.A1(new_n639), .A2(new_n645), .A3(new_n538), .A4(new_n598), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n473), .ZN(G24));
  AND3_X1   g461(.A1(new_n576), .A2(new_n546), .A3(new_n644), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n619), .A2(new_n640), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT99), .B(G125), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G27));
  NAND2_X1  g465(.A1(new_n406), .A2(KEYINPUT100), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n405), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(G469), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n416), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n417), .B1(new_n655), .B2(KEYINPUT101), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n464), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n422), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n459), .A2(new_n460), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT102), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n666));
  AOI211_X1 g480(.A(new_n666), .B(new_n663), .C1(new_n658), .C2(new_n659), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n634), .B(new_n619), .C1(new_n665), .C2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n284), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n592), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n290), .A2(new_n670), .A3(new_n291), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n633), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n674), .A2(KEYINPUT42), .A3(new_n351), .ZN(new_n675));
  INV_X1    g489(.A(new_n619), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n655), .A2(KEYINPUT101), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n418), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT101), .B1(new_n416), .B2(new_n655), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n666), .B1(new_n680), .B2(new_n663), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n660), .A2(KEYINPUT102), .A3(new_n664), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n676), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n668), .A2(new_n669), .B1(new_n675), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n213), .ZN(G33));
  OAI211_X1 g499(.A(new_n634), .B(new_n582), .C1(new_n665), .C2(new_n667), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G134), .ZN(G36));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n559), .A2(new_n530), .A3(KEYINPUT43), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n526), .A2(KEYINPUT105), .A3(new_n529), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT105), .B1(new_n526), .B2(new_n529), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n693), .A3(new_n559), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n547), .B1(new_n696), .B2(KEYINPUT106), .ZN(new_n697));
  INV_X1    g511(.A(new_n693), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n560), .A3(new_n691), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n689), .B1(new_n699), .B2(KEYINPUT43), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n576), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n688), .B1(new_n697), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n576), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n696), .B2(KEYINPUT106), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n572), .B1(new_n700), .B2(new_n701), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT44), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n600), .A2(new_n422), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n703), .A2(new_n707), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n652), .A2(KEYINPUT45), .A3(new_n654), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n711), .B(G469), .C1(KEYINPUT45), .C2(new_n407), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(KEYINPUT46), .A3(new_n418), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n416), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n713), .A2(KEYINPUT104), .A3(new_n416), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n712), .A2(new_n418), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n716), .B(new_n717), .C1(KEYINPUT46), .C2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n710), .A2(new_n719), .A3(new_n464), .A4(new_n608), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n703), .A2(new_n709), .A3(new_n707), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n721), .A2(KEYINPUT107), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n210), .ZN(G39));
  INV_X1    g538(.A(new_n709), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n676), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n719), .A2(new_n464), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n719), .A2(KEYINPUT47), .A3(new_n464), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n727), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n313), .A2(new_n351), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G140), .ZN(G42));
  AND3_X1   g549(.A1(new_n351), .A2(new_n662), .A3(new_n694), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(KEYINPUT108), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n623), .A2(new_n416), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT49), .Z(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n602), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  OR4_X1    g556(.A1(new_n597), .A2(new_n738), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n313), .A2(new_n351), .A3(new_n635), .A4(new_n624), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n646), .B1(new_n744), .B2(new_n636), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n616), .A2(KEYINPUT109), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n616), .A2(KEYINPUT109), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT110), .B1(new_n499), .B2(new_n615), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n499), .A2(new_n615), .A3(KEYINPUT110), .ZN(new_n749));
  OAI22_X1  g563(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n548), .A3(new_n549), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n540), .A2(new_n577), .A3(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n745), .A2(new_n752), .A3(new_n626), .A4(new_n641), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n420), .A2(new_n567), .A3(new_n464), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n600), .A2(new_n422), .A3(new_n499), .A4(new_n581), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n313), .A2(new_n576), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n704), .B1(new_n633), .B2(new_n594), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(KEYINPUT111), .A3(new_n754), .A4(new_n755), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n683), .A2(new_n648), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n686), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n753), .A2(new_n763), .A3(new_n684), .A4(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n464), .B(new_n704), .C1(new_n678), .C2(new_n679), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n461), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n769), .A2(new_n581), .A3(new_n598), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n595), .B1(new_n594), .B2(new_n589), .ZN(new_n771));
  INV_X1    g585(.A(new_n589), .ZN(new_n772));
  AOI211_X1 g586(.A(KEYINPUT96), .B(new_n772), .C1(new_n593), .C2(new_n292), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n768), .B(new_n770), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n583), .A2(new_n620), .A3(new_n649), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n766), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n759), .B(new_n465), .C1(new_n582), .C2(new_n619), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n774), .A3(new_n649), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n783), .B(new_n766), .C1(new_n778), .C2(new_n779), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n778), .B1(new_n783), .B2(new_n779), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n779), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n583), .A2(new_n620), .A3(new_n649), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(KEYINPUT52), .A3(new_n774), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n668), .A2(new_n669), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n675), .A2(new_n683), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n763), .ZN(new_n794));
  INV_X1    g608(.A(new_n646), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n637), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n641), .B1(new_n625), .B2(new_n544), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n540), .A2(new_n577), .A3(new_n751), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n790), .A2(new_n793), .A3(new_n794), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n765), .A2(new_n786), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n800), .A2(new_n802), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n753), .A2(new_n763), .A3(new_n684), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n313), .A2(new_n351), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n681), .B2(new_n682), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n810), .A2(new_n582), .B1(new_n758), .B2(new_n760), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n799), .A2(new_n793), .A3(new_n762), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n808), .A2(new_n786), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n806), .B1(new_n815), .B2(new_n764), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n805), .B1(new_n816), .B2(new_n804), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n739), .A2(new_n661), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n730), .A2(new_n731), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n696), .A2(new_n532), .A3(new_n645), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n709), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n624), .A2(new_n422), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n624), .A2(KEYINPUT116), .A3(new_n422), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n602), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT117), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(new_n828), .A3(new_n602), .A4(new_n825), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n820), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n739), .A2(new_n533), .A3(new_n664), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n833), .A2(new_n700), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n648), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n821), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n821), .A2(new_n837), .A3(new_n832), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n591), .A2(new_n596), .A3(new_n351), .A4(new_n833), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n615), .A3(new_n559), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n836), .A2(KEYINPUT51), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(KEYINPUT51), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n821), .A2(new_n832), .A3(new_n841), .A4(new_n835), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n674), .A2(new_n351), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n834), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT48), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(G952), .A3(new_n263), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n616), .B2(new_n840), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n842), .A2(new_n845), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n820), .A2(new_n640), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n817), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(G952), .A2(G953), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n854), .B(KEYINPUT119), .Z(new_n855));
  OAI21_X1  g669(.A(new_n743), .B1(new_n853), .B2(new_n855), .ZN(G75));
  NOR2_X1   g670(.A1(new_n803), .A2(new_n283), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT56), .B1(new_n857), .B2(G210), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n452), .A2(new_n454), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(new_n449), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT55), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n858), .A2(new_n861), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n263), .A2(G952), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT120), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(G51));
  NOR3_X1   g680(.A1(new_n803), .A2(new_n283), .A3(new_n712), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT121), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n786), .A2(new_n807), .A3(KEYINPUT53), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT52), .B1(new_n788), .B2(new_n774), .ZN(new_n870));
  AND4_X1   g684(.A1(KEYINPUT52), .A2(new_n782), .A3(new_n774), .A4(new_n649), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n802), .B1(new_n812), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n804), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n417), .B(KEYINPUT57), .Z(new_n876));
  OAI22_X1  g690(.A1(new_n875), .A2(new_n876), .B1(new_n415), .B2(new_n414), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n864), .B1(new_n868), .B2(new_n877), .ZN(G54));
  NAND3_X1  g692(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .ZN(new_n879));
  INV_X1    g693(.A(new_n523), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n882), .A3(new_n864), .ZN(G60));
  NAND2_X1  g697(.A1(new_n552), .A2(new_n554), .ZN(new_n884));
  XNOR2_X1  g698(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n556), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n884), .B1(new_n817), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n886), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n875), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n889), .A3(new_n865), .ZN(G63));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n891));
  XNOR2_X1  g705(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n345), .A2(new_n283), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n891), .B1(new_n874), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n894), .ZN(new_n896));
  AOI211_X1 g710(.A(KEYINPUT124), .B(new_n896), .C1(new_n869), .C2(new_n873), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n574), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n865), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT124), .B1(new_n803), .B2(new_n896), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n874), .A2(new_n891), .A3(new_n894), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n343), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n898), .A2(new_n902), .A3(KEYINPUT61), .A4(new_n899), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(G66));
  INV_X1    g721(.A(G224), .ZN(new_n908));
  OAI21_X1  g722(.A(G953), .B1(new_n535), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n799), .B2(G953), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n859), .B1(G898), .B2(new_n263), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(G69));
  NAND2_X1  g726(.A1(new_n233), .A2(new_n237), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n515), .ZN(new_n914));
  INV_X1    g728(.A(new_n723), .ZN(new_n915));
  INV_X1    g729(.A(new_n728), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n769), .A2(new_n598), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n608), .A3(new_n846), .A4(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n734), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n793), .A2(new_n686), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(KEYINPUT125), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n776), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n914), .B1(new_n924), .B2(new_n263), .ZN(new_n925));
  OAI21_X1  g739(.A(G953), .B1(new_n580), .B2(G227), .ZN(new_n926));
  INV_X1    g740(.A(G227), .ZN(new_n927));
  OAI21_X1  g741(.A(G953), .B1(new_n927), .B2(new_n580), .ZN(new_n928));
  INV_X1    g742(.A(new_n914), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n723), .B1(new_n732), .B2(new_n733), .ZN(new_n930));
  INV_X1    g744(.A(new_n611), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT62), .B1(new_n931), .B2(new_n776), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n611), .A2(new_n933), .A3(new_n788), .ZN(new_n934));
  INV_X1    g748(.A(new_n750), .ZN(new_n935));
  OR4_X1    g749(.A1(new_n809), .A2(new_n935), .A3(new_n609), .A4(new_n725), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n930), .A2(new_n932), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n929), .B1(new_n937), .B2(new_n263), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n925), .A2(new_n926), .B1(new_n928), .B2(new_n938), .ZN(G72));
  NAND3_X1  g753(.A1(new_n919), .A2(new_n923), .A3(new_n799), .ZN(new_n940));
  NAND2_X1  g754(.A1(G472), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT63), .Z(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT126), .Z(new_n943));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n303), .A2(new_n268), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n279), .B1(new_n260), .B2(new_n261), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n943), .B1(new_n937), .B2(new_n753), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(KEYINPUT127), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n932), .A2(new_n934), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n951), .A2(new_n799), .A3(new_n930), .A4(new_n936), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n952), .B2(new_n943), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n946), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n942), .ZN(new_n955));
  NOR4_X1   g769(.A1(new_n816), .A2(new_n955), .A3(new_n947), .A4(new_n945), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n954), .A2(new_n864), .A3(new_n956), .ZN(G57));
endmodule


