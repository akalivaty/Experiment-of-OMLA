//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n188), .A2(G128), .A3(new_n190), .A4(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n195), .B1(new_n190), .B2(new_n192), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(G146), .ZN(new_n199));
  AOI21_X1  g013(.A(G128), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n196), .A2(new_n200), .A3(KEYINPUT66), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n199), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n197), .A2(G143), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n202), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n193), .B1(new_n201), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G134), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G131), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n214), .B2(G137), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n215), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n216), .A2(new_n224), .A3(G131), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n211), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n230));
  INV_X1    g044(.A(G113), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT2), .A2(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT69), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G116), .B(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT69), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n236), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n234), .A2(new_n235), .A3(new_n243), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n220), .A2(new_n215), .A3(new_n221), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n223), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n188), .A2(KEYINPUT0), .A3(G128), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  OR2_X1    g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n203), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n228), .A2(new_n248), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(G237), .A2(G953), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G210), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n259), .B(KEYINPUT27), .Z(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n193), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT66), .B1(new_n196), .B2(new_n200), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n205), .A2(new_n209), .A3(new_n202), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT30), .B(new_n256), .C1(new_n269), .C2(new_n226), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n228), .A2(KEYINPUT70), .A3(KEYINPUT30), .A4(new_n256), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n211), .A2(KEYINPUT67), .A3(new_n227), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n269), .B2(new_n226), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n276), .A3(new_n256), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n272), .A2(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT71), .B1(new_n279), .B2(new_n247), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n273), .A2(new_n272), .ZN(new_n282));
  AND4_X1   g096(.A1(KEYINPUT71), .A2(new_n281), .A3(new_n282), .A4(new_n247), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n265), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n282), .A3(new_n247), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT71), .A4(new_n247), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT31), .A3(new_n265), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n257), .B(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n277), .A2(new_n247), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n286), .A2(new_n292), .B1(new_n295), .B2(new_n262), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT32), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n295), .A2(new_n262), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT31), .B1(new_n291), .B2(new_n265), .ZN(new_n301));
  AOI211_X1 g115(.A(new_n285), .B(new_n264), .C1(new_n289), .C2(new_n290), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT32), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n297), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n295), .B2(new_n262), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n257), .B1(new_n280), .B2(new_n283), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(new_n262), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n250), .A2(new_n223), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n255), .A2(new_n252), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n211), .B2(new_n227), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n313), .A2(new_n248), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n262), .A2(new_n306), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n257), .A2(KEYINPUT28), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n313), .B2(new_n248), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n314), .B(new_n315), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G902), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT72), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(KEYINPUT72), .A3(new_n320), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G472), .B1(new_n309), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n316), .A2(new_n318), .ZN(new_n327));
  INV_X1    g141(.A(new_n294), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n329), .B2(new_n263), .ZN(new_n330));
  INV_X1    g144(.A(new_n257), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n289), .B2(new_n290), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n332), .B2(new_n263), .ZN(new_n333));
  INV_X1    g147(.A(new_n323), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(new_n321), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G472), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n299), .A2(new_n305), .B1(new_n326), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G125), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G140), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT16), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n342), .A2(KEYINPUT16), .A3(G140), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G146), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G125), .B(G140), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n197), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n237), .A2(G128), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n237), .A2(G128), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n350), .B(new_n351), .C1(new_n352), .C2(KEYINPUT23), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n353), .A2(G110), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n355));
  INV_X1    g169(.A(new_n352), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(new_n351), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT24), .B(G110), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  OAI22_X1  g173(.A1(new_n354), .A2(new_n355), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n354), .A2(new_n355), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n349), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n353), .A2(G110), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT74), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n344), .A2(new_n345), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n197), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n366), .A2(new_n346), .B1(new_n357), .B2(new_n359), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT22), .B(G137), .ZN(new_n370));
  INV_X1    g184(.A(G953), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n371), .A2(G221), .A3(G234), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n370), .B(new_n372), .Z(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n362), .A2(new_n368), .A3(new_n373), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G902), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT25), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(G234), .B2(new_n320), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n187), .B1(new_n339), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n303), .A2(new_n304), .A3(new_n297), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n304), .B1(new_n303), .B2(new_n297), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n337), .B1(new_n336), .B2(G472), .ZN(new_n389));
  INV_X1    g203(.A(G472), .ZN(new_n390));
  AOI211_X1 g204(.A(KEYINPUT73), .B(new_n390), .C1(new_n333), .C2(new_n335), .ZN(new_n391));
  OAI22_X1  g205(.A1(new_n387), .A2(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n385), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(KEYINPUT76), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n348), .B(new_n197), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n258), .A2(G143), .A3(G214), .ZN(new_n400));
  AOI21_X1  g214(.A(G143), .B1(new_n258), .B2(G214), .ZN(new_n401));
  OAI211_X1 g215(.A(KEYINPUT18), .B(G131), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n258), .A2(G214), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n194), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n258), .A2(G143), .A3(G214), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT18), .A2(G131), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n402), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G131), .B1(new_n400), .B2(new_n401), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(new_n222), .A3(new_n405), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(KEYINPUT17), .B(G131), .C1(new_n400), .C2(new_n401), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n366), .A2(new_n413), .A3(new_n346), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n398), .B(new_n408), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT88), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n341), .A2(new_n343), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT19), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n348), .A2(new_n417), .A3(KEYINPUT19), .ZN(new_n421));
  AOI21_X1  g235(.A(G146), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT89), .B1(new_n422), .B2(new_n347), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT19), .B1(new_n348), .B2(new_n417), .ZN(new_n424));
  AND4_X1   g238(.A1(new_n417), .A2(new_n341), .A3(new_n343), .A4(KEYINPUT19), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n197), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT89), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n346), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n409), .A2(new_n410), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n408), .ZN(new_n431));
  INV_X1    g245(.A(new_n398), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n416), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT20), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT90), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT90), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(KEYINPUT20), .C1(new_n433), .C2(new_n435), .ZN(new_n439));
  OR3_X1    g253(.A1(new_n433), .A2(KEYINPUT20), .A3(new_n435), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT15), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(KEYINPUT92), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(KEYINPUT92), .B2(new_n443), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n194), .A2(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n204), .A2(G143), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(new_n214), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n239), .A2(KEYINPUT14), .A3(G122), .ZN(new_n451));
  XNOR2_X1  g265(.A(G116), .B(G122), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(G107), .B(new_n451), .C1(new_n453), .C2(KEYINPUT14), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n450), .B(new_n454), .C1(G107), .C2(new_n453), .ZN(new_n455));
  INV_X1    g269(.A(G107), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n452), .B(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n449), .A2(new_n214), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT13), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n448), .B1(new_n447), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT91), .ZN(new_n461));
  INV_X1    g275(.A(new_n447), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(KEYINPUT13), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n447), .A2(KEYINPUT91), .A3(new_n459), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n457), .B(new_n458), .C1(new_n465), .C2(new_n214), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT9), .B(G234), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n467), .A2(new_n380), .A3(G953), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n455), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n455), .B2(new_n466), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n320), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n455), .A2(new_n466), .ZN(new_n475));
  INV_X1    g289(.A(new_n468), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(G902), .B1(new_n477), .B2(new_n469), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT93), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n446), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n445), .B1(new_n478), .B2(KEYINPUT93), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n408), .B1(new_n412), .B2(new_n414), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n483), .A2(new_n432), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n320), .B1(new_n484), .B2(new_n416), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G475), .ZN(new_n486));
  NAND2_X1  g300(.A1(G234), .A2(G237), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n487), .A2(G952), .A3(new_n371), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n487), .A2(G902), .A3(G953), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT21), .B(G898), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AND4_X1   g306(.A1(new_n441), .A2(new_n482), .A3(new_n486), .A4(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G214), .B1(G237), .B2(G902), .ZN(new_n494));
  OAI21_X1  g308(.A(G210), .B1(G237), .B2(G902), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT3), .B1(new_n397), .B2(G107), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT3), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n456), .A3(G104), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n397), .A2(G107), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT4), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n501), .A2(new_n502), .A3(G101), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n245), .B2(new_n246), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n501), .B2(G101), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT78), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n507));
  INV_X1    g321(.A(G101), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT77), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT77), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G101), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n506), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n509), .A2(new_n511), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n501), .A2(KEYINPUT78), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n505), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n234), .A2(new_n235), .A3(new_n243), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT69), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT5), .B1(new_n518), .B2(new_n241), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n238), .A2(KEYINPUT5), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(new_n231), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n517), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n456), .A2(G104), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n508), .B1(new_n523), .B2(new_n500), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n499), .A2(new_n500), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n525), .A2(new_n506), .A3(new_n512), .A4(new_n497), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT78), .B1(new_n501), .B2(new_n514), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n504), .A2(new_n516), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G110), .B(G122), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n496), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n530), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n529), .B2(KEYINPUT83), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n504), .A2(new_n516), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n522), .A2(new_n528), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n534), .A2(KEYINPUT83), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n531), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n371), .A2(G224), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT85), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n311), .A2(G125), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT84), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT84), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n311), .A2(new_n543), .A3(G125), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n269), .A2(new_n342), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND4_X1   g361(.A1(new_n540), .A2(new_n546), .A3(new_n542), .A4(new_n544), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n534), .A2(new_n535), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT83), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n529), .A2(KEYINPUT83), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n496), .A4(new_n532), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n537), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT86), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT86), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n537), .A2(new_n554), .A3(new_n549), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n530), .B(KEYINPUT8), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n522), .A2(new_n528), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT87), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n243), .A2(KEYINPUT5), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n517), .B1(new_n521), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n562), .A2(new_n563), .B1(new_n528), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n561), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n545), .B2(new_n546), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n546), .A2(new_n541), .A3(new_n569), .ZN(new_n571));
  OAI22_X1  g385(.A1(new_n570), .A2(new_n571), .B1(new_n550), .B2(new_n532), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n320), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n495), .B1(new_n559), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n495), .ZN(new_n576));
  AOI211_X1 g390(.A(new_n576), .B(new_n573), .C1(new_n556), .C2(new_n558), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n493), .B(new_n494), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G221), .ZN(new_n580));
  INV_X1    g394(.A(new_n467), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n320), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n193), .B(new_n205), .C1(new_n189), .C2(new_n199), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n528), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n503), .A2(new_n311), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n516), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n211), .A2(KEYINPUT10), .A3(new_n528), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n590), .A2(new_n251), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT79), .B1(new_n211), .B2(new_n528), .ZN(new_n592));
  INV_X1    g406(.A(new_n524), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n513), .B2(new_n515), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT79), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n269), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n592), .A2(new_n596), .A3(new_n584), .ZN(new_n597));
  NOR2_X1   g411(.A1(KEYINPUT80), .A2(KEYINPUT12), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n597), .A2(new_n251), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n597), .B2(new_n251), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n591), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(G110), .B(G140), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n371), .A2(G227), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n590), .A2(new_n251), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n590), .A2(new_n251), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n606), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n603), .A2(new_n606), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(G469), .B1(new_n610), .B2(G902), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT81), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT82), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n600), .B2(new_n602), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n597), .A2(new_n251), .A3(new_n599), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n594), .A2(new_n269), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n616), .A2(KEYINPUT79), .B1(new_n528), .B2(new_n583), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n310), .B1(new_n617), .B2(new_n596), .ZN(new_n618));
  OAI211_X1 g432(.A(KEYINPUT82), .B(new_n615), .C1(new_n618), .C2(new_n601), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n614), .A2(new_n609), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n591), .A2(new_n607), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n606), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G469), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n611), .A2(new_n612), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n603), .A2(new_n606), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n609), .A2(new_n607), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n624), .B1(new_n628), .B2(new_n320), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT81), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n582), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n579), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n395), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n514), .ZN(G3));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n393), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n296), .B2(G902), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n636), .B1(new_n298), .B2(new_n296), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n478), .A2(new_n442), .ZN(new_n639));
  NAND2_X1  g453(.A1(G478), .A2(G902), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT33), .B1(new_n470), .B2(new_n471), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n477), .A2(new_n642), .A3(new_n469), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n639), .B(new_n640), .C1(new_n644), .C2(new_n442), .ZN(new_n645));
  AOI211_X1 g459(.A(new_n491), .B(new_n645), .C1(new_n441), .C2(new_n486), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n646), .B(new_n494), .C1(new_n575), .C2(new_n577), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT94), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n559), .A2(new_n574), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n576), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n559), .A2(new_n495), .A3(new_n574), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n653), .A2(KEYINPUT94), .A3(new_n494), .A4(new_n646), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n638), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  XNOR2_X1  g472(.A(new_n491), .B(KEYINPUT96), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n494), .B(new_n659), .C1(new_n575), .C2(new_n577), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n440), .A2(KEYINPUT95), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n440), .A2(KEYINPUT95), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n661), .A2(new_n439), .A3(new_n437), .A4(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n482), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n486), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n638), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT97), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT35), .B(G107), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  AOI21_X1  g484(.A(new_n390), .B1(new_n303), .B2(new_n320), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n296), .A2(new_n298), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n374), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n369), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n383), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n382), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n673), .A2(new_n631), .A3(new_n579), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT37), .B(G110), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT98), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n678), .B(new_n680), .ZN(G12));
  INV_X1    g495(.A(new_n494), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n651), .B2(new_n652), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n489), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n488), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n485), .B2(G475), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n663), .A2(new_n664), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AND4_X1   g506(.A1(new_n392), .A2(new_n692), .A3(new_n631), .A4(new_n677), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n204), .ZN(G30));
  XNOR2_X1  g508(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n653), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n441), .A2(new_n486), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n482), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n696), .A2(new_n682), .A3(new_n677), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n299), .A2(new_n305), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n332), .A2(new_n262), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n331), .A2(new_n263), .ZN(new_n704));
  AOI21_X1  g518(.A(G902), .B1(new_n704), .B2(new_n314), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(G472), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n687), .B(KEYINPUT39), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n631), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n701), .A2(new_n708), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  AOI211_X1 g528(.A(new_n688), .B(new_n645), .C1(new_n441), .C2(new_n486), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n715), .B(new_n494), .C1(new_n575), .C2(new_n577), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT100), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n653), .A2(KEYINPUT100), .A3(new_n494), .A4(new_n715), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n720), .A2(new_n392), .A3(new_n631), .A4(new_n677), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT101), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n326), .A2(new_n338), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n702), .A2(new_n723), .B1(new_n382), .B2(new_n676), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT101), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n631), .A4(new_n720), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G146), .ZN(G48));
  OR2_X1    g542(.A1(new_n623), .A2(new_n624), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n623), .A2(new_n624), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n582), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n655), .A2(new_n392), .A3(new_n393), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  NAND4_X1  g549(.A1(new_n392), .A2(new_n393), .A3(new_n666), .A4(new_n732), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n385), .B1(new_n702), .B2(new_n723), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(KEYINPUT102), .A3(new_n666), .A4(new_n732), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT103), .B(G116), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G18));
  NAND4_X1  g557(.A1(new_n392), .A2(new_n579), .A3(new_n677), .A4(new_n732), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  NAND2_X1  g559(.A1(new_n683), .A2(new_n699), .ZN(new_n746));
  INV_X1    g560(.A(new_n582), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n729), .A2(new_n747), .A3(new_n730), .A4(new_n659), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n263), .B1(new_n293), .B2(new_n314), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n286), .B2(new_n292), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT104), .B1(new_n751), .B2(new_n298), .ZN(new_n752));
  INV_X1    g566(.A(new_n750), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n301), .B2(new_n302), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n297), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n636), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n757), .A3(new_n393), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  INV_X1    g573(.A(new_n715), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n755), .B1(new_n754), .B2(new_n297), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n671), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n677), .A4(new_n756), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n636), .A2(new_n752), .A3(new_n677), .A4(new_n756), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT105), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n760), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n732), .A2(new_n683), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  NOR2_X1   g584(.A1(new_n582), .A2(new_n682), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n651), .A2(new_n652), .A3(new_n771), .ZN(new_n772));
  AOI211_X1 g586(.A(G469), .B(G902), .C1(new_n620), .C2(new_n622), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n629), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT106), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n575), .A2(new_n577), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n730), .A2(new_n611), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT106), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n771), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n392), .A3(new_n393), .A4(new_n715), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n715), .A4(new_n780), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G131), .ZN(G33));
  AND3_X1   g600(.A1(new_n739), .A2(new_n690), .A3(new_n780), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n214), .ZN(G36));
  OAI21_X1  g602(.A(G469), .B1(new_n610), .B2(KEYINPUT45), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(KEYINPUT45), .B2(new_n610), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(G469), .A2(G902), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n730), .B1(new_n794), .B2(KEYINPUT46), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n793), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n747), .B(new_n709), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n645), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n698), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT43), .Z(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n637), .A3(new_n677), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n653), .A2(new_n682), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n797), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(new_n212), .ZN(G39));
  NAND4_X1  g622(.A1(new_n339), .A2(new_n385), .A3(new_n715), .A4(new_n805), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n747), .B1(new_n795), .B2(new_n796), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(KEYINPUT47), .B(new_n747), .C1(new_n795), .C2(new_n796), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n809), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(new_n340), .ZN(G42));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n393), .A2(new_n757), .A3(new_n800), .A4(new_n488), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n682), .A3(new_n696), .A4(new_n732), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT50), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT112), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n805), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT110), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n812), .A2(new_n813), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n731), .A2(new_n747), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT111), .Z(new_n825));
  OAI21_X1  g639(.A(new_n822), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n819), .A2(KEYINPUT112), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n820), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n488), .A2(new_n800), .A3(new_n732), .A4(new_n805), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n764), .A2(new_n766), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT113), .ZN(new_n832));
  INV_X1    g646(.A(new_n708), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n393), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n732), .A2(new_n488), .A3(new_n805), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n698), .A3(new_n645), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n816), .B1(new_n828), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n829), .A2(new_n739), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT48), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n371), .A2(G952), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n817), .B2(new_n768), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n697), .A2(new_n798), .ZN(new_n844));
  INV_X1    g658(.A(new_n836), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n841), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT114), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n838), .A2(new_n819), .A3(new_n816), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n839), .A2(new_n847), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(KEYINPUT115), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(KEYINPUT115), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NOR4_X1   g668(.A1(new_n635), .A2(new_n637), .A3(new_n844), .A4(new_n660), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n395), .B2(new_n632), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n698), .A2(new_n664), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n660), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n673), .A2(new_n858), .A3(new_n393), .A4(new_n631), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n678), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT109), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT109), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n859), .A2(new_n678), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n663), .A2(new_n482), .A3(new_n689), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n653), .A2(new_n682), .A3(new_n865), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n392), .A2(new_n631), .A3(new_n677), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n767), .B2(new_n780), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n856), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n787), .B1(new_n783), .B2(new_n784), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n733), .A2(new_n758), .A3(new_n744), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n741), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT108), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n741), .A3(KEYINPUT108), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n869), .A2(new_n870), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n677), .A2(new_n582), .A3(new_n688), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n683), .A3(new_n699), .A4(new_n777), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n833), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n722), .B2(new_n726), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n693), .B1(new_n767), .B2(new_n768), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n880), .A2(KEYINPUT52), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT52), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n854), .B1(new_n876), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n870), .A2(new_n856), .A3(new_n864), .A4(new_n868), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n887), .A2(new_n854), .A3(new_n872), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n880), .A2(new_n881), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n880), .A2(KEYINPUT52), .A3(new_n881), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n885), .A2(new_n886), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n887), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n871), .A2(new_n741), .A3(KEYINPUT108), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT108), .B1(new_n871), .B2(new_n741), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n893), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n854), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n887), .A2(new_n897), .A3(new_n898), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT53), .B1(new_n902), .B2(new_n893), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n895), .B1(new_n904), .B2(new_n886), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n852), .A2(new_n853), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(G952), .A2(G953), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n731), .B(KEYINPUT49), .Z(new_n908));
  NOR3_X1   g722(.A1(new_n799), .A2(new_n582), .A3(new_n682), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n696), .A3(new_n909), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n906), .A2(new_n907), .B1(new_n834), .B2(new_n910), .ZN(G75));
  NAND2_X1  g725(.A1(new_n885), .A2(new_n894), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(G210), .A3(G902), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n537), .A2(new_n554), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n549), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT55), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(KEYINPUT56), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n371), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT116), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n913), .A2(new_n922), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n916), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(KEYINPUT117), .B(new_n916), .C1(new_n925), .C2(new_n926), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n921), .B1(new_n929), .B2(new_n930), .ZN(G51));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n912), .A2(G902), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n792), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n620), .A2(new_n622), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n793), .B(KEYINPUT57), .Z(new_n937));
  AND3_X1   g751(.A1(new_n871), .A2(new_n741), .A3(KEYINPUT53), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n869), .A2(new_n870), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n884), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n903), .A2(new_n940), .A3(KEYINPUT54), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n886), .B1(new_n885), .B2(new_n894), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT118), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n936), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n937), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT54), .B1(new_n903), .B2(new_n940), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n895), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(KEYINPUT118), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n934), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n932), .B1(new_n950), .B2(new_n919), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n935), .B1(new_n948), .B2(KEYINPUT118), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n943), .A2(new_n944), .ZN(new_n953));
  OAI22_X1  g767(.A1(new_n952), .A2(new_n953), .B1(new_n792), .B2(new_n933), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(KEYINPUT119), .A3(new_n920), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(G54));
  NAND4_X1  g770(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(new_n433), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n433), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n919), .ZN(G60));
  XOR2_X1   g774(.A(new_n640), .B(KEYINPUT59), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n644), .B1(new_n905), .B2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n644), .B(new_n962), .C1(new_n941), .C2(new_n942), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n920), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT120), .ZN(new_n966));
  OR3_X1    g780(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n963), .B2(new_n965), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(G63));
  INV_X1    g783(.A(KEYINPUT122), .ZN(new_n970));
  XNOR2_X1  g784(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n380), .A2(new_n320), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n912), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n973), .ZN(new_n975));
  AOI211_X1 g789(.A(KEYINPUT122), .B(new_n975), .C1(new_n885), .C2(new_n894), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n919), .B1(new_n977), .B2(new_n377), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n900), .A2(new_n854), .B1(new_n893), .B2(new_n888), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT122), .B1(new_n980), .B2(new_n975), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n912), .A2(new_n970), .A3(new_n973), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n675), .B(KEYINPUT123), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n984), .ZN(new_n986));
  AOI211_X1 g800(.A(KEYINPUT124), .B(new_n986), .C1(new_n981), .C2(new_n982), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n978), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT61), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n978), .B(KEYINPUT61), .C1(new_n985), .C2(new_n987), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(G66));
  INV_X1    g806(.A(G224), .ZN(new_n993));
  OAI21_X1  g807(.A(G953), .B1(new_n490), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n856), .A2(new_n864), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n899), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n994), .B1(new_n997), .B2(G953), .ZN(new_n998));
  INV_X1    g812(.A(G898), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n914), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n998), .B(new_n1000), .Z(G69));
  NAND2_X1  g815(.A1(new_n420), .A2(new_n421), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n279), .B(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n797), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n339), .A2(new_n385), .A3(new_n746), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n807), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n809), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n823), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1006), .A2(new_n1008), .A3(new_n870), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n881), .A2(new_n727), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1009), .A2(G953), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n684), .A2(new_n371), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1003), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n857), .A2(new_n844), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n805), .A2(new_n1015), .ZN(new_n1016));
  AOI211_X1 g830(.A(new_n710), .B(new_n1016), .C1(new_n386), .C2(new_n394), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n814), .A2(new_n807), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1010), .A2(new_n713), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(KEYINPUT125), .B1(new_n1022), .B2(new_n371), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT125), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1024), .B1(new_n1022), .B2(new_n371), .ZN(new_n1025));
  OAI22_X1  g839(.A1(new_n1014), .A2(new_n1023), .B1(new_n1025), .B2(new_n1003), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n371), .B1(G227), .B2(G900), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT126), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(KEYINPUT127), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT127), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1026), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1027), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1030), .B(new_n1032), .C1(new_n1026), .C2(new_n1033), .ZN(G72));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1037), .B1(new_n1038), .B2(new_n997), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n291), .A2(new_n704), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n920), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n308), .A2(new_n262), .ZN(new_n1042));
  AOI211_X1 g856(.A(new_n1037), .B(new_n904), .C1(new_n284), .C2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1036), .B1(new_n1022), .B2(new_n996), .ZN(new_n1044));
  AOI211_X1 g858(.A(new_n1041), .B(new_n1043), .C1(new_n703), .C2(new_n1044), .ZN(G57));
endmodule


