//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G231gat), .A2(G233gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G1gat), .B2(new_n205), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G57gat), .B(G64gat), .Z(new_n211));
  AND2_X1   g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(KEYINPUT9), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G71gat), .B(G78gat), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n213), .B(new_n214), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT21), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n210), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n216), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n218), .B2(new_n219), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n204), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n219), .ZN(new_n225));
  INV_X1    g024(.A(new_n220), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n227), .A2(G231gat), .A3(G233gat), .A4(new_n221), .ZN(new_n228));
  XNOR2_X1  g027(.A(G127gat), .B(G155gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(G211gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n224), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n224), .B2(new_n228), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n203), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(new_n228), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n230), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(new_n202), .A3(new_n232), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT100), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n241));
  XNOR2_X1  g040(.A(G134gat), .B(G162gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G85gat), .ZN(new_n245));
  INV_X1    g044(.A(G92gat), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT98), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT98), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(G85gat), .A3(G92gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT7), .ZN(new_n250));
  NAND2_X1  g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251));
  AOI22_X1  g050(.A1(KEYINPUT8), .A2(new_n251), .B1(new_n245), .B2(new_n246), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT7), .ZN(new_n253));
  OAI211_X1 g052(.A(KEYINPUT98), .B(new_n253), .C1(new_n245), .C2(new_n246), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G99gat), .B(G106gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n257), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT99), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT99), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n255), .A2(new_n261), .A3(new_n257), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT93), .ZN(new_n264));
  NOR2_X1   g063(.A1(G29gat), .A2(G36gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(KEYINPUT14), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G29gat), .A2(G36gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT14), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n271), .B(KEYINPUT92), .C1(G29gat), .C2(G36gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G43gat), .B(G50gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(KEYINPUT15), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(KEYINPUT15), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n274), .A2(KEYINPUT15), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n273), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n264), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n280), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(KEYINPUT93), .A3(new_n275), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n263), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G190gat), .B(G218gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(KEYINPUT94), .B(KEYINPUT17), .Z(new_n291));
  NAND3_X1  g090(.A1(new_n283), .A2(new_n281), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n282), .A2(KEYINPUT17), .A3(new_n275), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n292), .A2(new_n293), .A3(new_n262), .A4(new_n260), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n286), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n290), .B1(new_n286), .B2(new_n294), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n244), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n297), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(new_n243), .A3(new_n295), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n239), .A2(new_n240), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n235), .A2(new_n238), .ZN(new_n303));
  INV_X1    g102(.A(new_n301), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT100), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n308));
  NAND2_X1  g107(.A1(G227gat), .A2(G233gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n311));
  INV_X1    g110(.A(G127gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G134gat), .ZN(new_n313));
  INV_X1    g112(.A(G134gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G127gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT69), .B1(new_n312), .B2(G134gat), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT70), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n317), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n320));
  XNOR2_X1  g119(.A(G127gat), .B(G134gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n319), .B(new_n320), .C1(new_n321), .C2(new_n311), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323));
  XOR2_X1   g122(.A(G113gat), .B(G120gat), .Z(new_n324));
  AOI22_X1  g123(.A1(new_n318), .A2(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n326));
  AND2_X1   g125(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n326), .B(G113gat), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G113gat), .ZN(new_n330));
  OR2_X1    g129(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(KEYINPUT71), .A2(G120gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G120gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT72), .B1(new_n334), .B2(G113gat), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n329), .B(new_n321), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT73), .B(KEYINPUT1), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n325), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT67), .ZN(new_n342));
  NAND2_X1  g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT67), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n344), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346));
  INV_X1    g145(.A(G169gat), .ZN(new_n347));
  INV_X1    g146(.A(G176gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n342), .A2(new_n343), .A3(new_n345), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT68), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT27), .B(G183gat), .ZN(new_n356));
  INV_X1    g155(.A(G190gat), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n355), .B(new_n357), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n354), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n350), .A2(new_n364), .A3(new_n351), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT66), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT28), .A3(new_n361), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n353), .A2(new_n363), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n347), .A2(new_n348), .ZN(new_n370));
  AND2_X1   g169(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n371));
  NOR2_X1   g170(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n347), .B(new_n348), .C1(KEYINPUT64), .C2(KEYINPUT23), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n343), .ZN(new_n375));
  OR2_X1    g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT24), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT65), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n378), .A3(new_n351), .ZN(new_n379));
  AND2_X1   g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(KEYINPUT65), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT25), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT25), .B1(new_n385), .B2(KEYINPUT24), .ZN(new_n386));
  INV_X1    g185(.A(new_n343), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT64), .B(KEYINPUT23), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(new_n370), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n380), .A2(new_n377), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n386), .A2(new_n389), .A3(new_n374), .A4(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n340), .A2(new_n369), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n324), .A2(new_n323), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n314), .A2(G127gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n312), .A2(G134gat), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT69), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n320), .B1(new_n397), .B2(new_n319), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n316), .A2(KEYINPUT70), .A3(new_n317), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n333), .A2(new_n335), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n401), .A2(new_n321), .A3(new_n329), .A4(new_n337), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n369), .A2(new_n392), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n310), .B1(new_n393), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT74), .B(KEYINPUT33), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(KEYINPUT32), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G15gat), .B(G43gat), .Z(new_n408));
  XNOR2_X1  g207(.A(G71gat), .B(G99gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n405), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(KEYINPUT32), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT75), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT75), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n404), .A2(new_n414), .A3(KEYINPUT32), .A4(new_n411), .ZN(new_n415));
  AOI221_X4 g214(.A(new_n308), .B1(new_n407), .B2(new_n410), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n308), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n415), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n407), .A2(new_n410), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n369), .A2(new_n392), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n400), .A2(new_n402), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n340), .A2(new_n369), .A3(new_n392), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(new_n310), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n416), .A2(new_n420), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT32), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n425), .B2(new_n310), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n414), .B1(new_n430), .B2(new_n411), .ZN(new_n431));
  INV_X1    g230(.A(new_n415), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n419), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n308), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n417), .A3(new_n419), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n426), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n307), .B1(new_n428), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT36), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G50gat), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(KEYINPUT78), .ZN(new_n442));
  XNOR2_X1  g241(.A(G197gat), .B(G204gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G211gat), .B(G218gat), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n442), .B(new_n443), .C1(KEYINPUT79), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(KEYINPUT79), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT3), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G148gat), .ZN(new_n450));
  INV_X1    g249(.A(G141gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT83), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G141gat), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n450), .A2(G141gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT84), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT83), .B(G141gat), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n459), .B(new_n456), .C1(new_n460), .C2(new_n450), .ZN(new_n461));
  INV_X1    g260(.A(G155gat), .ZN(new_n462));
  INV_X1    g261(.A(G162gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(G155gat), .A2(G162gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT2), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n458), .A2(new_n461), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n450), .A2(G141gat), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n467), .B1(new_n457), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n464), .A2(new_n466), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n449), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n465), .A2(new_n468), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT3), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n473), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n447), .B1(new_n448), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(G22gat), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n482), .ZN(new_n484));
  INV_X1    g283(.A(G22gat), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n484), .B(new_n485), .C1(new_n475), .C2(new_n449), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n440), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n486), .A3(new_n440), .ZN(new_n489));
  OAI211_X1 g288(.A(G228gat), .B(G233gat), .C1(new_n482), .C2(KEYINPUT86), .ZN(new_n490));
  XOR2_X1   g289(.A(G78gat), .B(G106gat), .Z(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT31), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n492), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n488), .A2(new_n489), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  INV_X1    g295(.A(new_n489), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(new_n487), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n479), .A2(new_n400), .A3(new_n473), .A4(new_n402), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n340), .A2(new_n475), .A3(KEYINPUT4), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT3), .B1(new_n469), .B2(new_n474), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n481), .A2(new_n506), .A3(new_n422), .ZN(new_n507));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n505), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n501), .A2(new_n509), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n503), .A2(new_n512), .A3(new_n507), .A4(new_n504), .ZN(new_n513));
  INV_X1    g312(.A(new_n501), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n340), .A2(new_n475), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(KEYINPUT5), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT85), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT85), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n513), .A2(new_n516), .A3(new_n519), .A4(KEYINPUT5), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n511), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522));
  XNOR2_X1  g321(.A(G1gat), .B(G29gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G85gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT0), .B(G57gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n524), .B(new_n525), .Z(new_n526));
  NOR3_X1   g325(.A1(new_n521), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n518), .A2(new_n520), .ZN(new_n528));
  INV_X1    g327(.A(new_n511), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n526), .ZN(new_n531));
  AOI211_X1 g330(.A(new_n531), .B(new_n511), .C1(new_n518), .C2(new_n520), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n527), .B1(new_n533), .B2(new_n522), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT82), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G226gat), .A2(G233gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n421), .A2(new_n448), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n369), .A2(new_n392), .A3(G226gat), .A4(G233gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n447), .ZN(new_n542));
  XOR2_X1   g341(.A(G64gat), .B(G92gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G36gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT80), .B(G8gat), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n544), .B(new_n545), .Z(new_n546));
  INV_X1    g345(.A(new_n447), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n539), .A2(new_n547), .A3(new_n540), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n535), .A2(KEYINPUT82), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n537), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n549), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n542), .A2(new_n548), .ZN(new_n555));
  INV_X1    g354(.A(new_n546), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n557), .A2(KEYINPUT81), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(KEYINPUT81), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n552), .B(new_n554), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n500), .B1(new_n534), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n427), .B1(new_n416), .B2(new_n420), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n434), .A2(new_n426), .A3(new_n435), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n307), .A3(KEYINPUT36), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n439), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT87), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT89), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n530), .A2(new_n532), .A3(KEYINPUT6), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(new_n527), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n527), .A2(new_n569), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n555), .A2(KEYINPUT37), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n574), .B1(new_n576), .B2(new_n546), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(KEYINPUT90), .A3(new_n556), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n555), .A2(KEYINPUT37), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n553), .B1(new_n580), .B2(KEYINPUT38), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n579), .A2(new_n582), .A3(new_n556), .A4(new_n575), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n571), .A2(new_n573), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n505), .A2(new_n507), .ZN(new_n585));
  OR2_X1    g384(.A1(KEYINPUT88), .A2(KEYINPUT39), .ZN(new_n586));
  NAND2_X1  g385(.A1(KEYINPUT88), .A2(KEYINPUT39), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n585), .A2(new_n509), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n514), .A2(new_n515), .A3(new_n509), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n509), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT39), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n588), .B(new_n526), .C1(new_n589), .C2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT40), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n530), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n560), .A4(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n584), .A2(new_n499), .A3(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n439), .A2(new_n561), .A3(KEYINPUT87), .A4(new_n565), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n568), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n499), .A2(new_n562), .A3(new_n563), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT35), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n534), .A2(new_n560), .ZN(new_n605));
  INV_X1    g404(.A(new_n560), .ZN(new_n606));
  INV_X1    g405(.A(new_n532), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n595), .A2(new_n607), .A3(new_n522), .ZN(new_n608));
  INV_X1    g407(.A(new_n527), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT89), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n601), .B(new_n606), .C1(new_n610), .C2(new_n572), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n604), .A2(new_n605), .B1(new_n611), .B2(new_n603), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n306), .B1(new_n600), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n260), .A2(new_n215), .A3(new_n262), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n213), .B(new_n214), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(new_n259), .A3(new_n258), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n263), .A2(KEYINPUT10), .A3(new_n618), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n615), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n614), .B1(new_n616), .B2(new_n619), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n627), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n624), .A2(KEYINPUT101), .A3(new_n627), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n208), .B(G8gat), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n635), .A2(KEYINPUT95), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(KEYINPUT95), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n292), .A2(new_n636), .A3(new_n637), .A4(new_n293), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n283), .A2(new_n281), .A3(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(G229gat), .A2(G233gat), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT18), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n640), .B(KEYINPUT13), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n639), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n635), .B1(new_n283), .B2(new_n281), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n638), .A2(KEYINPUT18), .A3(new_n639), .A4(new_n640), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n651));
  XNOR2_X1  g450(.A(G169gat), .B(G197gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G113gat), .B(G141gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT12), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n643), .A2(new_n656), .A3(new_n648), .A4(new_n649), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n634), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n613), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n534), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g465(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n206), .A2(new_n209), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n664), .A2(new_n560), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G8gat), .B1(new_n663), .B2(new_n606), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(new_n564), .ZN(new_n675));
  AOI21_X1  g474(.A(G15gat), .B1(new_n664), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT36), .B1(new_n564), .B2(new_n307), .ZN(new_n678));
  AOI211_X1 g477(.A(KEYINPUT77), .B(new_n438), .C1(new_n562), .C2(new_n563), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n439), .A2(KEYINPUT102), .A3(new_n565), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(G15gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT103), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n676), .B1(new_n664), .B2(new_n684), .ZN(G1326gat));
  NOR2_X1   g484(.A1(new_n663), .A2(new_n499), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(new_n485), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  AOI21_X1  g488(.A(new_n301), .B1(new_n600), .B2(new_n612), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n662), .A2(new_n303), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n534), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n693), .A2(G29gat), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n611), .A2(new_n603), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n605), .A2(KEYINPUT35), .A3(new_n601), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n598), .A2(new_n561), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n680), .A2(new_n681), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n697), .B1(new_n703), .B2(new_n301), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n600), .A2(new_n612), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(KEYINPUT44), .A3(new_n304), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n692), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n694), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n696), .A2(new_n708), .ZN(G1328gat));
  NOR3_X1   g508(.A1(new_n693), .A2(G36gat), .A3(new_n606), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n707), .B2(new_n606), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n711), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(G1329gat));
  INV_X1    g514(.A(G43gat), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n690), .A2(new_n716), .A3(new_n675), .A4(new_n692), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT106), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT47), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G43gat), .B1(new_n707), .B2(new_n702), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n718), .B(new_n721), .C1(new_n719), .C2(KEYINPUT47), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1330gat));
  NOR3_X1   g524(.A1(new_n693), .A2(G50gat), .A3(new_n499), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n704), .A2(new_n500), .A3(new_n692), .A4(new_n706), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(G50gat), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g528(.A1(new_n302), .A2(new_n305), .A3(new_n661), .A4(new_n634), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n703), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n534), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n560), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n737), .B(new_n738), .Z(G1333gat));
  AOI21_X1  g538(.A(G71gat), .B1(new_n733), .B2(new_n675), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n682), .A2(G71gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n733), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g542(.A1(new_n733), .A2(new_n500), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n239), .A2(new_n660), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n704), .A2(new_n634), .A3(new_n706), .A4(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747), .B2(new_n694), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n598), .A2(new_n561), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n612), .B1(new_n682), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(new_n304), .A3(new_n746), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n750), .A2(KEYINPUT51), .A3(new_n304), .A4(new_n746), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n534), .A2(new_n245), .A3(new_n634), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT108), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n748), .B1(new_n756), .B2(new_n758), .ZN(G1336gat));
  AOI21_X1  g558(.A(new_n633), .B1(new_n753), .B2(new_n754), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n246), .A3(new_n560), .ZN(new_n761));
  OAI21_X1  g560(.A(G92gat), .B1(new_n747), .B2(new_n606), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT52), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n761), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1337gat));
  AOI21_X1  g566(.A(KEYINPUT44), .B1(new_n750), .B2(new_n304), .ZN(new_n768));
  AOI211_X1 g567(.A(new_n697), .B(new_n301), .C1(new_n600), .C2(new_n612), .ZN(new_n769));
  INV_X1    g568(.A(new_n746), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n771), .A2(G99gat), .A3(new_n634), .A4(new_n682), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n760), .A2(new_n675), .ZN(new_n773));
  OAI211_X1 g572(.A(KEYINPUT109), .B(new_n772), .C1(new_n773), .C2(G99gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n775));
  AOI21_X1  g574(.A(G99gat), .B1(new_n760), .B2(new_n675), .ZN(new_n776));
  INV_X1    g575(.A(G99gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n747), .A2(new_n777), .A3(new_n702), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n774), .A2(new_n779), .ZN(G1338gat));
  NAND4_X1  g579(.A1(new_n771), .A2(KEYINPUT110), .A3(new_n634), .A4(new_n500), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n747), .B2(new_n499), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n783), .A3(G106gat), .ZN(new_n784));
  AOI211_X1 g583(.A(G106gat), .B(new_n633), .C1(new_n753), .C2(new_n754), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT53), .B1(new_n785), .B2(new_n500), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G106gat), .B1(new_n747), .B2(new_n499), .ZN(new_n788));
  INV_X1    g587(.A(G106gat), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n755), .A2(new_n789), .A3(new_n634), .A4(new_n500), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(new_n792), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n620), .A2(new_n615), .A3(new_n621), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n622), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT111), .A4(new_n615), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n627), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n622), .B2(new_n794), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT112), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n800), .A2(new_n805), .A3(KEYINPUT55), .A4(new_n802), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n640), .B1(new_n638), .B2(new_n639), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n646), .A2(new_n647), .A3(new_n645), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n655), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n298), .A2(new_n300), .A3(new_n659), .A4(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n624), .A2(new_n627), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n800), .A2(new_n802), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n807), .A2(new_n808), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n804), .A3(new_n806), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT113), .B1(new_n819), .B2(new_n812), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n817), .A2(new_n660), .A3(new_n804), .A4(new_n806), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n631), .A2(new_n659), .A3(new_n632), .A4(new_n811), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n304), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT114), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n301), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n820), .A4(new_n818), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n825), .A2(new_n829), .A3(new_n303), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n302), .A2(new_n305), .A3(new_n661), .A4(new_n633), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n602), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n694), .A2(new_n560), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n661), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(new_n330), .ZN(G1340gat));
  INV_X1    g635(.A(new_n834), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n634), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G120gat), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n327), .A2(new_n328), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n838), .ZN(G1341gat));
  NOR3_X1   g640(.A1(new_n834), .A2(new_n312), .A3(new_n303), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n844));
  AOI21_X1  g643(.A(G127gat), .B1(new_n837), .B2(new_n239), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G1342gat));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n314), .A3(new_n304), .A4(new_n833), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n850), .B2(KEYINPUT56), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n848), .A2(new_n849), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n848), .A2(new_n849), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n852), .A2(KEYINPUT117), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n834), .B2(new_n301), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(G1343gat));
  AOI21_X1  g658(.A(new_n499), .B1(new_n830), .B2(new_n831), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n702), .A2(new_n833), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n303), .B1(new_n821), .B2(new_n824), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n499), .B1(new_n831), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n862), .B(new_n863), .C1(new_n861), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n661), .ZN(new_n867));
  INV_X1    g666(.A(new_n460), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT118), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n860), .A2(new_n863), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n451), .A3(new_n660), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n872), .B1(new_n867), .B2(new_n868), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n869), .A2(new_n873), .A3(KEYINPUT58), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  OAI221_X1 g674(.A(new_n872), .B1(KEYINPUT118), .B2(new_n875), .C1(new_n867), .C2(new_n868), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1344gat));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n450), .A3(new_n634), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n866), .B2(new_n633), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n450), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n863), .B(KEYINPUT119), .Z(new_n882));
  NOR2_X1   g681(.A1(new_n819), .A2(new_n812), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n303), .B1(new_n824), .B2(new_n883), .ZN(new_n884));
  AOI211_X1 g683(.A(KEYINPUT57), .B(new_n499), .C1(new_n831), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n830), .A2(new_n831), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n500), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n885), .B1(new_n887), .B2(KEYINPUT57), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n634), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n879), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n878), .B1(new_n881), .B2(new_n890), .ZN(G1345gat));
  OAI21_X1  g690(.A(new_n462), .B1(new_n870), .B2(new_n303), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n303), .A2(new_n462), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT120), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n892), .B1(new_n866), .B2(new_n894), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT121), .Z(G1346gat));
  OAI21_X1  g695(.A(new_n463), .B1(new_n870), .B2(new_n301), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n304), .A2(G162gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n866), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n534), .A2(new_n606), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n832), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n660), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n634), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g705(.A1(new_n832), .A2(new_n239), .A3(new_n901), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT123), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(KEYINPUT123), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(G183gat), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n902), .A2(new_n239), .A3(new_n356), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT60), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n910), .A2(new_n911), .A3(new_n915), .A4(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1350gat));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n304), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G190gat), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n918), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(KEYINPUT61), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n919), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n923), .B(new_n925), .C1(G190gat), .C2(new_n918), .ZN(G1351gat));
  NAND2_X1  g725(.A1(new_n702), .A2(new_n901), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n888), .A2(KEYINPUT126), .A3(new_n660), .A4(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n831), .A2(new_n884), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n861), .A3(new_n500), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n932), .B(new_n928), .C1(new_n860), .C2(new_n861), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n661), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n929), .A2(G197gat), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n887), .A2(new_n927), .ZN(new_n936));
  INV_X1    g735(.A(G197gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n937), .A3(new_n660), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n935), .A2(KEYINPUT127), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1352gat));
  NOR4_X1   g742(.A1(new_n887), .A2(G204gat), .A3(new_n633), .A4(new_n927), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT62), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n888), .A2(new_n634), .A3(new_n928), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G204gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1353gat));
  OAI21_X1  g747(.A(G211gat), .B1(new_n933), .B2(new_n303), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT63), .Z(new_n950));
  INV_X1    g749(.A(G211gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n936), .A2(new_n951), .A3(new_n239), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n933), .B2(new_n301), .ZN(new_n954));
  INV_X1    g753(.A(G218gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n936), .A2(new_n955), .A3(new_n304), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1355gat));
endmodule


