//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n216), .A2(KEYINPUT64), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n205), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n208), .B1(new_n212), .B2(new_n213), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XOR2_X1   g0032(.A(G87), .B(G97), .Z(new_n233));
  XOR2_X1   g0033(.A(G107), .B(G116), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  NAND3_X1  g0039(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n240));
  AND3_X1   g0040(.A1(new_n240), .A2(KEYINPUT69), .A3(new_n209), .ZN(new_n241));
  AOI21_X1  g0041(.A(KEYINPUT69), .B1(new_n240), .B2(new_n209), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g0043(.A1(G20), .A2(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G68), .ZN(new_n245));
  AOI22_X1  g0045(.A1(new_n244), .A2(G50), .B1(G20), .B2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n210), .A2(G33), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT11), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT75), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n243), .A2(new_n249), .A3(KEYINPUT11), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n256));
  INV_X1    g0056(.A(KEYINPUT12), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT77), .ZN(new_n258));
  INV_X1    g0058(.A(G13), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n259), .A2(new_n210), .A3(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n245), .ZN(new_n261));
  MUX2_X1   g0061(.A(new_n256), .B(new_n258), .S(new_n261), .Z(new_n262));
  AND2_X1   g0062(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n252), .A2(new_n254), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT75), .ZN(new_n265));
  INV_X1    g0065(.A(new_n242), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n240), .A2(KEYINPUT69), .A3(new_n209), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n259), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G20), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n268), .A2(G68), .A3(new_n270), .A4(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT76), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n263), .A2(new_n265), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT78), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT78), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n263), .A2(new_n277), .A3(new_n265), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n284), .A3(G274), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT74), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  AND2_X1   g0087(.A1(G1), .A2(G13), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n283), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT74), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(new_n282), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n284), .A2(KEYINPUT65), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT65), .B1(new_n284), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g0095(.A(G238), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n299));
  INV_X1    g0099(.A(G226), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT66), .ZN(new_n302));
  AND2_X1   g0102(.A1(KEYINPUT3), .A2(G33), .ZN(new_n303));
  NOR2_X1   g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT3), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(KEYINPUT66), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n301), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT73), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n305), .A2(new_n310), .A3(G232), .A4(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT73), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n301), .A2(new_n305), .A3(new_n310), .A4(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n284), .ZN(new_n318));
  AOI211_X1 g0118(.A(KEYINPUT13), .B(new_n297), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n318), .ZN(new_n321));
  INV_X1    g0121(.A(new_n297), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G190), .ZN(new_n325));
  OAI21_X1  g0125(.A(G200), .B1(new_n319), .B2(new_n323), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n279), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(G169), .B1(new_n319), .B2(new_n323), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT14), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(G169), .C1(new_n319), .C2(new_n323), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT79), .B1(new_n324), .B2(G179), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT79), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NOR4_X1   g0134(.A1(new_n319), .A2(new_n323), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n329), .B(new_n331), .C1(new_n332), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n279), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n327), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n303), .A2(new_n304), .A3(new_n302), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT66), .B1(new_n308), .B2(new_n309), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n298), .A2(new_n299), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(G222), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(G223), .A3(G1698), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n344), .C1(new_n247), .C2(new_n341), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n318), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT68), .ZN(new_n347));
  INV_X1    g0147(.A(new_n285), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n294), .A2(new_n295), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(G226), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(new_n346), .B2(new_n350), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n334), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n243), .A2(new_n260), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n272), .A2(G50), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT70), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT8), .B(G58), .ZN(new_n359));
  INV_X1    g0159(.A(G150), .ZN(new_n360));
  INV_X1    g0160(.A(new_n244), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n359), .A2(new_n248), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G50), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n210), .B1(new_n201), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n243), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n358), .B(new_n365), .C1(G50), .C2(new_n270), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n346), .A2(new_n350), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT68), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(new_n351), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n354), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(G190), .B1(new_n352), .B2(new_n353), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(G200), .A3(new_n351), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n366), .B(KEYINPUT9), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n373), .A2(new_n374), .A3(new_n375), .A4(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n372), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n359), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n244), .B1(G20), .B2(G77), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n248), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n243), .B1(new_n247), .B2(new_n260), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n355), .A2(G77), .A3(new_n272), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n305), .A2(new_n310), .A3(G232), .A4(new_n342), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n305), .A2(new_n310), .A3(G238), .A4(G1698), .ZN(new_n389));
  INV_X1    g0189(.A(G107), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n388), .B(new_n389), .C1(new_n341), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n318), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n348), .B1(new_n349), .B2(G244), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT71), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n392), .B2(new_n393), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n387), .B1(new_n397), .B2(G200), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT72), .B(G190), .C1(new_n395), .C2(new_n396), .ZN(new_n399));
  OAI21_X1  g0199(.A(G190), .B1(new_n395), .B2(new_n396), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n398), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n359), .B1(new_n271), .B2(G20), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n355), .A2(new_n404), .B1(new_n260), .B2(new_n359), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  NOR4_X1   g0206(.A1(new_n303), .A2(new_n304), .A3(new_n406), .A4(G20), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(G20), .B1(new_n305), .B2(new_n310), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(KEYINPUT7), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G68), .ZN(new_n411));
  INV_X1    g0211(.A(G58), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n245), .ZN(new_n413));
  OAI21_X1  g0213(.A(G20), .B1(new_n413), .B2(new_n201), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n244), .A2(G159), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT16), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n303), .A2(new_n304), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT7), .B1(new_n419), .B2(new_n210), .ZN(new_n420));
  OAI21_X1  g0220(.A(G68), .B1(new_n420), .B2(new_n407), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(KEYINPUT16), .A3(new_n417), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n243), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n405), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT67), .ZN(new_n425));
  INV_X1    g0225(.A(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(G223), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G226), .A2(G1698), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n419), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G87), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n307), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n318), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT80), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n284), .A2(new_n293), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(G232), .B1(new_n289), .B2(new_n282), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n434), .A2(new_n435), .A3(new_n334), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n429), .A2(new_n430), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n308), .A2(new_n309), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n433), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n334), .B(new_n437), .C1(new_n441), .C2(new_n284), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT80), .ZN(new_n443));
  AOI21_X1  g0243(.A(G169), .B1(new_n434), .B2(new_n437), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n438), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n424), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT18), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n424), .A2(new_n448), .A3(new_n445), .ZN(new_n449));
  INV_X1    g0249(.A(G190), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n434), .A2(new_n450), .A3(new_n437), .ZN(new_n451));
  INV_X1    g0251(.A(G232), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n284), .A2(new_n293), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n285), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n433), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n342), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n419), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n457), .B2(new_n318), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n451), .B1(new_n458), .B2(G200), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n405), .C1(new_n418), .C2(new_n423), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT17), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n416), .B1(new_n410), .B2(G68), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n243), .B(new_n422), .C1(new_n463), .C2(KEYINPUT16), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(KEYINPUT17), .A3(new_n405), .A4(new_n459), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n447), .A2(new_n449), .A3(new_n462), .A4(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n334), .B1(new_n395), .B2(new_n396), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n392), .A2(new_n393), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT71), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n369), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n471), .A3(new_n387), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n403), .A2(new_n466), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n338), .A2(new_n380), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n281), .A2(G1), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G257), .A3(new_n284), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n289), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(new_n480), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n305), .A2(new_n310), .A3(G250), .A4(G1698), .ZN(new_n487));
  AND2_X1   g0287(.A1(KEYINPUT4), .A2(G244), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n305), .A2(new_n310), .A3(new_n342), .A4(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  OAI21_X1  g0290(.A(G244), .B1(new_n303), .B2(new_n304), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n427), .A2(new_n428), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n487), .A2(new_n489), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n318), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n486), .A2(new_n496), .A3(new_n334), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT82), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n486), .A2(new_n496), .A3(new_n499), .A4(new_n334), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n390), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n390), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G97), .A2(G107), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n502), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(G20), .B1(G77), .B2(new_n244), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n210), .B1(new_n339), .B2(new_n340), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n407), .B1(new_n509), .B2(new_n406), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n510), .B2(new_n390), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n243), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n260), .A2(new_n503), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n271), .A2(G33), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n270), .B(new_n514), .C1(new_n241), .C2(new_n242), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n515), .B2(new_n503), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n486), .A2(new_n496), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n512), .A2(new_n517), .B1(new_n518), .B2(new_n369), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n501), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(G200), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n516), .B1(new_n511), .B2(new_n243), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n450), .C2(new_n518), .ZN(new_n523));
  INV_X1    g0323(.A(new_n383), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(new_n270), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n268), .A2(new_n270), .A3(new_n524), .A4(new_n514), .ZN(new_n527));
  AOI21_X1  g0327(.A(G20), .B1(new_n308), .B2(new_n309), .ZN(new_n528));
  XNOR2_X1  g0328(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n528), .A2(G68), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n505), .A2(new_n432), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT84), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT84), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT19), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n313), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n537), .B2(G20), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n526), .B(new_n527), .C1(new_n539), .C2(new_n268), .ZN(new_n540));
  OAI211_X1 g0340(.A(G244), .B(G1698), .C1(new_n303), .C2(new_n304), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT83), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n440), .A2(KEYINPUT83), .A3(G244), .A4(G1698), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n440), .A2(new_n342), .A3(G238), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n318), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n271), .A2(G45), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n549), .A2(G250), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n284), .ZN(new_n551));
  INV_X1    g0351(.A(new_n289), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n549), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n548), .A2(new_n334), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n547), .B2(new_n318), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n540), .B(new_n555), .C1(G169), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n548), .A2(G190), .A3(new_n554), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n268), .B1(new_n531), .B2(new_n538), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n515), .A2(new_n432), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n559), .A2(new_n560), .A3(new_n525), .ZN(new_n561));
  INV_X1    g0361(.A(G200), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n558), .B(new_n561), .C1(new_n562), .C2(new_n556), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n520), .A2(new_n523), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT86), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n260), .A2(new_n390), .ZN(new_n567));
  XNOR2_X1  g0367(.A(new_n567), .B(KEYINPUT25), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n515), .A2(new_n390), .ZN(new_n569));
  OR2_X1    g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n432), .A2(KEYINPUT22), .A3(G20), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n305), .A2(new_n310), .A3(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n210), .B(G87), .C1(new_n303), .C2(new_n304), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT22), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n546), .A2(G20), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n210), .B2(G107), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n390), .A2(KEYINPUT23), .A3(G20), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT24), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n575), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n570), .B1(new_n585), .B2(new_n243), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n479), .A2(G264), .A3(new_n284), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n483), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n440), .A2(new_n342), .A3(G250), .ZN(new_n589));
  AND2_X1   g0389(.A1(G257), .A2(G1698), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n303), .B2(new_n304), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT85), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT85), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n440), .A2(new_n593), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(G33), .A2(G294), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n589), .A2(new_n592), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n588), .B1(new_n596), .B2(new_n318), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n334), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(G169), .B2(new_n597), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n566), .B1(new_n586), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT87), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n597), .B2(new_n450), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G200), .B2(new_n597), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n597), .A2(new_n601), .A3(new_n450), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n586), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n597), .A2(G169), .ZN(new_n606));
  AOI211_X1 g0406(.A(G179), .B(new_n588), .C1(new_n318), .C2(new_n596), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n575), .A2(new_n583), .A3(new_n580), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n583), .B1(new_n575), .B2(new_n580), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n243), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n568), .A2(new_n569), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n608), .A2(new_n613), .A3(KEYINPUT86), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n600), .A2(new_n605), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(G116), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n269), .A2(G20), .A3(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n240), .A2(new_n209), .B1(G20), .B2(new_n616), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n494), .B(new_n210), .C1(G33), .C2(new_n503), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n618), .A2(KEYINPUT20), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT20), .B1(new_n618), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n515), .A2(new_n616), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT21), .ZN(new_n626));
  INV_X1    g0426(.A(G303), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n305), .B2(new_n310), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n427), .A2(G257), .A3(new_n428), .ZN(new_n629));
  NAND2_X1  g0429(.A1(G264), .A2(G1698), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n419), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n318), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n482), .A2(new_n476), .B1(new_n288), .B2(new_n283), .ZN(new_n633));
  INV_X1    g0433(.A(new_n478), .ZN(new_n634));
  NAND2_X1  g0434(.A1(KEYINPUT5), .A2(G41), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n549), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n633), .A2(G270), .B1(new_n289), .B2(new_n636), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n626), .B(new_n369), .C1(new_n632), .C2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n632), .A2(G179), .A3(new_n637), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n625), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n632), .A2(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G169), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n626), .B1(new_n642), .B2(new_n624), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(G200), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n646), .B(new_n624), .C1(new_n450), .C2(new_n641), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NOR4_X1   g0448(.A1(new_n475), .A2(new_n565), .A3(new_n615), .A4(new_n648), .ZN(G372));
  INV_X1    g0449(.A(KEYINPUT91), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n462), .A2(new_n465), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n332), .A2(new_n335), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n329), .A2(new_n331), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n337), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n279), .A2(new_n325), .A3(new_n326), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n473), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n652), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n424), .A2(new_n448), .A3(new_n445), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n448), .B1(new_n424), .B2(new_n445), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n650), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n377), .A2(new_n379), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n336), .A2(new_n337), .B1(new_n656), .B2(new_n473), .ZN(new_n665));
  OAI211_X1 g0465(.A(KEYINPUT91), .B(new_n661), .C1(new_n665), .C2(new_n652), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(new_n371), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n520), .A2(new_n523), .A3(new_n564), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n586), .A2(new_n599), .A3(KEYINPUT88), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT88), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n608), .B2(new_n613), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n645), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT89), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n669), .A2(new_n673), .A3(new_n674), .A4(new_n605), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n520), .A2(new_n564), .A3(new_n523), .A4(new_n605), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT88), .B1(new_n586), .B2(new_n599), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n608), .A2(new_n613), .A3(new_n671), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n644), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT89), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n557), .A2(new_n563), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n520), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n564), .A2(KEYINPUT26), .A3(new_n501), .A4(new_n519), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n557), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT90), .ZN(new_n688));
  INV_X1    g0488(.A(new_n557), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n684), .B2(new_n685), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n681), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n668), .B1(new_n475), .B2(new_n693), .ZN(G369));
  INV_X1    g0494(.A(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n269), .A2(new_n695), .A3(new_n210), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT92), .ZN(new_n697));
  INV_X1    g0497(.A(G213), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n269), .A2(new_n210), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(G343), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT93), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n624), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT94), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n644), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n648), .B2(new_n705), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT95), .Z(new_n708));
  INV_X1    g0508(.A(new_n703), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n613), .A3(new_n608), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n586), .A2(new_n703), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n615), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(G330), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n677), .A2(new_n678), .A3(new_n703), .ZN(new_n714));
  INV_X1    g0514(.A(new_n615), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n645), .A2(new_n709), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n713), .A2(new_n714), .A3(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n206), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n532), .A2(G116), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n213), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  INV_X1    g0525(.A(G330), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n703), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n518), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n596), .A2(new_n318), .B1(G264), .B2(new_n633), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n556), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n729), .A2(new_n731), .A3(KEYINPUT30), .A4(new_n639), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n597), .A2(G179), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n548), .A2(new_n554), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n518), .A3(new_n734), .A4(new_n641), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n632), .A2(new_n637), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(G179), .A3(new_n556), .A4(new_n730), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n739), .B2(new_n518), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n728), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  AND4_X1   g0542(.A1(new_n643), .A2(new_n640), .A3(new_n647), .A4(new_n703), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n600), .A3(new_n614), .A4(new_n605), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n742), .B1(new_n744), .B2(new_n565), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(KEYINPUT96), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT96), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n748), .B(new_n737), .C1(new_n739), .C2(new_n518), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n736), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n727), .B1(new_n750), .B2(new_n703), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n726), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT29), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n693), .B2(new_n709), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n600), .A2(new_n614), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n676), .B1(new_n755), .B2(new_n645), .ZN(new_n756));
  OAI211_X1 g0556(.A(KEYINPUT29), .B(new_n703), .C1(new_n687), .C2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n752), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n725), .B1(new_n758), .B2(G1), .ZN(G364));
  NOR2_X1   g0559(.A1(new_n259), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n271), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OR3_X1    g0562(.A1(new_n720), .A2(new_n762), .A3(KEYINPUT97), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT97), .B1(new_n720), .B2(new_n762), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n708), .B2(G330), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n708), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT98), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n210), .A2(new_n334), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n450), .A2(new_n562), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n562), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G326), .A2(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n210), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n771), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n770), .A2(new_n782), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n778), .B1(new_n627), .B2(new_n780), .C1(new_n781), .C2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n450), .A2(G179), .A3(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n210), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n341), .B(new_n784), .C1(G294), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n779), .A2(new_n782), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G329), .ZN(new_n791));
  INV_X1    g0591(.A(new_n770), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n792), .A2(new_n450), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G322), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n779), .A2(new_n774), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(G283), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n341), .ZN(new_n800));
  INV_X1    g0600(.A(new_n780), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G87), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n794), .B2(new_n412), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n800), .B(new_n803), .C1(G97), .C2(new_n787), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n783), .A2(new_n247), .B1(new_n797), .B2(new_n390), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n772), .A2(new_n363), .B1(new_n775), .B2(new_n245), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT32), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n789), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n790), .A2(KEYINPUT32), .A3(G159), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n805), .B(new_n806), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n788), .A2(new_n799), .B1(new_n804), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n209), .B1(G20), .B2(new_n369), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n766), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n813), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT99), .Z(new_n820));
  NOR2_X1   g0620(.A1(new_n800), .A2(new_n719), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n821), .A2(G355), .B1(new_n616), .B2(new_n719), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n238), .A2(G45), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n719), .A2(new_n440), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(G45), .C2(new_n213), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n820), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n815), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n818), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n708), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n769), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  NAND2_X1  g0631(.A1(new_n709), .A2(new_n387), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n472), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n398), .A2(new_n399), .A3(new_n402), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n833), .A2(new_n834), .B1(new_n473), .B2(new_n709), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n693), .B2(new_n709), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n691), .B1(new_n686), .B2(new_n557), .ZN(new_n837));
  AOI211_X1 g0637(.A(KEYINPUT90), .B(new_n689), .C1(new_n684), .C2(new_n685), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n675), .B(new_n680), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n472), .A2(new_n832), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n403), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n709), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n752), .B1(new_n836), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n763), .B2(new_n764), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n836), .A2(new_n752), .A3(new_n844), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n772), .A2(new_n627), .B1(new_n789), .B2(new_n781), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G294), .B2(new_n793), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n341), .B1(G97), .B2(new_n787), .ZN(new_n851));
  INV_X1    g0651(.A(new_n783), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G116), .A2(new_n852), .B1(new_n798), .B2(G87), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G107), .A2(new_n801), .B1(new_n776), .B2(G283), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n850), .A2(new_n851), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT100), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G150), .A2(new_n776), .B1(new_n852), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  XNOR2_X1  g0658(.A(KEYINPUT101), .B(G143), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n857), .B1(new_n858), .B2(new_n772), .C1(new_n794), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT34), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n440), .B1(new_n789), .B2(new_n863), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n780), .A2(new_n363), .B1(new_n797), .B2(new_n245), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n864), .B(new_n865), .C1(G58), .C2(new_n787), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n860), .A2(new_n861), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n856), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n855), .A2(KEYINPUT100), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n813), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n813), .A2(new_n816), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n765), .B1(new_n247), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n473), .A2(new_n709), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n403), .B2(new_n840), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n871), .B(new_n873), .C1(new_n875), .C2(new_n817), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n848), .A2(new_n876), .ZN(G384));
  AOI211_X1 g0677(.A(new_n616), .B(new_n212), .C1(new_n507), .C2(KEYINPUT35), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(KEYINPUT35), .B2(new_n507), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  OR3_X1    g0680(.A1(new_n213), .A2(new_n247), .A3(new_n413), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n363), .A2(G68), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n271), .B(G13), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n667), .A2(new_n371), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT29), .B1(new_n839), .B2(new_n703), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n757), .A2(new_n338), .A3(new_n380), .A4(new_n474), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT102), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT102), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n703), .B1(new_n687), .B2(new_n756), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n475), .B1(new_n891), .B2(KEYINPUT29), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n754), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n885), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n697), .A2(new_n700), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n662), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT16), .B1(new_n421), .B2(new_n417), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n405), .B1(new_n423), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n895), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n661), .B2(new_n651), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n445), .A2(new_n899), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n460), .A3(new_n901), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n424), .A2(new_n900), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n446), .A2(new_n906), .A3(new_n907), .A4(new_n460), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n897), .B1(new_n902), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n901), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n466), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n905), .A2(new_n908), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT39), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n336), .A2(new_n337), .A3(new_n703), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n906), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n446), .A2(new_n906), .A3(new_n460), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT37), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n466), .A2(new_n920), .B1(new_n922), .B2(new_n908), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n914), .B1(new_n923), .B2(KEYINPUT38), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n917), .A2(new_n919), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n472), .A2(new_n709), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n843), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n929), .B1(new_n693), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n337), .A2(new_n709), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n655), .A2(new_n656), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n337), .B(new_n709), .C1(new_n327), .C2(new_n336), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n896), .B(new_n927), .C1(new_n936), .C2(new_n916), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n894), .B(new_n937), .Z(new_n938));
  NAND4_X1  g0738(.A1(new_n640), .A2(new_n647), .A3(new_n643), .A4(new_n703), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n615), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n739), .A2(new_n518), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n596), .A2(new_n318), .ZN(new_n942));
  INV_X1    g0742(.A(new_n588), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND4_X1   g0744(.A1(new_n334), .A2(new_n734), .A3(new_n944), .A4(new_n641), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n941), .A2(KEYINPUT30), .B1(new_n945), .B2(new_n518), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n729), .A2(new_n731), .A3(new_n639), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n748), .B1(new_n947), .B2(new_n737), .ZN(new_n948));
  INV_X1    g0748(.A(new_n749), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n940), .A2(new_n669), .B1(new_n950), .B2(new_n728), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n835), .B1(new_n951), .B2(new_n751), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n935), .A2(new_n915), .A3(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT40), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n935), .A2(new_n924), .A3(new_n952), .A4(KEYINPUT40), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n475), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n951), .A2(new_n751), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n957), .A2(new_n960), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(G330), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n938), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n271), .B2(new_n760), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n938), .A2(new_n963), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n884), .B1(new_n965), .B2(new_n966), .ZN(G367));
  INV_X1    g0767(.A(new_n820), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n206), .B2(new_n383), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n231), .A2(new_n719), .A3(new_n440), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n766), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G294), .A2(new_n776), .B1(new_n790), .B2(G317), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n781), .B2(new_n772), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n794), .A2(new_n627), .B1(new_n797), .B2(new_n503), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT46), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n780), .B2(new_n616), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n975), .B(new_n977), .C1(new_n390), .C2(new_n786), .ZN(new_n978));
  INV_X1    g0778(.A(G283), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n419), .B1(new_n783), .B2(new_n979), .ZN(new_n980));
  NOR4_X1   g0780(.A1(new_n973), .A2(new_n974), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n793), .A2(G150), .B1(G50), .B2(new_n852), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n772), .B2(new_n859), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n341), .B1(new_n245), .B2(new_n786), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n797), .A2(new_n247), .B1(new_n789), .B2(new_n858), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n412), .A2(new_n780), .B1(new_n775), .B2(new_n808), .ZN(new_n986));
  NOR4_X1   g0786(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT47), .Z(new_n989));
  AOI21_X1  g0789(.A(new_n971), .B1(new_n989), .B2(new_n813), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n703), .A2(new_n561), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n564), .B(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n990), .B1(new_n993), .B2(new_n828), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n708), .A2(G330), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n717), .B1(new_n712), .B2(new_n716), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n995), .B(new_n996), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n758), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n717), .A2(new_n714), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n520), .B(new_n523), .C1(new_n522), .C2(new_n703), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n501), .A2(new_n519), .A3(new_n709), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT45), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n999), .A2(new_n1002), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT44), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(new_n713), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n713), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n758), .B1(new_n998), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n720), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n762), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1002), .A2(new_n717), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT42), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n755), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n523), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n709), .B1(new_n1018), .B2(new_n520), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n1015), .B2(KEYINPUT42), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1016), .A2(new_n1020), .B1(KEYINPUT43), .B2(new_n993), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n713), .A2(new_n1002), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n994), .B1(new_n1014), .B2(new_n1025), .ZN(G387));
  NAND2_X1  g0826(.A1(new_n997), .A2(new_n762), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT103), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n997), .A2(KEYINPUT103), .A3(new_n762), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n712), .A2(new_n828), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n381), .A2(new_n363), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n722), .B(new_n281), .C1(new_n245), .C2(new_n247), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n824), .B1(new_n1033), .B2(new_n1034), .C1(new_n228), .C2(new_n281), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n722), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n821), .A2(new_n1036), .B1(new_n390), .B2(new_n719), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(KEYINPUT104), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n968), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT104), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n766), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n794), .A2(new_n363), .B1(new_n783), .B2(new_n245), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n381), .B2(new_n776), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n780), .A2(new_n247), .B1(new_n789), .B2(new_n360), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT105), .Z(new_n1045));
  NOR2_X1   g0845(.A1(new_n772), .A2(new_n808), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT106), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n786), .A2(new_n383), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n419), .B(new_n1048), .C1(G97), .C2(new_n798), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n440), .B1(new_n790), .B2(G326), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n793), .A2(G317), .B1(new_n773), .B2(G322), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n627), .B2(new_n783), .C1(new_n781), .C2(new_n775), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT108), .Z(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  INV_X1    g0857(.A(G294), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n786), .A2(new_n979), .B1(new_n780), .B2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT107), .Z(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT49), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1051), .B1(new_n616), .B2(new_n797), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1050), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1041), .B1(new_n1065), .B2(new_n813), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n997), .A2(new_n758), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n998), .A2(new_n720), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(G393));
  NAND3_X1  g0870(.A1(new_n1008), .A2(KEYINPUT109), .A3(new_n1009), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT109), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1007), .A2(new_n1072), .A3(new_n713), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT110), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n761), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n1075), .B2(new_n1074), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1071), .A2(new_n998), .A3(new_n1073), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1078), .B(new_n720), .C1(new_n998), .C2(new_n1010), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n235), .A2(new_n824), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n968), .B(new_n1080), .C1(new_n503), .C2(new_n206), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n766), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT111), .Z(new_n1083));
  OAI22_X1  g0883(.A1(new_n775), .A2(new_n627), .B1(new_n797), .B2(new_n390), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n341), .B(new_n1084), .C1(G116), .C2(new_n787), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G283), .A2(new_n801), .B1(new_n790), .B2(G322), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n1058), .C2(new_n783), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n793), .A2(G311), .B1(new_n773), .B2(G317), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n780), .A2(new_n245), .B1(new_n789), .B2(new_n859), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n419), .B(new_n1091), .C1(G87), .C2(new_n798), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT112), .Z(new_n1093));
  AOI22_X1  g0893(.A1(new_n793), .A2(G159), .B1(new_n773), .B2(G150), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT51), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n787), .A2(G77), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n363), .B2(new_n775), .C1(new_n359), .C2(new_n783), .ZN(new_n1097));
  OR3_X1    g0897(.A1(new_n1093), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1090), .B1(new_n1098), .B2(KEYINPUT113), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(KEYINPUT113), .B2(new_n1098), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1083), .B1(new_n1100), .B2(new_n813), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1002), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n828), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1077), .A2(new_n1079), .A3(new_n1103), .ZN(G390));
  NAND3_X1  g0904(.A1(new_n959), .A2(G330), .A3(new_n875), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n935), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n928), .B1(new_n839), .B2(new_n843), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n933), .A2(new_n934), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n918), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n917), .A2(new_n926), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n924), .A2(new_n918), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n929), .B1(new_n890), .B2(new_n842), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n935), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1107), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n752), .A2(new_n935), .A3(new_n875), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1119), .B(new_n1115), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n958), .A2(G330), .A3(new_n959), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n889), .B1(new_n754), .B2(new_n892), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n886), .A2(KEYINPUT102), .A3(new_n887), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n668), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT31), .B1(new_n950), .B2(new_n709), .ZN(new_n1126));
  OAI211_X1 g0926(.A(G330), .B(new_n875), .C1(new_n745), .C2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n933), .A3(new_n934), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1109), .B2(new_n1105), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n931), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1109), .A2(new_n1105), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1114), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(new_n1118), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1125), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n721), .B1(new_n1121), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1115), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1118), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1107), .B2(new_n1138), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n894), .A2(new_n1122), .A3(new_n1134), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1140), .A2(KEYINPUT114), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(KEYINPUT114), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1137), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n872), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n794), .A2(new_n863), .B1(new_n797), .B2(new_n363), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n800), .B(new_n1146), .C1(G159), .C2(new_n787), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n801), .A2(G150), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT53), .ZN(new_n1149));
  INV_X1    g0949(.A(G128), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT54), .B(G143), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n772), .A2(new_n1150), .B1(new_n783), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n775), .A2(new_n858), .B1(new_n789), .B2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1149), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n800), .A2(new_n802), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT116), .Z(new_n1157));
  OAI221_X1 g0957(.A(new_n1096), .B1(new_n245), .B2(new_n797), .C1(new_n1058), .C2(new_n789), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n772), .A2(new_n979), .B1(new_n783), .B2(new_n503), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n794), .A2(new_n616), .B1(new_n775), .B2(new_n390), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1147), .A2(new_n1155), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n766), .B1(new_n381), .B2(new_n1145), .C1(new_n1162), .C2(new_n814), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1111), .B2(new_n816), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT115), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1140), .B2(new_n761), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1121), .A2(KEYINPUT115), .A3(new_n762), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1164), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1144), .A2(new_n1168), .ZN(G378));
  XNOR2_X1  g0969(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n366), .A2(new_n900), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n380), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n380), .A2(new_n1172), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1171), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1175), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n1173), .A3(new_n1170), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT117), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n728), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n744), .A2(new_n565), .B1(new_n750), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n875), .B1(new_n1182), .B2(new_n1126), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n933), .B2(new_n934), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT40), .B1(new_n1184), .B2(new_n915), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n956), .A2(G330), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1179), .B(new_n1180), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n955), .A2(KEYINPUT117), .A3(G330), .A4(new_n956), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1179), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n924), .A2(KEYINPUT40), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n726), .B1(new_n1191), .B2(new_n1184), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT117), .B1(new_n1192), .B2(new_n955), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1187), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n937), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n937), .B(new_n1187), .C1(new_n1190), .C2(new_n1193), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n762), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n765), .B1(new_n363), .B2(new_n872), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n794), .A2(new_n1150), .B1(new_n772), .B2(new_n1153), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1151), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G132), .A2(new_n776), .B1(new_n801), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n360), .B2(new_n786), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1201), .B(new_n1204), .C1(G137), .C2(new_n852), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n307), .B(new_n280), .C1(new_n797), .C2(new_n808), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G124), .B2(new_n790), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n419), .A2(new_n280), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n798), .A2(G58), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n383), .B2(new_n783), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1212), .B(new_n1214), .C1(G77), .C2(new_n801), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n245), .B2(new_n786), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n794), .A2(new_n390), .B1(new_n789), .B2(new_n979), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n772), .A2(new_n616), .B1(new_n775), .B2(new_n503), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(KEYINPUT58), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(KEYINPUT58), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1212), .B(new_n363), .C1(G33), .C2(G41), .ZN(new_n1222));
  AND4_X1   g1022(.A1(new_n1211), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1200), .B1(new_n814), .B2(new_n1223), .C1(new_n1179), .C2(new_n817), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1199), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1197), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1180), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n937), .B1(new_n1229), .B2(new_n1187), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT57), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1125), .B1(new_n1121), .B2(new_n1136), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT118), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1125), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT118), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1235), .A2(new_n1198), .A3(new_n1236), .A4(KEYINPUT57), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1138), .A2(new_n1107), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1136), .A2(new_n1239), .A3(new_n1139), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1240), .A2(new_n1234), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n720), .B1(new_n1241), .B2(KEYINPUT57), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1226), .B1(new_n1238), .B2(new_n1242), .ZN(G375));
  INV_X1    g1043(.A(KEYINPUT119), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1244), .B(new_n1134), .C1(new_n894), .C2(new_n1122), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT119), .B1(new_n1125), .B2(new_n1135), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n1013), .A3(new_n1141), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n935), .A2(new_n817), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT120), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n765), .B1(new_n245), .B2(new_n872), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n786), .A2(new_n363), .B1(new_n783), .B2(new_n360), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT121), .Z(new_n1253));
  AOI22_X1  g1053(.A1(new_n793), .A2(G137), .B1(new_n776), .B2(new_n1202), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1150), .B2(new_n789), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G132), .A2(new_n773), .B1(new_n801), .B2(G159), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n440), .A3(new_n1213), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1253), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n772), .A2(new_n1058), .B1(new_n775), .B2(new_n616), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G107), .B2(new_n852), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(G77), .A2(new_n798), .B1(new_n790), .B2(G303), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1261), .B1(new_n503), .B2(new_n780), .C1(new_n979), .C2(new_n794), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1262), .A2(new_n341), .A3(new_n1048), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1258), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1250), .B(new_n1251), .C1(new_n814), .C2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1135), .B2(new_n761), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1248), .A2(new_n1267), .ZN(G381));
  NOR3_X1   g1068(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT122), .Z(new_n1270));
  OR2_X1    g1070(.A1(G375), .A2(G378), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G390), .A2(G387), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  OR4_X1    g1073(.A1(G381), .A2(new_n1270), .A3(new_n1271), .A4(new_n1273), .ZN(G407));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(G343), .C2(new_n1271), .ZN(G409));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n698), .A2(G343), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G378), .B(new_n1226), .C1(new_n1238), .C2(new_n1242), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1241), .A2(new_n1013), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1144), .B(new_n1168), .C1(new_n1279), .C2(new_n1225), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1277), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1277), .ZN(new_n1282));
  INV_X1    g1082(.A(G2897), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1125), .A2(new_n1135), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1244), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1125), .A2(KEYINPUT119), .A3(new_n1135), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1134), .B1(new_n894), .B2(new_n1122), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n721), .B1(new_n1291), .B2(KEYINPUT60), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G384), .B1(new_n1293), .B2(new_n1267), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1295), .B(new_n1266), .C1(new_n1290), .C2(new_n1292), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1285), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n720), .B1(new_n1286), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n1247), .B2(new_n1289), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1295), .B1(new_n1300), .B2(new_n1266), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1293), .A2(G384), .A3(new_n1267), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1284), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1297), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1276), .B1(new_n1281), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(KEYINPUT126), .B(new_n1276), .C1(new_n1281), .C2(new_n1304), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1281), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT62), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1281), .A2(new_n1312), .A3(new_n1309), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1307), .A2(new_n1308), .A3(new_n1311), .A4(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(G393), .B(new_n830), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G390), .A2(G387), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1273), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1317), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1315), .B1(new_n1319), .B2(new_n1272), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1314), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1297), .A2(new_n1303), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT125), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1323), .B(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT124), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1281), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1281), .A2(new_n1326), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1325), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1310), .A2(KEYINPUT123), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(KEYINPUT63), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1321), .A2(KEYINPUT61), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1310), .A2(KEYINPUT123), .A3(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1329), .A2(new_n1331), .A3(new_n1332), .A4(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1322), .A2(new_n1335), .ZN(G405));
  NAND3_X1  g1136(.A1(G375), .A2(new_n1144), .A3(new_n1168), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1278), .ZN(new_n1338));
  OR2_X1    g1138(.A1(new_n1338), .A2(new_n1309), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1318), .A2(new_n1320), .A3(KEYINPUT127), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1338), .A2(new_n1309), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1339), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT127), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(new_n1343), .A3(new_n1321), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1321), .A2(new_n1343), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1345), .A2(new_n1339), .A3(new_n1340), .A4(new_n1341), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(G402));
endmodule


