//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n463), .A2(new_n468), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n468), .B2(G112), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n475), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT66), .A2(G114), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT66), .A2(G114), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT67), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2105), .C1(new_n484), .C2(new_n485), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n468), .C1(new_n461), .C2(new_n462), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n468), .B(new_n497), .C1(new_n461), .C2(new_n462), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n492), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n502), .B(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G62), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n505), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n509), .A2(new_n511), .A3(G543), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(KEYINPUT68), .ZN(new_n519));
  OAI221_X1 g094(.A(KEYINPUT68), .B1(new_n515), .B2(new_n516), .C1(new_n513), .C2(new_n514), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n508), .B1(new_n519), .B2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND3_X1  g098(.A1(new_n512), .A2(G89), .A3(new_n505), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n509), .A2(new_n511), .A3(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(G51), .B1(new_n505), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n525), .B1(new_n524), .B2(new_n527), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  NAND3_X1  g109(.A1(new_n512), .A2(G90), .A3(new_n505), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OAI221_X1 g112(.A(new_n535), .B1(new_n536), .B2(new_n516), .C1(new_n537), .C2(new_n501), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  XOR2_X1   g114(.A(KEYINPUT71), .B(G43), .Z(new_n540));
  NAND2_X1  g115(.A1(new_n529), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n513), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n501), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT72), .ZN(G176));
  XOR2_X1   g124(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n550));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  AOI22_X1  g128(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(new_n501), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n509), .A2(new_n511), .A3(G53), .A4(G543), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT74), .B1(new_n513), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n512), .A2(new_n562), .A3(G91), .A4(new_n505), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n559), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  NAND2_X1  g141(.A1(new_n529), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n568));
  INV_X1    g143(.A(G87), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n567), .B(new_n568), .C1(new_n513), .C2(new_n569), .ZN(G288));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n513), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n512), .A2(KEYINPUT76), .A3(G86), .A4(new_n505), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(G48), .A2(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n509), .A2(new_n511), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n509), .A2(new_n511), .A3(new_n576), .A4(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g156(.A1(KEYINPUT5), .A2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(KEYINPUT5), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G61), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n584), .A2(new_n585), .B1(G73), .B2(G543), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n505), .A2(KEYINPUT75), .A3(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n581), .B1(new_n588), .B2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n575), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n529), .A2(G47), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n591), .B1(new_n513), .B2(new_n592), .C1(new_n501), .C2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n513), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n512), .A2(KEYINPUT10), .A3(G92), .A4(new_n505), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n582), .A2(new_n583), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  INV_X1    g180(.A(G543), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n603), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI221_X1 g184(.A(KEYINPUT79), .B1(new_n605), .B2(new_n606), .C1(new_n603), .C2(new_n604), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(G651), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n529), .A2(G54), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n602), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n597), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n597), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(G299), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n617), .B2(G168), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(new_n617), .B2(G168), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n614), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n478), .A2(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n478), .A2(G135), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT80), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n474), .A2(G123), .ZN(new_n635));
  NOR2_X1   g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(G2096), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n631), .A2(new_n632), .A3(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT14), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n647), .A2(new_n654), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n655), .A2(new_n656), .A3(G14), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  OR3_X1    g238(.A1(new_n660), .A2(new_n658), .A3(new_n661), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n658), .A3(new_n661), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n639), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2100), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT81), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n674), .A2(new_n676), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n672), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n677), .A3(new_n672), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n678), .B1(new_n677), .B2(new_n672), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT86), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n693), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT33), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1976), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n693), .A2(G6), .ZN(new_n704));
  INV_X1    g279(.A(G305), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n693), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n698), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT85), .B(KEYINPUT34), .Z(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n478), .A2(G131), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(G95), .A2(G2105), .ZN(new_n718));
  INV_X1    g293(.A(G2104), .ZN(new_n719));
  INV_X1    g294(.A(G107), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G2105), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n474), .A2(G119), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n714), .B1(new_n724), .B2(new_n713), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT84), .Z(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n726), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n693), .A2(G24), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n594), .B(KEYINPUT78), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n693), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1986), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n711), .A2(new_n712), .A3(new_n729), .A4(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n713), .A2(G33), .ZN(new_n739));
  NAND2_X1  g314(.A1(G115), .A2(G2104), .ZN(new_n740));
  INV_X1    g315(.A(G127), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n463), .B2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n468), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n743), .B2(new_n742), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n748), .A2(new_n749), .B1(new_n478), .B2(G139), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n739), .B1(new_n751), .B2(new_n713), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT90), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(G2072), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT91), .ZN(new_n755));
  NAND2_X1  g330(.A1(G168), .A2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT94), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G16), .B2(G21), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT95), .B(G1966), .Z(new_n759));
  AND2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n693), .A2(G5), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G171), .B2(new_n693), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G1961), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT97), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n474), .A2(G129), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND3_X1  g342(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n478), .A2(G141), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n765), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(new_n713), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n771), .A2(KEYINPUT93), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(KEYINPUT93), .ZN(new_n773));
  OAI22_X1  g348(.A1(new_n772), .A2(new_n773), .B1(G29), .B2(G32), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n764), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n758), .A2(new_n759), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n760), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n753), .A2(G2072), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT92), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT31), .B(G11), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT96), .ZN(new_n784));
  INV_X1    g359(.A(G28), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n785), .B2(KEYINPUT30), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT30), .B2(new_n785), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n787), .C1(new_n638), .C2(new_n713), .ZN(new_n788));
  INV_X1    g363(.A(G1961), .ZN(new_n789));
  INV_X1    g364(.A(new_n762), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n713), .B1(KEYINPUT24), .B2(G34), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(KEYINPUT24), .B2(G34), .ZN(new_n793));
  INV_X1    g368(.A(G160), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2084), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n693), .A2(G19), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n546), .B2(new_n693), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1341), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n713), .A2(G35), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G162), .B2(new_n713), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT29), .B(G2090), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n791), .A2(new_n796), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G164), .A2(G29), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G27), .B2(G29), .ZN(new_n806));
  INV_X1    g381(.A(G2078), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n474), .A2(G128), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n478), .A2(G140), .ZN(new_n810));
  NOR2_X1   g385(.A1(G104), .A2(G2105), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G29), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n713), .A2(G26), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT28), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G2067), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n806), .A2(new_n807), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n808), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n693), .A2(G20), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT23), .Z(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(G299), .B2(G16), .ZN(new_n824));
  INV_X1    g399(.A(G1956), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n693), .A2(G4), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n614), .B2(new_n693), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT87), .B(G1348), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT88), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  NOR4_X1   g406(.A1(new_n804), .A2(new_n821), .A3(new_n826), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n755), .A2(new_n780), .A3(new_n782), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n738), .A2(new_n833), .ZN(G311));
  OR2_X1    g409(.A1(new_n738), .A2(new_n833), .ZN(G150));
  INV_X1    g410(.A(new_n546), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT99), .B(G93), .Z(new_n837));
  INV_X1    g412(.A(G55), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n513), .A2(new_n837), .B1(new_n838), .B2(new_n516), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  INV_X1    g416(.A(G80), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n603), .A2(new_n841), .B1(new_n842), .B2(new_n606), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI221_X1 g420(.A(KEYINPUT98), .B1(new_n842), .B2(new_n606), .C1(new_n603), .C2(new_n841), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(G651), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n836), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n546), .A2(new_n847), .A3(new_n840), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n614), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n856), .B2(new_n855), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT101), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n848), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(G145));
  XNOR2_X1  g437(.A(new_n499), .B(new_n813), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n770), .ZN(new_n864));
  INV_X1    g439(.A(new_n751), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n723), .B(KEYINPUT102), .ZN(new_n869));
  INV_X1    g444(.A(new_n628), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n723), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n628), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n474), .A2(G130), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n478), .A2(G142), .ZN(new_n876));
  OR2_X1    g451(.A1(G106), .A2(G2105), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n877), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n871), .A2(new_n874), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n871), .B2(new_n874), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n868), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n866), .B(new_n867), .C1(new_n881), .C2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n638), .B(G160), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G162), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n871), .A2(new_n874), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n879), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n871), .A2(new_n874), .A3(new_n880), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n866), .A3(new_n867), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n868), .A2(new_n883), .A3(new_n893), .ZN(new_n897));
  INV_X1    g472(.A(new_n888), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n889), .A2(new_n890), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n889), .A2(KEYINPUT104), .A3(new_n899), .A4(new_n890), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT40), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(G395));
  XNOR2_X1  g481(.A(new_n851), .B(new_n623), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n613), .A2(new_n564), .A3(new_n559), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n600), .A2(new_n601), .B1(G54), .B2(new_n529), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n561), .A2(new_n563), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n909), .B(new_n611), .C1(new_n910), .C2(new_n558), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(G299), .A2(new_n614), .A3(KEYINPUT105), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n907), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n917), .B(KEYINPUT106), .Z(new_n918));
  INV_X1    g493(.A(new_n907), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n908), .A2(new_n911), .A3(KEYINPUT107), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n613), .A2(new_n559), .A3(new_n922), .A4(new_n564), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n920), .B1(KEYINPUT41), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n918), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(G290), .A2(new_n705), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n732), .A2(G305), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G303), .B(G288), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(G303), .B(new_n700), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT42), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n926), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n926), .A2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n848), .A2(new_n617), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n939), .ZN(G331));
  NAND2_X1  g516(.A1(G168), .A2(G171), .ZN(new_n942));
  OAI21_X1  g517(.A(G301), .B1(new_n532), .B2(new_n533), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n851), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n942), .A2(new_n849), .A3(new_n850), .A4(new_n943), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n851), .A3(KEYINPUT108), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n951), .A3(new_n947), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n944), .A2(new_n851), .A3(KEYINPUT109), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n925), .A2(new_n950), .B1(new_n916), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n955), .B2(new_n934), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n916), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT41), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n921), .A2(new_n958), .A3(new_n923), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n913), .B2(new_n914), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n949), .B(new_n948), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n934), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n934), .A2(new_n957), .A3(new_n961), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n924), .A2(new_n958), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n958), .B2(new_n915), .ZN(new_n969));
  INV_X1    g544(.A(new_n954), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n948), .A2(new_n949), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n969), .A2(new_n970), .B1(new_n916), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n890), .B(new_n967), .C1(new_n972), .C2(new_n934), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n966), .B1(KEYINPUT43), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n964), .A2(new_n977), .A3(new_n890), .A4(new_n967), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n956), .A2(KEYINPUT110), .A3(new_n977), .A4(new_n964), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n975), .B1(new_n973), .B2(KEYINPUT43), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n982), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n976), .B1(new_n985), .B2(new_n986), .ZN(G397));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n499), .B2(new_n988), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n467), .A2(new_n472), .A3(G40), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n813), .B(G2067), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT112), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n770), .B(G1996), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n723), .A2(new_n728), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n724), .A2(new_n727), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(G290), .B(G1986), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n992), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1002));
  AND3_X1   g577(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT45), .B(new_n988), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n990), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n989), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1002), .B1(new_n1007), .B2(new_n807), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT124), .B(G2078), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1007), .A2(KEYINPUT53), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n988), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n499), .A2(KEYINPUT113), .A3(new_n988), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1013), .A2(KEYINPUT114), .A3(new_n1015), .A4(new_n1014), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1018), .A2(new_n990), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n1008), .B(new_n1010), .C1(new_n1021), .C2(new_n789), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1022), .A2(KEYINPUT125), .A3(G301), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT125), .B1(new_n1022), .B2(G301), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT45), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1026), .A2(new_n1006), .A3(new_n1027), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1008), .B(new_n1028), .C1(new_n1021), .C2(new_n789), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1025), .B1(new_n1029), .B2(G301), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1024), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT126), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n1022), .B2(G301), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1008), .B1(new_n1021), .B2(new_n789), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1010), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1029), .A2(G301), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1023), .A2(new_n1031), .B1(new_n1039), .B2(KEYINPUT54), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1014), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n990), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n825), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT56), .B(G2072), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1007), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G299), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n559), .A2(KEYINPUT57), .A3(new_n564), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1013), .A2(new_n990), .A3(new_n1015), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2067), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1021), .B2(new_n829), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1052), .B1(new_n1055), .B2(new_n613), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1043), .A2(new_n1050), .A3(new_n1045), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(KEYINPUT122), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1043), .A2(new_n1050), .A3(new_n1060), .A4(new_n1045), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(new_n1052), .A3(KEYINPUT61), .A4(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n613), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1064));
  INV_X1    g639(.A(new_n1057), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1050), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1068), .A2(KEYINPUT120), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT58), .B(G1341), .Z(new_n1070));
  AND2_X1   g645(.A1(new_n1053), .A2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1006), .A2(new_n989), .A3(G1996), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n546), .B(new_n1069), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1996), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1074), .A2(new_n1007), .B1(new_n1053), .B2(new_n1070), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1068), .A2(KEYINPUT120), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1075), .A2(new_n836), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1073), .B1(new_n1077), .B2(new_n1069), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1062), .A2(new_n1063), .A3(new_n1067), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1021), .A2(new_n829), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1054), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT60), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1083), .B(new_n1054), .C1(new_n1021), .C2(new_n829), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1082), .A2(new_n1084), .A3(new_n613), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1058), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT49), .ZN(new_n1087));
  INV_X1    g662(.A(G1981), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n575), .A2(new_n589), .A3(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n513), .A2(new_n572), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1088), .B1(new_n589), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1089), .B1(new_n1092), .B2(KEYINPUT117), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n501), .B1(new_n586), .B2(new_n587), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1094), .A2(new_n581), .A3(new_n1090), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1088), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1087), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1092), .A2(KEYINPUT117), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1095), .B2(new_n1088), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1099), .A2(KEYINPUT49), .A3(new_n1100), .A4(new_n1089), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1053), .A2(G8), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n700), .A2(G1976), .ZN(new_n1104));
  INV_X1    g679(.A(G1976), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT52), .B1(G288), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1053), .A2(G8), .A3(new_n1104), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1108), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT116), .B1(new_n1108), .B2(KEYINPUT52), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1103), .B(new_n1107), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT55), .ZN(new_n1112));
  AND3_X1   g687(.A1(G303), .A2(new_n1112), .A3(G8), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(G303), .B2(G8), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n697), .B1(new_n1006), .B2(new_n989), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1042), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1014), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1116), .B1(new_n1119), .B2(G2090), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1115), .B1(new_n1120), .B2(G8), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1111), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n990), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(G2090), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(KEYINPUT115), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1116), .B1(new_n1125), .B2(KEYINPUT115), .ZN(new_n1127));
  OAI211_X1 g702(.A(G8), .B(new_n1115), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1123), .A2(G2084), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(G1966), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n1026), .B2(new_n1006), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(G168), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1130), .B1(new_n1135), .B2(G8), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(G286), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT51), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1135), .A2(G8), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1129), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1086), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1040), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1137), .A2(G8), .A3(G168), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1122), .A2(new_n1128), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT63), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1111), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(G8), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1115), .A2(KEYINPUT119), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI221_X1 g729(.A(G8), .B1(KEYINPUT119), .B2(new_n1115), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1149), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1029), .A2(G301), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1122), .A2(new_n1158), .A3(new_n1128), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1130), .B1(new_n1137), .B2(G286), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1135), .A2(G8), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT62), .B1(new_n1162), .B2(new_n1136), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1136), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1164), .B(new_n1165), .C1(new_n1161), .C2(new_n1160), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1159), .A2(new_n1163), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1128), .A2(new_n1111), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1103), .A2(new_n1105), .A3(new_n700), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1089), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1168), .B1(new_n1102), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1157), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1001), .B1(new_n1144), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n996), .A2(new_n727), .A3(new_n724), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n813), .A2(G2067), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n991), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n999), .A2(new_n992), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n992), .A2(new_n686), .A3(new_n732), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT48), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1176), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT47), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n992), .B1(new_n994), .B2(new_n770), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n992), .A2(KEYINPUT46), .A3(new_n1074), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT46), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1184), .B1(new_n991), .B2(G1996), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT127), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1180), .B1(new_n1181), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1188), .B1(new_n1181), .B2(new_n1187), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1173), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g765(.A1(new_n902), .A2(new_n903), .ZN(new_n1192));
  NOR4_X1   g766(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n1192), .A2(new_n974), .A3(new_n1193), .ZN(G225));
  INV_X1    g768(.A(G225), .ZN(G308));
endmodule


