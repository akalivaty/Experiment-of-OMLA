

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811;

  BUF_X1 U376 ( .A(n700), .Z(n355) );
  INV_X1 U377 ( .A(KEYINPUT82), .ZN(n357) );
  AND2_X1 U378 ( .A1(n453), .A2(n454), .ZN(n424) );
  OR2_X1 U379 ( .A1(n634), .A2(n675), .ZN(n482) );
  AND2_X1 U380 ( .A1(n425), .A2(n738), .ZN(n633) );
  AND2_X1 U381 ( .A1(n471), .A2(n522), .ZN(n521) );
  XNOR2_X1 U382 ( .A(n488), .B(KEYINPUT19), .ZN(n664) );
  XNOR2_X1 U383 ( .A(n401), .B(n566), .ZN(n663) );
  XNOR2_X1 U384 ( .A(n593), .B(n483), .ZN(n747) );
  XNOR2_X1 U385 ( .A(n430), .B(n530), .ZN(n796) );
  INV_X1 U386 ( .A(KEYINPUT75), .ZN(n428) );
  INV_X1 U387 ( .A(G116), .ZN(n413) );
  AND2_X2 U388 ( .A1(n790), .A2(n697), .ZN(n494) );
  NOR2_X2 U389 ( .A1(n727), .A2(KEYINPUT73), .ZN(n465) );
  XNOR2_X2 U390 ( .A(n356), .B(n469), .ZN(n808) );
  NAND2_X2 U391 ( .A1(n422), .A2(n420), .ZN(n356) );
  XNOR2_X1 U392 ( .A(n698), .B(n357), .ZN(n359) );
  NOR2_X2 U393 ( .A1(n635), .A2(n644), .ZN(n636) );
  NAND2_X1 U394 ( .A1(n646), .A2(n630), .ZN(n631) );
  XNOR2_X2 U395 ( .A(n487), .B(n370), .ZN(n646) );
  NAND2_X1 U396 ( .A1(n358), .A2(n443), .ZN(n612) );
  AND2_X1 U397 ( .A1(n444), .A2(n683), .ZN(n358) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n582) );
  XOR2_X1 U399 ( .A(G137), .B(G140), .Z(n571) );
  INV_X1 U400 ( .A(G953), .ZN(n798) );
  AND2_X2 U401 ( .A1(n688), .A2(n514), .ZN(n513) );
  XNOR2_X2 U402 ( .A(n429), .B(KEYINPUT38), .ZN(n755) );
  INV_X2 U403 ( .A(G104), .ZN(n492) );
  INV_X2 U404 ( .A(G143), .ZN(n508) );
  XNOR2_X2 U405 ( .A(n417), .B(n418), .ZN(n665) );
  NAND2_X2 U406 ( .A1(n403), .A2(n535), .ZN(n698) );
  XNOR2_X2 U407 ( .A(n404), .B(n501), .ZN(n403) );
  XNOR2_X2 U408 ( .A(n796), .B(G146), .ZN(n414) );
  XNOR2_X1 U409 ( .A(n623), .B(KEYINPUT102), .ZN(n651) );
  INV_X1 U410 ( .A(KEYINPUT23), .ZN(n526) );
  NAND2_X1 U411 ( .A1(n516), .A2(n513), .ZN(n404) );
  AND2_X1 U412 ( .A1(n673), .A2(n461), .ZN(n460) );
  NAND2_X1 U413 ( .A1(n687), .A2(n719), .ZN(n449) );
  NAND2_X1 U414 ( .A1(n406), .A2(n405), .ZN(n768) );
  XNOR2_X1 U415 ( .A(n482), .B(KEYINPUT78), .ZN(n635) );
  XNOR2_X1 U416 ( .A(n447), .B(n476), .ZN(n443) );
  BUF_X1 U417 ( .A(n616), .Z(n429) );
  XNOR2_X1 U418 ( .A(n509), .B(n533), .ZN(n616) );
  NAND2_X1 U419 ( .A1(n705), .A2(n695), .ZN(n509) );
  XNOR2_X1 U420 ( .A(n475), .B(n577), .ZN(n742) );
  NOR2_X1 U421 ( .A1(n776), .A2(G902), .ZN(n401) );
  XNOR2_X1 U422 ( .A(n549), .B(n364), .ZN(n506) );
  XNOR2_X1 U423 ( .A(n526), .B(G110), .ZN(n574) );
  XNOR2_X1 U424 ( .A(n594), .B(KEYINPUT10), .ZN(n570) );
  NAND2_X1 U425 ( .A1(n503), .A2(n772), .ZN(n360) );
  BUF_X1 U426 ( .A(n769), .Z(n361) );
  NAND2_X1 U427 ( .A1(n503), .A2(n772), .ZN(n502) );
  XNOR2_X1 U428 ( .A(n637), .B(KEYINPUT33), .ZN(n769) );
  AND2_X1 U429 ( .A1(n738), .A2(n737), .ZN(n415) );
  NOR2_X1 U430 ( .A1(n742), .A2(n741), .ZN(n737) );
  XNOR2_X1 U431 ( .A(G902), .B(KEYINPUT15), .ZN(n695) );
  OR2_X1 U432 ( .A1(n710), .A2(G902), .ZN(n475) );
  INV_X1 U433 ( .A(G472), .ZN(n483) );
  INV_X1 U434 ( .A(KEYINPUT76), .ZN(n476) );
  NAND2_X1 U435 ( .A1(n427), .A2(n416), .ZN(n447) );
  INV_X1 U436 ( .A(n660), .ZN(n416) );
  INV_X1 U437 ( .A(KEYINPUT74), .ZN(n418) );
  AND2_X1 U438 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U439 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n563) );
  INV_X1 U440 ( .A(KEYINPUT16), .ZN(n491) );
  XNOR2_X1 U441 ( .A(n604), .B(n459), .ZN(n498) );
  NAND2_X1 U442 ( .A1(n683), .A2(n409), .ZN(n408) );
  NOR2_X1 U443 ( .A1(n412), .A2(n410), .ZN(n409) );
  NAND2_X1 U444 ( .A1(n677), .A2(n411), .ZN(n410) );
  INV_X1 U445 ( .A(KEYINPUT86), .ZN(n438) );
  XNOR2_X1 U446 ( .A(n663), .B(n532), .ZN(n738) );
  XNOR2_X1 U447 ( .A(n632), .B(KEYINPUT66), .ZN(n532) );
  XOR2_X1 U448 ( .A(G134), .B(G122), .Z(n549) );
  NAND2_X1 U449 ( .A1(n369), .A2(n484), .ZN(n772) );
  INV_X1 U450 ( .A(n698), .ZN(n484) );
  AND2_X1 U451 ( .A1(n675), .A2(n479), .ZN(n678) );
  XNOR2_X1 U452 ( .A(n631), .B(KEYINPUT22), .ZN(n644) );
  XNOR2_X1 U453 ( .A(n446), .B(n445), .ZN(n444) );
  NOR2_X1 U454 ( .A1(n452), .A2(n490), .ZN(n489) );
  INV_X1 U455 ( .A(n425), .ZN(n490) );
  AND2_X1 U456 ( .A1(n580), .A2(n737), .ZN(n427) );
  BUF_X1 U457 ( .A(n742), .Z(n425) );
  XNOR2_X1 U458 ( .A(n747), .B(n486), .ZN(n675) );
  INV_X1 U459 ( .A(KEYINPUT6), .ZN(n486) );
  NAND2_X1 U460 ( .A1(n395), .A2(G472), .ZN(n383) );
  INV_X1 U461 ( .A(n709), .ZN(n388) );
  XNOR2_X1 U462 ( .A(n705), .B(n708), .ZN(n709) );
  NAND2_X1 U463 ( .A1(n682), .A2(KEYINPUT72), .ZN(n451) );
  XNOR2_X1 U464 ( .A(n448), .B(n371), .ZN(n688) );
  NAND2_X1 U465 ( .A1(n436), .A2(n450), .ZN(n435) );
  NAND2_X1 U466 ( .A1(n682), .A2(n674), .ZN(n450) );
  INV_X1 U467 ( .A(KEYINPUT103), .ZN(n510) );
  INV_X1 U468 ( .A(n662), .ZN(n523) );
  INV_X1 U469 ( .A(KEYINPUT18), .ZN(n507) );
  XNOR2_X1 U470 ( .A(n595), .B(KEYINPUT17), .ZN(n474) );
  INV_X1 U471 ( .A(KEYINPUT77), .ZN(n595) );
  OR2_X1 U472 ( .A1(G902), .A2(G237), .ZN(n611) );
  AND2_X1 U473 ( .A1(n747), .A2(n662), .ZN(n519) );
  XNOR2_X1 U474 ( .A(KEYINPUT13), .B(G475), .ZN(n545) );
  XNOR2_X1 U475 ( .A(KEYINPUT69), .B(G134), .ZN(n531) );
  NOR2_X1 U476 ( .A1(n396), .A2(n372), .ZN(n527) );
  XNOR2_X1 U477 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U478 ( .A(G107), .B(G101), .ZN(n558) );
  INV_X1 U479 ( .A(G104), .ZN(n557) );
  XNOR2_X1 U480 ( .A(G116), .B(G137), .ZN(n586) );
  INV_X1 U481 ( .A(KEYINPUT95), .ZN(n585) );
  XOR2_X1 U482 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n584) );
  XNOR2_X1 U483 ( .A(n468), .B(n602), .ZN(n783) );
  XNOR2_X1 U484 ( .A(n600), .B(n491), .ZN(n601) );
  XNOR2_X1 U485 ( .A(n498), .B(n570), .ZN(n499) );
  NAND2_X1 U486 ( .A1(n415), .A2(n675), .ZN(n637) );
  NAND2_X1 U487 ( .A1(G237), .A2(G234), .ZN(n554) );
  NAND2_X1 U488 ( .A1(n362), .A2(KEYINPUT41), .ZN(n405) );
  AND2_X1 U489 ( .A1(n408), .A2(n407), .ZN(n406) );
  XNOR2_X1 U490 ( .A(n612), .B(KEYINPUT39), .ZN(n687) );
  XNOR2_X1 U491 ( .A(n679), .B(n438), .ZN(n437) );
  NOR2_X1 U492 ( .A1(n689), .A2(n440), .ZN(n439) );
  INV_X1 U493 ( .A(KEYINPUT34), .ZN(n638) );
  XNOR2_X1 U494 ( .A(n473), .B(n472), .ZN(n685) );
  INV_X1 U495 ( .A(KEYINPUT108), .ZN(n472) );
  NAND2_X1 U496 ( .A1(n524), .A2(n580), .ZN(n473) );
  AND2_X1 U497 ( .A1(n572), .A2(G217), .ZN(n504) );
  NAND2_X1 U498 ( .A1(n359), .A2(n496), .ZN(n495) );
  INV_X1 U499 ( .A(n681), .ZN(n515) );
  AND2_X1 U500 ( .A1(n443), .A2(n444), .ZN(n668) );
  INV_X1 U501 ( .A(KEYINPUT106), .ZN(n469) );
  AND2_X1 U502 ( .A1(n489), .A2(n421), .ZN(n420) );
  AND2_X1 U503 ( .A1(n646), .A2(n427), .ZN(n621) );
  NOR2_X1 U504 ( .A1(n675), .A2(n477), .ZN(n419) );
  NAND2_X1 U505 ( .A1(n382), .A2(n386), .ZN(n381) );
  XNOR2_X1 U506 ( .A(n383), .B(n373), .ZN(n382) );
  INV_X1 U507 ( .A(KEYINPUT60), .ZN(n377) );
  XNOR2_X1 U508 ( .A(n380), .B(n363), .ZN(n379) );
  INV_X1 U509 ( .A(KEYINPUT56), .ZN(n384) );
  NAND2_X1 U510 ( .A1(n387), .A2(n386), .ZN(n385) );
  XNOR2_X1 U511 ( .A(n389), .B(n388), .ZN(n387) );
  XNOR2_X1 U512 ( .A(n390), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U513 ( .A1(n391), .A2(G953), .ZN(n390) );
  XNOR2_X1 U514 ( .A(n392), .B(KEYINPUT118), .ZN(n391) );
  OR2_X1 U515 ( .A1(n774), .A2(n775), .ZN(n392) );
  INV_X1 U516 ( .A(n756), .ZN(n677) );
  OR2_X1 U517 ( .A1(n412), .A2(n756), .ZN(n362) );
  XNOR2_X1 U518 ( .A(KEYINPUT59), .B(n704), .ZN(n363) );
  XOR2_X1 U519 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n364) );
  NOR2_X1 U520 ( .A1(n478), .A2(n684), .ZN(n365) );
  INV_X1 U521 ( .A(n525), .ZN(n452) );
  XNOR2_X1 U522 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n366) );
  AND2_X1 U523 ( .A1(n495), .A2(n697), .ZN(n367) );
  AND2_X1 U524 ( .A1(n683), .A2(n677), .ZN(n368) );
  XNOR2_X1 U525 ( .A(n565), .B(G469), .ZN(n566) );
  NOR2_X1 U526 ( .A1(n790), .A2(n697), .ZN(n369) );
  INV_X1 U527 ( .A(G902), .ZN(n550) );
  XOR2_X1 U528 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n370) );
  XOR2_X1 U529 ( .A(KEYINPUT84), .B(KEYINPUT46), .Z(n371) );
  INV_X1 U530 ( .A(KEYINPUT41), .ZN(n411) );
  AND2_X1 U531 ( .A1(n650), .A2(n684), .ZN(n719) );
  INV_X1 U532 ( .A(n719), .ZN(n480) );
  OR2_X1 U533 ( .A1(n695), .A2(KEYINPUT2), .ZN(n372) );
  XOR2_X1 U534 ( .A(n355), .B(n699), .Z(n373) );
  OR2_X1 U535 ( .A1(n695), .A2(KEYINPUT81), .ZN(n374) );
  XNOR2_X1 U536 ( .A(n499), .B(n543), .ZN(n500) );
  AND2_X1 U537 ( .A1(KEYINPUT85), .A2(KEYINPUT44), .ZN(n375) );
  XNOR2_X1 U538 ( .A(n703), .B(n702), .ZN(n782) );
  INV_X1 U539 ( .A(n782), .ZN(n386) );
  NAND2_X1 U540 ( .A1(n376), .A2(G478), .ZN(n715) );
  NAND2_X1 U541 ( .A1(n376), .A2(G210), .ZN(n389) );
  XNOR2_X2 U542 ( .A(n502), .B(KEYINPUT65), .ZN(n376) );
  XNOR2_X1 U543 ( .A(n378), .B(n377), .ZN(G60) );
  NAND2_X1 U544 ( .A1(n379), .A2(n386), .ZN(n378) );
  NAND2_X1 U545 ( .A1(n395), .A2(G475), .ZN(n380) );
  XNOR2_X1 U546 ( .A(n381), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U547 ( .A(n385), .B(n384), .ZN(G51) );
  XNOR2_X2 U548 ( .A(n360), .B(KEYINPUT65), .ZN(n395) );
  BUF_X1 U549 ( .A(n753), .Z(n393) );
  XNOR2_X1 U550 ( .A(n698), .B(KEYINPUT82), .ZN(n394) );
  XNOR2_X1 U551 ( .A(n658), .B(n657), .ZN(n396) );
  XNOR2_X1 U552 ( .A(n658), .B(n657), .ZN(n790) );
  INV_X1 U553 ( .A(n429), .ZN(n440) );
  NOR2_X1 U554 ( .A1(n458), .A2(KEYINPUT85), .ZN(n457) );
  NAND2_X1 U555 ( .A1(n655), .A2(n654), .ZN(n458) );
  BUF_X1 U556 ( .A(n738), .Z(n477) );
  NAND2_X1 U557 ( .A1(n462), .A2(n460), .ZN(n432) );
  NAND2_X1 U558 ( .A1(n512), .A2(n506), .ZN(n399) );
  NAND2_X1 U559 ( .A1(n397), .A2(n398), .ZN(n400) );
  NAND2_X1 U560 ( .A1(n399), .A2(n400), .ZN(n505) );
  INV_X1 U561 ( .A(n512), .ZN(n397) );
  INV_X1 U562 ( .A(n506), .ZN(n398) );
  XNOR2_X2 U563 ( .A(n505), .B(n504), .ZN(n714) );
  AND2_X2 U564 ( .A1(n462), .A2(n460), .ZN(n402) );
  XNOR2_X1 U565 ( .A(n551), .B(G478), .ZN(n627) );
  NAND2_X1 U566 ( .A1(n402), .A2(n435), .ZN(n423) );
  NAND2_X1 U567 ( .A1(n810), .A2(n811), .ZN(n448) );
  NAND2_X1 U568 ( .A1(n755), .A2(KEYINPUT41), .ZN(n407) );
  INV_X1 U569 ( .A(n365), .ZN(n412) );
  XNOR2_X2 U570 ( .A(n413), .B(G107), .ZN(n603) );
  XNOR2_X1 U571 ( .A(n414), .B(n564), .ZN(n776) );
  XNOR2_X1 U572 ( .A(n414), .B(n592), .ZN(n700) );
  AND2_X1 U573 ( .A1(n415), .A2(n452), .ZN(n749) );
  NOR2_X2 U574 ( .A1(n659), .A2(KEYINPUT47), .ZN(n417) );
  XNOR2_X2 U575 ( .A(n753), .B(KEYINPUT80), .ZN(n659) );
  XNOR2_X2 U576 ( .A(n511), .B(n510), .ZN(n753) );
  NAND2_X1 U577 ( .A1(n422), .A2(n419), .ZN(n653) );
  INV_X1 U578 ( .A(n477), .ZN(n421) );
  INV_X1 U579 ( .A(n644), .ZN(n422) );
  NAND2_X1 U580 ( .A1(n423), .A2(n431), .ZN(n516) );
  XOR2_X2 U581 ( .A(KEYINPUT32), .B(n636), .Z(n809) );
  INV_X1 U582 ( .A(n663), .ZN(n580) );
  NAND2_X1 U583 ( .A1(n424), .A2(n455), .ZN(n485) );
  NAND2_X1 U584 ( .A1(n457), .A2(n456), .ZN(n455) );
  NAND2_X1 U585 ( .A1(n426), .A2(n696), .ZN(n503) );
  NAND2_X1 U586 ( .A1(n493), .A2(n497), .ZN(n426) );
  XNOR2_X2 U587 ( .A(n428), .B(G110), .ZN(n600) );
  XNOR2_X2 U588 ( .A(n441), .B(n563), .ZN(n430) );
  XNOR2_X1 U589 ( .A(n430), .B(n507), .ZN(n598) );
  NAND2_X1 U590 ( .A1(n433), .A2(n432), .ZN(n431) );
  NAND2_X1 U591 ( .A1(n434), .A2(n451), .ZN(n433) );
  NAND2_X1 U592 ( .A1(n517), .A2(n674), .ZN(n434) );
  NAND2_X1 U593 ( .A1(n517), .A2(KEYINPUT72), .ZN(n436) );
  XNOR2_X1 U594 ( .A(n439), .B(n437), .ZN(n680) );
  XNOR2_X1 U595 ( .A(n603), .B(n441), .ZN(n512) );
  XNOR2_X2 U596 ( .A(n508), .B(G128), .ZN(n441) );
  INV_X1 U597 ( .A(KEYINPUT30), .ZN(n445) );
  NAND2_X1 U598 ( .A1(n747), .A2(n677), .ZN(n446) );
  XNOR2_X2 U599 ( .A(n449), .B(KEYINPUT40), .ZN(n810) );
  NAND2_X1 U600 ( .A1(n656), .A2(n375), .ZN(n453) );
  NAND2_X1 U601 ( .A1(n458), .A2(KEYINPUT85), .ZN(n454) );
  NAND2_X1 U602 ( .A1(n656), .A2(KEYINPUT44), .ZN(n456) );
  NAND2_X1 U603 ( .A1(n645), .A2(n809), .ZN(n656) );
  XNOR2_X1 U604 ( .A(n459), .B(n531), .ZN(n530) );
  XNOR2_X2 U605 ( .A(KEYINPUT68), .B(G131), .ZN(n459) );
  NAND2_X1 U606 ( .A1(n727), .A2(KEYINPUT73), .ZN(n461) );
  AND2_X2 U607 ( .A1(n464), .A2(n463), .ZN(n462) );
  NAND2_X1 U608 ( .A1(n665), .A2(KEYINPUT73), .ZN(n463) );
  NAND2_X1 U609 ( .A1(n466), .A2(n465), .ZN(n464) );
  INV_X1 U610 ( .A(n665), .ZN(n466) );
  NAND2_X1 U611 ( .A1(n467), .A2(n652), .ZN(n655) );
  XNOR2_X1 U612 ( .A(n649), .B(KEYINPUT98), .ZN(n467) );
  NAND2_X1 U613 ( .A1(n606), .A2(n607), .ZN(n610) );
  XNOR2_X1 U614 ( .A(n605), .B(n601), .ZN(n468) );
  NAND2_X1 U615 ( .A1(n525), .A2(n523), .ZN(n471) );
  XNOR2_X2 U616 ( .A(n492), .B(G122), .ZN(n604) );
  NAND2_X1 U617 ( .A1(n720), .A2(n731), .ZN(n649) );
  NAND2_X1 U618 ( .A1(n622), .A2(n525), .ZN(n720) );
  XNOR2_X1 U619 ( .A(n598), .B(n599), .ZN(n607) );
  XNOR2_X1 U620 ( .A(n594), .B(n474), .ZN(n597) );
  NOR2_X1 U621 ( .A1(n700), .A2(G902), .ZN(n593) );
  BUF_X1 U622 ( .A(n627), .Z(n478) );
  NAND2_X1 U623 ( .A1(n680), .A2(n477), .ZN(n681) );
  NOR2_X1 U624 ( .A1(n676), .A2(n480), .ZN(n479) );
  NAND2_X1 U625 ( .A1(n714), .A2(n550), .ZN(n551) );
  XNOR2_X2 U626 ( .A(n481), .B(KEYINPUT101), .ZN(n623) );
  NAND2_X1 U627 ( .A1(n627), .A2(n640), .ZN(n481) );
  XNOR2_X1 U628 ( .A(n529), .B(n795), .ZN(n710) );
  NAND2_X1 U629 ( .A1(n769), .A2(n646), .ZN(n639) );
  NAND2_X1 U630 ( .A1(n394), .A2(n697), .ZN(n497) );
  NAND2_X1 U631 ( .A1(n485), .A2(n536), .ZN(n658) );
  NAND2_X1 U632 ( .A1(n664), .A2(n620), .ZN(n487) );
  NAND2_X1 U633 ( .A1(n616), .A2(n677), .ZN(n488) );
  NOR2_X1 U634 ( .A1(n494), .A2(n374), .ZN(n493) );
  INV_X1 U635 ( .A(n396), .ZN(n496) );
  NAND2_X1 U636 ( .A1(n500), .A2(n550), .ZN(n546) );
  INV_X1 U637 ( .A(n500), .ZN(n704) );
  INV_X1 U638 ( .A(KEYINPUT48), .ZN(n501) );
  INV_X1 U639 ( .A(n755), .ZN(n683) );
  XNOR2_X1 U640 ( .A(n597), .B(n596), .ZN(n599) );
  XNOR2_X2 U641 ( .A(G146), .B(G125), .ZN(n594) );
  NOR2_X2 U642 ( .A1(n651), .A2(n719), .ZN(n511) );
  NAND2_X1 U643 ( .A1(n515), .A2(KEYINPUT70), .ZN(n514) );
  NAND2_X1 U644 ( .A1(n681), .A2(n682), .ZN(n517) );
  NAND2_X1 U645 ( .A1(n521), .A2(n518), .ZN(n524) );
  NAND2_X1 U646 ( .A1(n520), .A2(n519), .ZN(n518) );
  INV_X1 U647 ( .A(n676), .ZN(n520) );
  NAND2_X1 U648 ( .A1(n676), .A2(n523), .ZN(n522) );
  INV_X1 U649 ( .A(n747), .ZN(n525) );
  NAND2_X1 U650 ( .A1(n359), .A2(n527), .ZN(n694) );
  XNOR2_X1 U651 ( .A(n528), .B(n576), .ZN(n529) );
  XNOR2_X1 U652 ( .A(n575), .B(n366), .ZN(n528) );
  AND2_X1 U653 ( .A1(G210), .A2(n611), .ZN(n533) );
  XOR2_X1 U654 ( .A(n545), .B(n544), .Z(n534) );
  NOR2_X1 U655 ( .A1(n736), .A2(n693), .ZN(n535) );
  OR2_X1 U656 ( .A1(n656), .A2(KEYINPUT44), .ZN(n536) );
  INV_X1 U657 ( .A(KEYINPUT72), .ZN(n674) );
  XNOR2_X1 U658 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U659 ( .A(n588), .B(n587), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n560), .B(n559), .ZN(n562) );
  XNOR2_X1 U661 ( .A(n591), .B(n602), .ZN(n592) );
  XNOR2_X1 U662 ( .A(G134), .B(KEYINPUT114), .ZN(n613) );
  NAND2_X1 U663 ( .A1(n582), .A2(G214), .ZN(n538) );
  XNOR2_X1 U664 ( .A(G143), .B(G140), .ZN(n537) );
  XNOR2_X1 U665 ( .A(n538), .B(n537), .ZN(n542) );
  XNOR2_X1 U666 ( .A(G113), .B(KEYINPUT12), .ZN(n540) );
  XNOR2_X1 U667 ( .A(KEYINPUT99), .B(KEYINPUT11), .ZN(n539) );
  XNOR2_X1 U668 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U669 ( .A(n542), .B(n541), .ZN(n543) );
  INV_X1 U670 ( .A(KEYINPUT100), .ZN(n544) );
  XNOR2_X2 U671 ( .A(n546), .B(n534), .ZN(n640) );
  NAND2_X1 U672 ( .A1(n798), .A2(G234), .ZN(n548) );
  XNOR2_X1 U673 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n547) );
  XNOR2_X1 U674 ( .A(n548), .B(n547), .ZN(n572) );
  NOR2_X1 U675 ( .A1(G900), .A2(n798), .ZN(n552) );
  NAND2_X1 U676 ( .A1(n552), .A2(G902), .ZN(n553) );
  NAND2_X1 U677 ( .A1(G952), .A2(n798), .ZN(n617) );
  NAND2_X1 U678 ( .A1(n553), .A2(n617), .ZN(n556) );
  XOR2_X1 U679 ( .A(n554), .B(KEYINPUT14), .Z(n766) );
  INV_X1 U680 ( .A(n766), .ZN(n555) );
  NAND2_X1 U681 ( .A1(n556), .A2(n555), .ZN(n660) );
  XOR2_X1 U682 ( .A(n571), .B(n600), .Z(n560) );
  NAND2_X1 U683 ( .A1(G227), .A2(n798), .ZN(n561) );
  XNOR2_X1 U684 ( .A(n562), .B(n561), .ZN(n564) );
  INV_X1 U685 ( .A(KEYINPUT71), .ZN(n565) );
  XOR2_X1 U686 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n569) );
  NAND2_X1 U687 ( .A1(n695), .A2(G234), .ZN(n567) );
  XNOR2_X1 U688 ( .A(n567), .B(KEYINPUT20), .ZN(n578) );
  NAND2_X1 U689 ( .A1(n578), .A2(G217), .ZN(n568) );
  XNOR2_X1 U690 ( .A(n569), .B(n568), .ZN(n577) );
  XNOR2_X1 U691 ( .A(n570), .B(n571), .ZN(n795) );
  NAND2_X1 U692 ( .A1(G221), .A2(n572), .ZN(n576) );
  XNOR2_X1 U693 ( .A(G128), .B(G119), .ZN(n573) );
  XNOR2_X1 U694 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U695 ( .A1(G221), .A2(n578), .ZN(n579) );
  XNOR2_X1 U696 ( .A(KEYINPUT21), .B(n579), .ZN(n741) );
  NAND2_X1 U697 ( .A1(n611), .A2(G214), .ZN(n581) );
  XNOR2_X1 U698 ( .A(KEYINPUT91), .B(n581), .ZN(n756) );
  NAND2_X1 U699 ( .A1(n582), .A2(G210), .ZN(n583) );
  XNOR2_X1 U700 ( .A(n584), .B(n583), .ZN(n588) );
  XOR2_X1 U701 ( .A(G101), .B(G113), .Z(n590) );
  XNOR2_X1 U702 ( .A(KEYINPUT3), .B(G119), .ZN(n589) );
  XNOR2_X1 U703 ( .A(n590), .B(n589), .ZN(n602) );
  NAND2_X1 U704 ( .A1(G224), .A2(n798), .ZN(n596) );
  XNOR2_X1 U705 ( .A(n604), .B(n603), .ZN(n605) );
  INV_X1 U706 ( .A(n783), .ZN(n606) );
  INV_X1 U707 ( .A(n607), .ZN(n608) );
  NAND2_X1 U708 ( .A1(n608), .A2(n783), .ZN(n609) );
  NAND2_X1 U709 ( .A1(n610), .A2(n609), .ZN(n705) );
  AND2_X1 U710 ( .A1(n651), .A2(n687), .ZN(n693) );
  XOR2_X1 U711 ( .A(n613), .B(n693), .Z(G36) );
  XOR2_X1 U712 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n615) );
  XNOR2_X1 U713 ( .A(G107), .B(KEYINPUT110), .ZN(n614) );
  XNOR2_X1 U714 ( .A(n615), .B(n614), .ZN(n625) );
  NOR2_X1 U715 ( .A1(G898), .A2(n798), .ZN(n784) );
  NAND2_X1 U716 ( .A1(n784), .A2(G902), .ZN(n618) );
  AND2_X1 U717 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U718 ( .A1(n619), .A2(n766), .ZN(n620) );
  XNOR2_X1 U719 ( .A(n621), .B(KEYINPUT94), .ZN(n622) );
  INV_X1 U720 ( .A(n623), .ZN(n730) );
  NOR2_X1 U721 ( .A1(n720), .A2(n730), .ZN(n624) );
  XOR2_X1 U722 ( .A(n625), .B(n624), .Z(G9) );
  INV_X1 U723 ( .A(n741), .ZN(n626) );
  NAND2_X1 U724 ( .A1(n640), .A2(n626), .ZN(n628) );
  NOR2_X1 U725 ( .A1(n628), .A2(n478), .ZN(n629) );
  XNOR2_X1 U726 ( .A(KEYINPUT104), .B(n629), .ZN(n630) );
  INV_X1 U727 ( .A(KEYINPUT1), .ZN(n632) );
  XNOR2_X1 U728 ( .A(n633), .B(KEYINPUT105), .ZN(n634) );
  XNOR2_X1 U729 ( .A(n639), .B(n638), .ZN(n641) );
  INV_X1 U730 ( .A(n640), .ZN(n684) );
  AND2_X1 U731 ( .A1(n478), .A2(n684), .ZN(n666) );
  NAND2_X1 U732 ( .A1(n641), .A2(n666), .ZN(n643) );
  XOR2_X1 U733 ( .A(KEYINPUT83), .B(KEYINPUT35), .Z(n642) );
  XNOR2_X1 U734 ( .A(n643), .B(n642), .ZN(n807) );
  NOR2_X1 U735 ( .A1(n807), .A2(n808), .ZN(n645) );
  XNOR2_X1 U736 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n648) );
  NAND2_X1 U737 ( .A1(n646), .A2(n749), .ZN(n647) );
  XNOR2_X1 U738 ( .A(n648), .B(n647), .ZN(n731) );
  INV_X1 U739 ( .A(n478), .ZN(n650) );
  INV_X1 U740 ( .A(n659), .ZN(n652) );
  NOR2_X1 U741 ( .A1(n425), .A2(n653), .ZN(n718) );
  INV_X1 U742 ( .A(n718), .ZN(n654) );
  INV_X1 U743 ( .A(KEYINPUT45), .ZN(n657) );
  XOR2_X1 U744 ( .A(KEYINPUT28), .B(KEYINPUT107), .Z(n662) );
  NOR2_X1 U745 ( .A1(n741), .A2(n660), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n742), .A2(n661), .ZN(n676) );
  NAND2_X1 U747 ( .A1(n664), .A2(n685), .ZN(n727) );
  NAND2_X1 U748 ( .A1(n727), .A2(KEYINPUT47), .ZN(n672) );
  AND2_X1 U749 ( .A1(n429), .A2(n666), .ZN(n667) );
  NAND2_X1 U750 ( .A1(n668), .A2(n667), .ZN(n726) );
  AND2_X1 U751 ( .A1(n753), .A2(KEYINPUT47), .ZN(n669) );
  XNOR2_X1 U752 ( .A(n669), .B(KEYINPUT79), .ZN(n670) );
  AND2_X1 U753 ( .A1(n726), .A2(n670), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n689) );
  INV_X1 U755 ( .A(KEYINPUT36), .ZN(n679) );
  INV_X1 U756 ( .A(KEYINPUT70), .ZN(n682) );
  NAND2_X1 U757 ( .A1(n685), .A2(n768), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n686), .B(KEYINPUT42), .ZN(n811) );
  NOR2_X1 U759 ( .A1(n689), .A2(n477), .ZN(n691) );
  INV_X1 U760 ( .A(KEYINPUT43), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n691), .B(n690), .ZN(n692) );
  AND2_X1 U762 ( .A1(n692), .A2(n440), .ZN(n736) );
  NAND2_X1 U763 ( .A1(n694), .A2(KEYINPUT81), .ZN(n696) );
  INV_X1 U764 ( .A(KEYINPUT2), .ZN(n697) );
  XOR2_X1 U765 ( .A(KEYINPUT89), .B(KEYINPUT62), .Z(n699) );
  INV_X1 U766 ( .A(G952), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n701), .A2(G953), .ZN(n703) );
  INV_X1 U768 ( .A(KEYINPUT90), .ZN(n702) );
  XNOR2_X1 U769 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n707) );
  XNOR2_X1 U770 ( .A(KEYINPUT55), .B(KEYINPUT87), .ZN(n706) );
  XNOR2_X1 U771 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n376), .A2(G217), .ZN(n712) );
  XNOR2_X1 U773 ( .A(n710), .B(KEYINPUT122), .ZN(n711) );
  XNOR2_X1 U774 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U775 ( .A1(n713), .A2(n782), .ZN(G66) );
  XNOR2_X1 U776 ( .A(n714), .B(n715), .ZN(n716) );
  NAND2_X1 U777 ( .A1(n716), .A2(n386), .ZN(n717) );
  XNOR2_X1 U778 ( .A(n717), .B(KEYINPUT121), .ZN(G63) );
  XOR2_X1 U779 ( .A(G101), .B(n718), .Z(G3) );
  NOR2_X1 U780 ( .A1(n720), .A2(n480), .ZN(n722) );
  XNOR2_X1 U781 ( .A(G104), .B(KEYINPUT109), .ZN(n721) );
  XNOR2_X1 U782 ( .A(n722), .B(n721), .ZN(G6) );
  NOR2_X1 U783 ( .A1(n727), .A2(n730), .ZN(n724) );
  XNOR2_X1 U784 ( .A(KEYINPUT111), .B(KEYINPUT29), .ZN(n723) );
  XNOR2_X1 U785 ( .A(n724), .B(n723), .ZN(n725) );
  XOR2_X1 U786 ( .A(G128), .B(n725), .Z(G30) );
  XNOR2_X1 U787 ( .A(n726), .B(G143), .ZN(G45) );
  NOR2_X1 U788 ( .A1(n727), .A2(n480), .ZN(n728) );
  XOR2_X1 U789 ( .A(G146), .B(n728), .Z(G48) );
  NOR2_X1 U790 ( .A1(n731), .A2(n480), .ZN(n729) );
  XOR2_X1 U791 ( .A(G113), .B(n729), .Z(G15) );
  NOR2_X1 U792 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U793 ( .A(KEYINPUT112), .B(n732), .Z(n733) );
  XNOR2_X1 U794 ( .A(G116), .B(n733), .ZN(G18) );
  XOR2_X1 U795 ( .A(KEYINPUT37), .B(KEYINPUT113), .Z(n735) );
  XNOR2_X1 U796 ( .A(G125), .B(n515), .ZN(n734) );
  XNOR2_X1 U797 ( .A(n735), .B(n734), .ZN(G27) );
  XOR2_X1 U798 ( .A(G140), .B(n736), .Z(G42) );
  XOR2_X1 U799 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n740) );
  OR2_X1 U800 ( .A1(n477), .A2(n737), .ZN(n739) );
  XNOR2_X1 U801 ( .A(n740), .B(n739), .ZN(n745) );
  NAND2_X1 U802 ( .A1(n425), .A2(n741), .ZN(n743) );
  XOR2_X1 U803 ( .A(KEYINPUT49), .B(n743), .Z(n744) );
  NAND2_X1 U804 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U805 ( .A1(n452), .A2(n746), .ZN(n748) );
  NOR2_X1 U806 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U807 ( .A(n750), .B(KEYINPUT51), .ZN(n751) );
  XNOR2_X1 U808 ( .A(n751), .B(KEYINPUT116), .ZN(n752) );
  NAND2_X1 U809 ( .A1(n768), .A2(n752), .ZN(n762) );
  INV_X1 U810 ( .A(n393), .ZN(n754) );
  NAND2_X1 U811 ( .A1(n368), .A2(n754), .ZN(n759) );
  NAND2_X1 U812 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U813 ( .A1(n757), .A2(n365), .ZN(n758) );
  NAND2_X1 U814 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U815 ( .A1(n361), .A2(n760), .ZN(n761) );
  NAND2_X1 U816 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U817 ( .A(KEYINPUT52), .B(n763), .ZN(n764) );
  NAND2_X1 U818 ( .A1(n764), .A2(G952), .ZN(n765) );
  NOR2_X1 U819 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U820 ( .A(n767), .B(KEYINPUT117), .ZN(n771) );
  NAND2_X1 U821 ( .A1(n361), .A2(n768), .ZN(n770) );
  NAND2_X1 U822 ( .A1(n771), .A2(n770), .ZN(n775) );
  INV_X1 U823 ( .A(n772), .ZN(n773) );
  NOR2_X1 U824 ( .A1(n773), .A2(n367), .ZN(n774) );
  NAND2_X1 U825 ( .A1(n395), .A2(G469), .ZN(n780) );
  XOR2_X1 U826 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n778) );
  XNOR2_X1 U827 ( .A(n776), .B(KEYINPUT120), .ZN(n777) );
  XNOR2_X1 U828 ( .A(n778), .B(n777), .ZN(n779) );
  XNOR2_X1 U829 ( .A(n780), .B(n779), .ZN(n781) );
  NOR2_X1 U830 ( .A1(n782), .A2(n781), .ZN(G54) );
  NOR2_X1 U831 ( .A1(n784), .A2(n783), .ZN(n786) );
  XNOR2_X1 U832 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n785) );
  XNOR2_X1 U833 ( .A(n786), .B(n785), .ZN(n794) );
  XOR2_X1 U834 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n788) );
  NAND2_X1 U835 ( .A1(G224), .A2(G953), .ZN(n787) );
  XNOR2_X1 U836 ( .A(n788), .B(n787), .ZN(n789) );
  NAND2_X1 U837 ( .A1(n789), .A2(G898), .ZN(n792) );
  OR2_X1 U838 ( .A1(n396), .A2(G953), .ZN(n791) );
  NAND2_X1 U839 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U840 ( .A(n794), .B(n793), .Z(G69) );
  XNOR2_X1 U841 ( .A(n796), .B(n795), .ZN(n800) );
  XNOR2_X1 U842 ( .A(n394), .B(n800), .ZN(n799) );
  NAND2_X1 U843 ( .A1(n799), .A2(n798), .ZN(n806) );
  XNOR2_X1 U844 ( .A(G227), .B(n800), .ZN(n801) );
  XNOR2_X1 U845 ( .A(n801), .B(KEYINPUT126), .ZN(n802) );
  NAND2_X1 U846 ( .A1(n802), .A2(G900), .ZN(n803) );
  NAND2_X1 U847 ( .A1(G953), .A2(n803), .ZN(n804) );
  XOR2_X1 U848 ( .A(KEYINPUT127), .B(n804), .Z(n805) );
  NAND2_X1 U849 ( .A1(n806), .A2(n805), .ZN(G72) );
  XOR2_X1 U850 ( .A(n807), .B(G122), .Z(G24) );
  XOR2_X1 U851 ( .A(n808), .B(G110), .Z(G12) );
  XNOR2_X1 U852 ( .A(n809), .B(G119), .ZN(G21) );
  XNOR2_X1 U853 ( .A(n810), .B(G131), .ZN(G33) );
  XNOR2_X1 U854 ( .A(G137), .B(n811), .ZN(G39) );
endmodule

