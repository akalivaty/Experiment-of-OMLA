

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(n475), .B(KEYINPUT119), .ZN(n567) );
  XOR2_X2 U325 ( .A(n413), .B(n412), .Z(n583) );
  XNOR2_X1 U326 ( .A(n466), .B(KEYINPUT48), .ZN(n544) );
  XOR2_X1 U327 ( .A(n347), .B(n346), .Z(n518) );
  XNOR2_X1 U328 ( .A(KEYINPUT93), .B(n387), .ZN(n546) );
  XOR2_X1 U329 ( .A(n373), .B(n341), .Z(n292) );
  XOR2_X1 U330 ( .A(G211GAT), .B(KEYINPUT85), .Z(n293) );
  XOR2_X1 U331 ( .A(n429), .B(n428), .Z(n294) );
  XNOR2_X1 U332 ( .A(n461), .B(KEYINPUT47), .ZN(n462) );
  XNOR2_X1 U333 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U334 ( .A(n430), .B(n294), .ZN(n431) );
  XNOR2_X1 U335 ( .A(n342), .B(n292), .ZN(n344) );
  XNOR2_X1 U336 ( .A(n432), .B(n431), .ZN(n436) );
  NOR2_X1 U337 ( .A1(n515), .A2(n478), .ZN(n450) );
  INV_X1 U338 ( .A(KEYINPUT100), .ZN(n451) );
  XNOR2_X1 U339 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n476) );
  XNOR2_X1 U340 ( .A(n451), .B(G36GAT), .ZN(n452) );
  XNOR2_X1 U341 ( .A(n477), .B(n476), .ZN(G1350GAT) );
  XNOR2_X1 U342 ( .A(n453), .B(n452), .ZN(G1329GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n296) );
  XNOR2_X1 U344 ( .A(KEYINPUT73), .B(KEYINPUT9), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U346 ( .A(G92GAT), .B(G106GAT), .Z(n298) );
  XNOR2_X1 U347 ( .A(G134GAT), .B(G162GAT), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U349 ( .A(n300), .B(n299), .Z(n302) );
  XOR2_X1 U350 ( .A(G190GAT), .B(G218GAT), .Z(n343) );
  XOR2_X1 U351 ( .A(G99GAT), .B(G85GAT), .Z(n418) );
  XNOR2_X1 U352 ( .A(n343), .B(n418), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U354 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n304) );
  NAND2_X1 U355 ( .A1(G232GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U357 ( .A(n306), .B(n305), .Z(n313) );
  XOR2_X1 U358 ( .A(G29GAT), .B(KEYINPUT7), .Z(n308) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G36GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n310) );
  XOR2_X1 U361 ( .A(G50GAT), .B(KEYINPUT8), .Z(n309) );
  XOR2_X1 U362 ( .A(n310), .B(n309), .Z(n448) );
  INV_X1 U363 ( .A(n448), .ZN(n311) );
  XOR2_X1 U364 ( .A(n311), .B(KEYINPUT72), .Z(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n566) );
  XNOR2_X1 U366 ( .A(KEYINPUT36), .B(KEYINPUT97), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n566), .B(n314), .ZN(n587) );
  XOR2_X1 U368 ( .A(G113GAT), .B(G1GAT), .Z(n441) );
  XOR2_X1 U369 ( .A(KEYINPUT87), .B(KEYINPUT1), .Z(n316) );
  XNOR2_X1 U370 ( .A(G29GAT), .B(G85GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U372 ( .A(n441), .B(n317), .Z(n319) );
  NAND2_X1 U373 ( .A1(G225GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n331) );
  XOR2_X1 U375 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n321) );
  XNOR2_X1 U376 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U378 ( .A(KEYINPUT88), .B(KEYINPUT5), .Z(n323) );
  XNOR2_X1 U379 ( .A(KEYINPUT92), .B(KEYINPUT91), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U381 ( .A(n325), .B(n324), .Z(n329) );
  XNOR2_X1 U382 ( .A(G134GAT), .B(G127GAT), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n326), .B(KEYINPUT0), .ZN(n364) );
  XNOR2_X1 U384 ( .A(G120GAT), .B(G148GAT), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n327), .B(G57GAT), .ZN(n434) );
  XNOR2_X1 U386 ( .A(n364), .B(n434), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U389 ( .A(KEYINPUT2), .B(G162GAT), .Z(n333) );
  XNOR2_X1 U390 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U392 ( .A(G141GAT), .B(n334), .ZN(n378) );
  XNOR2_X1 U393 ( .A(n335), .B(n378), .ZN(n387) );
  XOR2_X1 U394 ( .A(G183GAT), .B(KEYINPUT17), .Z(n337) );
  XNOR2_X1 U395 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n363) );
  XNOR2_X1 U397 ( .A(G36GAT), .B(n363), .ZN(n342) );
  XNOR2_X1 U398 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n293), .B(n338), .ZN(n373) );
  XOR2_X1 U400 ( .A(G204GAT), .B(KEYINPUT74), .Z(n340) );
  NAND2_X1 U401 ( .A1(G226GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U403 ( .A(n344), .B(n343), .Z(n347) );
  XOR2_X1 U404 ( .A(G169GAT), .B(G8GAT), .Z(n440) );
  XNOR2_X1 U405 ( .A(G176GAT), .B(G92GAT), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n345), .B(G64GAT), .ZN(n433) );
  XNOR2_X1 U407 ( .A(n440), .B(n433), .ZN(n346) );
  XOR2_X1 U408 ( .A(n518), .B(KEYINPUT27), .Z(n389) );
  INV_X1 U409 ( .A(n389), .ZN(n382) );
  XOR2_X1 U410 ( .A(G120GAT), .B(G190GAT), .Z(n349) );
  XNOR2_X1 U411 ( .A(G43GAT), .B(G99GAT), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U413 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n351) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G113GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U416 ( .A(n353), .B(n352), .Z(n358) );
  XOR2_X1 U417 ( .A(KEYINPUT81), .B(G176GAT), .Z(n355) );
  NAND2_X1 U418 ( .A1(G227GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U420 ( .A(G15GAT), .B(n356), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U422 ( .A(KEYINPUT80), .B(KEYINPUT82), .Z(n360) );
  XNOR2_X1 U423 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U425 ( .A(n362), .B(n361), .Z(n366) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U427 ( .A(n366), .B(n365), .Z(n529) );
  XOR2_X1 U428 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n372) );
  XOR2_X1 U429 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n368) );
  XNOR2_X1 U430 ( .A(G22GAT), .B(G148GAT), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n370) );
  XNOR2_X1 U432 ( .A(G106GAT), .B(G78GAT), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n369), .B(G204GAT), .ZN(n427) );
  XNOR2_X1 U434 ( .A(n370), .B(n427), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n377) );
  XOR2_X1 U436 ( .A(G218GAT), .B(n373), .Z(n375) );
  NAND2_X1 U437 ( .A1(G228GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U439 ( .A(n377), .B(n376), .Z(n380) );
  XOR2_X1 U440 ( .A(G50GAT), .B(n378), .Z(n379) );
  XOR2_X1 U441 ( .A(n380), .B(n379), .Z(n388) );
  INV_X1 U442 ( .A(n388), .ZN(n471) );
  NAND2_X1 U443 ( .A1(n529), .A2(n471), .ZN(n381) );
  XNOR2_X1 U444 ( .A(n381), .B(KEYINPUT26), .ZN(n574) );
  NOR2_X1 U445 ( .A1(n382), .A2(n574), .ZN(n543) );
  INV_X1 U446 ( .A(n518), .ZN(n467) );
  INV_X1 U447 ( .A(n529), .ZN(n473) );
  NAND2_X1 U448 ( .A1(n467), .A2(n473), .ZN(n383) );
  NAND2_X1 U449 ( .A1(n383), .A2(n388), .ZN(n384) );
  XNOR2_X1 U450 ( .A(KEYINPUT25), .B(n384), .ZN(n385) );
  NOR2_X1 U451 ( .A1(n543), .A2(n385), .ZN(n386) );
  NOR2_X1 U452 ( .A1(n387), .A2(n386), .ZN(n392) );
  XOR2_X1 U453 ( .A(n388), .B(KEYINPUT28), .Z(n492) );
  NOR2_X1 U454 ( .A1(n546), .A2(n492), .ZN(n390) );
  NAND2_X1 U455 ( .A1(n390), .A2(n389), .ZN(n528) );
  NOR2_X1 U456 ( .A1(n473), .A2(n528), .ZN(n391) );
  NOR2_X1 U457 ( .A1(n392), .A2(n391), .ZN(n479) );
  XOR2_X1 U458 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n394) );
  XNOR2_X1 U459 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n393) );
  XNOR2_X1 U460 ( .A(n394), .B(n393), .ZN(n413) );
  XOR2_X1 U461 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n396) );
  XNOR2_X1 U462 ( .A(G8GAT), .B(KEYINPUT74), .ZN(n395) );
  XNOR2_X1 U463 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U464 ( .A(G64GAT), .B(G57GAT), .Z(n398) );
  XNOR2_X1 U465 ( .A(G1GAT), .B(G211GAT), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n400), .B(n399), .ZN(n411) );
  XOR2_X1 U468 ( .A(G15GAT), .B(G22GAT), .Z(n444) );
  XOR2_X1 U469 ( .A(G78GAT), .B(G155GAT), .Z(n402) );
  XNOR2_X1 U470 ( .A(G127GAT), .B(G183GAT), .ZN(n401) );
  XNOR2_X1 U471 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U472 ( .A(n444), .B(n403), .Z(n405) );
  NAND2_X1 U473 ( .A1(G231GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U475 ( .A(n406), .B(KEYINPUT15), .Z(n409) );
  XNOR2_X1 U476 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n407), .B(KEYINPUT66), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n419), .B(KEYINPUT14), .ZN(n408) );
  XNOR2_X1 U479 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n412) );
  NOR2_X1 U481 ( .A1(n479), .A2(n583), .ZN(n414) );
  XOR2_X1 U482 ( .A(KEYINPUT98), .B(n414), .Z(n415) );
  NOR2_X1 U483 ( .A1(n587), .A2(n415), .ZN(n416) );
  XOR2_X1 U484 ( .A(n416), .B(KEYINPUT37), .Z(n417) );
  XNOR2_X1 U485 ( .A(KEYINPUT99), .B(n417), .ZN(n515) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n420) );
  AND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n421) );
  NAND2_X1 U488 ( .A1(n420), .A2(n421), .ZN(n425) );
  INV_X1 U489 ( .A(n420), .ZN(n423) );
  INV_X1 U490 ( .A(n421), .ZN(n422) );
  NAND2_X1 U491 ( .A1(n423), .A2(n422), .ZN(n424) );
  NAND2_X1 U492 ( .A1(n425), .A2(n424), .ZN(n426) );
  XOR2_X1 U493 ( .A(n426), .B(KEYINPUT68), .Z(n432) );
  XNOR2_X1 U494 ( .A(n427), .B(KEYINPUT69), .ZN(n430) );
  XOR2_X1 U495 ( .A(KEYINPUT67), .B(KEYINPUT33), .Z(n429) );
  XNOR2_X1 U496 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n428) );
  XNOR2_X1 U497 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n578) );
  XOR2_X1 U499 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n438) );
  NAND2_X1 U500 ( .A1(G229GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U502 ( .A(n439), .B(KEYINPUT64), .Z(n443) );
  XNOR2_X1 U503 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U505 ( .A(n445), .B(n444), .Z(n447) );
  XNOR2_X1 U506 ( .A(G141GAT), .B(G197GAT), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U508 ( .A(n449), .B(n448), .Z(n502) );
  INV_X1 U509 ( .A(n502), .ZN(n575) );
  XOR2_X1 U510 ( .A(KEYINPUT65), .B(n575), .Z(n558) );
  NAND2_X1 U511 ( .A1(n578), .A2(n558), .ZN(n478) );
  XOR2_X1 U512 ( .A(KEYINPUT38), .B(n450), .Z(n500) );
  NOR2_X1 U513 ( .A1(n500), .A2(n518), .ZN(n453) );
  INV_X1 U514 ( .A(KEYINPUT45), .ZN(n455) );
  INV_X1 U515 ( .A(n583), .ZN(n480) );
  NOR2_X1 U516 ( .A1(n587), .A2(n480), .ZN(n454) );
  XNOR2_X1 U517 ( .A(n455), .B(n454), .ZN(n456) );
  NOR2_X1 U518 ( .A1(n558), .A2(n456), .ZN(n457) );
  NAND2_X1 U519 ( .A1(n578), .A2(n457), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n578), .B(KEYINPUT41), .ZN(n561) );
  NAND2_X1 U521 ( .A1(n575), .A2(n561), .ZN(n458) );
  XNOR2_X1 U522 ( .A(KEYINPUT46), .B(n458), .ZN(n460) );
  NOR2_X1 U523 ( .A1(n566), .A2(n583), .ZN(n459) );
  NAND2_X1 U524 ( .A1(n460), .A2(n459), .ZN(n463) );
  XNOR2_X1 U525 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n461) );
  NAND2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n544), .A2(n467), .ZN(n469) );
  XOR2_X1 U528 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n468) );
  XNOR2_X1 U529 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n546), .A2(n470), .ZN(n573) );
  NOR2_X1 U531 ( .A1(n471), .A2(n573), .ZN(n472) );
  XOR2_X1 U532 ( .A(KEYINPUT55), .B(n472), .Z(n474) );
  NAND2_X1 U533 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n567), .A2(n583), .ZN(n477) );
  INV_X1 U535 ( .A(n478), .ZN(n483) );
  NOR2_X1 U536 ( .A1(n566), .A2(n480), .ZN(n481) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n481), .Z(n482) );
  NOR2_X1 U538 ( .A1(n479), .A2(n482), .ZN(n503) );
  NAND2_X1 U539 ( .A1(n483), .A2(n503), .ZN(n493) );
  NOR2_X1 U540 ( .A1(n546), .A2(n493), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT34), .B(n484), .Z(n485) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U543 ( .A1(n518), .A2(n493), .ZN(n486) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  NOR2_X1 U545 ( .A1(n529), .A2(n493), .ZN(n491) );
  XOR2_X1 U546 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n488) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U549 ( .A(KEYINPUT94), .B(n489), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  INV_X1 U551 ( .A(n492), .ZN(n525) );
  NOR2_X1 U552 ( .A1(n525), .A2(n493), .ZN(n494) );
  XOR2_X1 U553 ( .A(G22GAT), .B(n494), .Z(G1327GAT) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n496) );
  NOR2_X1 U555 ( .A1(n546), .A2(n500), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U557 ( .A1(n500), .A2(n529), .ZN(n498) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n525), .A2(n500), .ZN(n501) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  NAND2_X1 U563 ( .A1(n502), .A2(n561), .ZN(n514) );
  INV_X1 U564 ( .A(n514), .ZN(n504) );
  NAND2_X1 U565 ( .A1(n504), .A2(n503), .ZN(n510) );
  NOR2_X1 U566 ( .A1(n546), .A2(n510), .ZN(n505) );
  XOR2_X1 U567 ( .A(n505), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n518), .A2(n510), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT102), .B(n507), .Z(n508) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U572 ( .A1(n529), .A2(n510), .ZN(n509) );
  XOR2_X1 U573 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U574 ( .A1(n525), .A2(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(KEYINPUT43), .B(KEYINPUT103), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U577 ( .A(G78GAT), .B(n513), .Z(G1335GAT) );
  OR2_X1 U578 ( .A1(n515), .A2(n514), .ZN(n524) );
  NOR2_X1 U579 ( .A1(n546), .A2(n524), .ZN(n516) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n516), .Z(n517) );
  XNOR2_X1 U581 ( .A(KEYINPUT104), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n524), .ZN(n519) );
  XOR2_X1 U583 ( .A(G92GAT), .B(n519), .Z(G1337GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n524), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(KEYINPUT105), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n527) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U591 ( .A(n527), .B(n526), .Z(G1339GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n533) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U594 ( .A1(n530), .A2(n544), .ZN(n531) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(n531), .Z(n539) );
  NAND2_X1 U596 ( .A1(n539), .A2(n558), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U600 ( .A1(n539), .A2(n561), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  NAND2_X1 U602 ( .A1(n539), .A2(n583), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U606 ( .A1(n566), .A2(n539), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U608 ( .A(G134GAT), .B(n542), .Z(G1343GAT) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n575), .A2(n555), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n547), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n549) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(KEYINPUT114), .B(n550), .Z(n552) );
  NAND2_X1 U617 ( .A1(n555), .A2(n561), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n555), .A2(n583), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT116), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  XOR2_X1 U622 ( .A(G162GAT), .B(KEYINPUT117), .Z(n557) );
  NAND2_X1 U623 ( .A1(n555), .A2(n566), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1347GAT) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n567), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n567), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(n570), .ZN(G1351GAT) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT124), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(n572), .Z(n577) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n584) );
  NAND2_X1 U641 ( .A1(n584), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  INV_X1 U643 ( .A(n584), .ZN(n586) );
  NOR2_X1 U644 ( .A1(n586), .A2(n578), .ZN(n582) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

