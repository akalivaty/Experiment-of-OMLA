

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n426) );
  NOR2_X1 U327 ( .A1(n546), .A2(n450), .ZN(n588) );
  AND2_X1 U328 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  AND2_X1 U329 ( .A1(n569), .A2(n582), .ZN(n385) );
  XNOR2_X1 U330 ( .A(n350), .B(n294), .ZN(n352) );
  XNOR2_X1 U331 ( .A(n352), .B(n399), .ZN(n353) );
  NOR2_X1 U332 ( .A1(n414), .A2(n413), .ZN(n415) );
  XNOR2_X1 U333 ( .A(n427), .B(n426), .ZN(n561) );
  XOR2_X1 U334 ( .A(KEYINPUT48), .B(n415), .Z(n547) );
  XNOR2_X1 U335 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U336 ( .A(n364), .B(n363), .ZN(n585) );
  XNOR2_X1 U337 ( .A(n411), .B(KEYINPUT41), .ZN(n569) );
  XOR2_X1 U338 ( .A(n383), .B(n382), .Z(n582) );
  XOR2_X1 U339 ( .A(n422), .B(n348), .Z(n524) );
  XNOR2_X1 U340 ( .A(n452), .B(G218GAT), .ZN(n453) );
  XNOR2_X1 U341 ( .A(n454), .B(n453), .ZN(G1355GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT10), .B(KEYINPUT77), .Z(n296) );
  XNOR2_X1 U343 ( .A(KEYINPUT11), .B(KEYINPUT78), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n313) );
  XOR2_X1 U345 ( .A(KEYINPUT9), .B(G92GAT), .Z(n298) );
  XNOR2_X1 U346 ( .A(G218GAT), .B(KEYINPUT79), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U348 ( .A(KEYINPUT80), .B(KEYINPUT65), .Z(n300) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(KEYINPUT76), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U351 ( .A(n302), .B(n301), .Z(n311) );
  XNOR2_X1 U352 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n303), .B(KEYINPUT7), .ZN(n371) );
  XOR2_X1 U354 ( .A(G106GAT), .B(n371), .Z(n305) );
  NAND2_X1 U355 ( .A1(G232GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U357 ( .A(G36GAT), .B(G190GAT), .Z(n416) );
  XOR2_X1 U358 ( .A(G85GAT), .B(KEYINPUT74), .Z(n350) );
  XOR2_X1 U359 ( .A(n416), .B(n350), .Z(n307) );
  XOR2_X1 U360 ( .A(G43GAT), .B(G134GAT), .Z(n337) );
  XOR2_X1 U361 ( .A(G50GAT), .B(G162GAT), .Z(n323) );
  XNOR2_X1 U362 ( .A(n337), .B(n323), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U366 ( .A(n313), .B(n312), .Z(n575) );
  XOR2_X1 U367 ( .A(KEYINPUT36), .B(n575), .Z(n486) );
  XNOR2_X1 U368 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n314), .B(KEYINPUT90), .ZN(n315) );
  XOR2_X1 U370 ( .A(n315), .B(KEYINPUT91), .Z(n317) );
  XNOR2_X1 U371 ( .A(G197GAT), .B(G218GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n421) );
  XOR2_X1 U373 ( .A(G78GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n354) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n320), .B(KEYINPUT2), .ZN(n436) );
  XNOR2_X1 U378 ( .A(n354), .B(n436), .ZN(n331) );
  XOR2_X1 U379 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n322) );
  XNOR2_X1 U380 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U382 ( .A(KEYINPUT92), .B(KEYINPUT23), .Z(n325) );
  XOR2_X1 U383 ( .A(G22GAT), .B(G155GAT), .Z(n390) );
  XNOR2_X1 U384 ( .A(n323), .B(n390), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U386 ( .A(n327), .B(n326), .Z(n329) );
  NAND2_X1 U387 ( .A1(G228GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n421), .B(n332), .ZN(n559) );
  XNOR2_X1 U391 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n333), .B(KEYINPUT18), .ZN(n334) );
  XOR2_X1 U393 ( .A(n334), .B(KEYINPUT17), .Z(n336) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(G176GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n422) );
  XOR2_X1 U396 ( .A(G113GAT), .B(G15GAT), .Z(n370) );
  XNOR2_X1 U397 ( .A(n370), .B(n337), .ZN(n347) );
  XOR2_X1 U398 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n339) );
  NAND2_X1 U399 ( .A1(G227GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U401 ( .A(n340), .B(G190GAT), .Z(n345) );
  XNOR2_X1 U402 ( .A(G99GAT), .B(G71GAT), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n341), .B(G120GAT), .ZN(n358) );
  XOR2_X1 U404 ( .A(G127GAT), .B(KEYINPUT86), .Z(n343) );
  XNOR2_X1 U405 ( .A(KEYINPUT0), .B(KEYINPUT85), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n437) );
  XNOR2_X1 U407 ( .A(n358), .B(n437), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n348) );
  INV_X1 U410 ( .A(n524), .ZN(n564) );
  NAND2_X1 U411 ( .A1(n559), .A2(n564), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n349), .B(KEYINPUT26), .ZN(n546) );
  XNOR2_X1 U413 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n351), .B(KEYINPUT71), .ZN(n399) );
  XOR2_X1 U415 ( .A(n353), .B(KEYINPUT32), .Z(n356) );
  XNOR2_X1 U416 ( .A(n354), .B(KEYINPUT72), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n364) );
  XNOR2_X1 U418 ( .A(G204GAT), .B(G92GAT), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n357), .B(G64GAT), .ZN(n419) );
  XNOR2_X1 U420 ( .A(n358), .B(n419), .ZN(n362) );
  XOR2_X1 U421 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n360) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  INV_X1 U424 ( .A(n585), .ZN(n411) );
  XOR2_X1 U425 ( .A(G197GAT), .B(G22GAT), .Z(n366) );
  XNOR2_X1 U426 ( .A(G36GAT), .B(G141GAT), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U428 ( .A(n367), .B(G50GAT), .Z(n369) );
  XOR2_X1 U429 ( .A(G1GAT), .B(G8GAT), .Z(n391) );
  XNOR2_X1 U430 ( .A(n391), .B(G43GAT), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n375) );
  XOR2_X1 U432 ( .A(n371), .B(n370), .Z(n373) );
  NAND2_X1 U433 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U435 ( .A(n375), .B(n374), .Z(n383) );
  XOR2_X1 U436 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n377) );
  XNOR2_X1 U437 ( .A(G169GAT), .B(KEYINPUT70), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U439 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n379) );
  XNOR2_X1 U440 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U443 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n404) );
  XOR2_X1 U445 ( .A(G127GAT), .B(G71GAT), .Z(n387) );
  XNOR2_X1 U446 ( .A(G15GAT), .B(G183GAT), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n403) );
  XOR2_X1 U448 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n389) );
  XNOR2_X1 U449 ( .A(G64GAT), .B(KEYINPUT82), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n395) );
  XOR2_X1 U451 ( .A(n390), .B(G78GAT), .Z(n393) );
  XNOR2_X1 U452 ( .A(n391), .B(G211GAT), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U454 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U457 ( .A(n398), .B(KEYINPUT81), .Z(n401) );
  XNOR2_X1 U458 ( .A(n399), .B(KEYINPUT12), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U460 ( .A(n403), .B(n402), .Z(n484) );
  INV_X1 U461 ( .A(n484), .ZN(n589) );
  NOR2_X1 U462 ( .A1(n404), .A2(n589), .ZN(n405) );
  INV_X1 U463 ( .A(n575), .ZN(n456) );
  NAND2_X1 U464 ( .A1(n405), .A2(n456), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n406), .B(KEYINPUT47), .ZN(n414) );
  XNOR2_X1 U466 ( .A(KEYINPUT111), .B(KEYINPUT45), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n407), .B(KEYINPUT64), .ZN(n409) );
  NOR2_X1 U468 ( .A1(n484), .A2(n486), .ZN(n408) );
  XOR2_X1 U469 ( .A(n409), .B(n408), .Z(n410) );
  NAND2_X1 U470 ( .A1(n411), .A2(n410), .ZN(n412) );
  NOR2_X1 U471 ( .A1(n582), .A2(n412), .ZN(n413) );
  XOR2_X1 U472 ( .A(n416), .B(G8GAT), .Z(n418) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n420) );
  XOR2_X1 U475 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U477 ( .A(n424), .B(n423), .Z(n496) );
  XNOR2_X1 U478 ( .A(n496), .B(KEYINPUT119), .ZN(n425) );
  AND2_X1 U479 ( .A1(n547), .A2(n425), .ZN(n427) );
  XOR2_X1 U480 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n429) );
  XNOR2_X1 U481 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n441) );
  XOR2_X1 U483 ( .A(G155GAT), .B(G120GAT), .Z(n431) );
  XNOR2_X1 U484 ( .A(G113GAT), .B(G1GAT), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U486 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n433) );
  XNOR2_X1 U487 ( .A(G57GAT), .B(KEYINPUT6), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U489 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n449) );
  NAND2_X1 U493 ( .A1(G225GAT), .A2(G233GAT), .ZN(n447) );
  XOR2_X1 U494 ( .A(G85GAT), .B(G162GAT), .Z(n443) );
  XNOR2_X1 U495 ( .A(G29GAT), .B(G148GAT), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U497 ( .A(G134GAT), .B(KEYINPUT79), .Z(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U500 ( .A(n449), .B(n448), .Z(n558) );
  INV_X1 U501 ( .A(n558), .ZN(n491) );
  NAND2_X1 U502 ( .A1(n561), .A2(n491), .ZN(n450) );
  INV_X1 U503 ( .A(n588), .ZN(n451) );
  NOR2_X1 U504 ( .A1(n486), .A2(n451), .ZN(n454) );
  XNOR2_X1 U505 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n452) );
  INV_X1 U506 ( .A(n582), .ZN(n455) );
  NOR2_X1 U507 ( .A1(n455), .A2(n585), .ZN(n488) );
  NAND2_X1 U508 ( .A1(n456), .A2(n589), .ZN(n459) );
  XNOR2_X1 U509 ( .A(KEYINPUT16), .B(KEYINPUT84), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n457), .B(KEYINPUT83), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n459), .B(n458), .ZN(n471) );
  XOR2_X1 U512 ( .A(n524), .B(KEYINPUT88), .Z(n460) );
  XOR2_X1 U513 ( .A(KEYINPUT28), .B(n559), .Z(n500) );
  INV_X1 U514 ( .A(n500), .ZN(n526) );
  XNOR2_X1 U515 ( .A(n496), .B(KEYINPUT27), .ZN(n461) );
  OR2_X1 U516 ( .A1(n491), .A2(n461), .ZN(n545) );
  NOR2_X1 U517 ( .A1(n526), .A2(n545), .ZN(n530) );
  NAND2_X1 U518 ( .A1(n460), .A2(n530), .ZN(n470) );
  NOR2_X1 U519 ( .A1(n546), .A2(n461), .ZN(n462) );
  XOR2_X1 U520 ( .A(KEYINPUT96), .B(n462), .Z(n467) );
  INV_X1 U521 ( .A(n496), .ZN(n521) );
  NAND2_X1 U522 ( .A1(n524), .A2(n521), .ZN(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT97), .B(n463), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n559), .A2(n464), .ZN(n465) );
  XNOR2_X1 U525 ( .A(KEYINPUT25), .B(n465), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n491), .A2(n468), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n483) );
  NAND2_X1 U529 ( .A1(n471), .A2(n483), .ZN(n507) );
  INV_X1 U530 ( .A(n507), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n488), .A2(n472), .ZN(n480) );
  NOR2_X1 U532 ( .A1(n491), .A2(n480), .ZN(n474) );
  XNOR2_X1 U533 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U535 ( .A(G1GAT), .B(n475), .Z(G1324GAT) );
  NOR2_X1 U536 ( .A1(n496), .A2(n480), .ZN(n477) );
  XNOR2_X1 U537 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(G1325GAT) );
  NOR2_X1 U539 ( .A1(n564), .A2(n480), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n500), .A2(n480), .ZN(n481) );
  XOR2_X1 U543 ( .A(KEYINPUT100), .B(n481), .Z(n482) );
  XNOR2_X1 U544 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  NAND2_X1 U545 ( .A1(n484), .A2(n483), .ZN(n485) );
  NOR2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(KEYINPUT37), .B(n487), .ZN(n519) );
  INV_X1 U548 ( .A(n519), .ZN(n489) );
  NAND2_X1 U549 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT38), .B(n490), .ZN(n501) );
  NOR2_X1 U551 ( .A1(n491), .A2(n501), .ZN(n495) );
  XOR2_X1 U552 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n493) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n501), .A2(n496), .ZN(n497) );
  XOR2_X1 U557 ( .A(G36GAT), .B(n497), .Z(G1329GAT) );
  NOR2_X1 U558 ( .A1(n501), .A2(n564), .ZN(n498) );
  XOR2_X1 U559 ( .A(KEYINPUT40), .B(n498), .Z(n499) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n501), .A2(n500), .ZN(n503) );
  XNOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT103), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U564 ( .A(G50GAT), .B(n504), .ZN(G1331GAT) );
  INV_X1 U565 ( .A(n569), .ZN(n505) );
  NOR2_X1 U566 ( .A1(n582), .A2(n505), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n506), .B(KEYINPUT105), .ZN(n518) );
  NOR2_X1 U568 ( .A1(n507), .A2(n518), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n508), .B(KEYINPUT106), .ZN(n515) );
  NAND2_X1 U570 ( .A1(n515), .A2(n558), .ZN(n512) );
  XOR2_X1 U571 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n510) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n515), .A2(n521), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n513), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n515), .A2(n524), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U580 ( .A1(n526), .A2(n515), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n558), .A2(n527), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT109), .Z(n523) );
  NAND2_X1 U586 ( .A1(n527), .A2(n521), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n527), .A2(n524), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U593 ( .A1(n547), .A2(n530), .ZN(n531) );
  NOR2_X1 U594 ( .A1(n564), .A2(n531), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n582), .A2(n541), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n532), .B(KEYINPUT112), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n535) );
  NAND2_X1 U599 ( .A1(n541), .A2(n569), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT113), .Z(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n539) );
  NAND2_X1 U604 ( .A1(n541), .A2(n589), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n575), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(KEYINPUT117), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n582), .A2(n556), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U617 ( .A1(n556), .A2(n569), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n589), .A2(n556), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n575), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  AND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT55), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n576) );
  NAND2_X1 U629 ( .A1(n576), .A2(n582), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n567) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT121), .B(n568), .Z(n571) );
  NAND2_X1 U635 ( .A1(n576), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n576), .A2(n589), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(n574), .ZN(G1350GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G190GAT), .B(n579), .ZN(G1351GAT) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n580), .B(KEYINPUT126), .ZN(n581) );
  XOR2_X1 U647 ( .A(KEYINPUT60), .B(n581), .Z(n584) );
  NAND2_X1 U648 ( .A1(n588), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  NAND2_X1 U651 ( .A1(n585), .A2(n588), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
endmodule

