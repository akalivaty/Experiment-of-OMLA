

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806;

  AND2_X1 U373 ( .A1(n387), .A2(n775), .ZN(n360) );
  AND2_X2 U374 ( .A1(n449), .A2(n448), .ZN(n625) );
  XNOR2_X2 U375 ( .A(n506), .B(G143), .ZN(n554) );
  XNOR2_X2 U376 ( .A(G128), .B(KEYINPUT64), .ZN(n506) );
  XNOR2_X2 U377 ( .A(n603), .B(n593), .ZN(n768) );
  NOR2_X1 U378 ( .A1(n607), .A2(n667), .ZN(n459) );
  NAND2_X1 U379 ( .A1(n355), .A2(n354), .ZN(n362) );
  AND2_X1 U380 ( .A1(n359), .A2(n356), .ZN(n355) );
  AND2_X1 U381 ( .A1(n357), .A2(n353), .ZN(n356) );
  AND2_X2 U382 ( .A1(n387), .A2(n371), .ZN(n774) );
  AND2_X1 U383 ( .A1(n371), .A2(G478), .ZN(n390) );
  NOR2_X1 U384 ( .A1(n626), .A2(n496), .ZN(n702) );
  NOR2_X1 U385 ( .A1(n757), .A2(n659), .ZN(n511) );
  NOR2_X1 U386 ( .A1(n680), .A2(n656), .ZN(n645) );
  NOR2_X1 U387 ( .A1(n619), .A2(n631), .ZN(n620) );
  INV_X1 U388 ( .A(n653), .ZN(n352) );
  XNOR2_X1 U389 ( .A(n499), .B(KEYINPUT67), .ZN(n727) );
  BUF_X1 U390 ( .A(G104), .Z(n587) );
  INV_X1 U391 ( .A(KEYINPUT120), .ZN(n361) );
  XNOR2_X1 U392 ( .A(n362), .B(n361), .ZN(G63) );
  NAND2_X1 U393 ( .A1(n390), .A2(n360), .ZN(n359) );
  AND2_X1 U394 ( .A1(n765), .A2(n371), .ZN(n363) );
  NAND2_X1 U395 ( .A1(n365), .A2(n364), .ZN(n370) );
  OR2_X1 U396 ( .A1(n764), .A2(KEYINPUT2), .ZN(n765) );
  NOR2_X1 U397 ( .A1(n684), .A2(n367), .ZN(n366) );
  INV_X1 U398 ( .A(n684), .ZN(n762) );
  AND2_X1 U399 ( .A1(n477), .A2(n393), .ZN(n473) );
  XNOR2_X1 U400 ( .A(n511), .B(n402), .ZN(n652) );
  XNOR2_X1 U401 ( .A(n624), .B(n623), .ZN(n721) );
  OR2_X1 U402 ( .A1(n406), .A2(n404), .ZN(n744) );
  OR2_X1 U403 ( .A1(n656), .A2(n655), .ZN(n673) );
  XNOR2_X1 U404 ( .A(n641), .B(n642), .ZN(n740) );
  XNOR2_X1 U405 ( .A(n430), .B(KEYINPUT6), .ZN(n653) );
  XNOR2_X1 U406 ( .A(n579), .B(n578), .ZN(n646) );
  AND2_X1 U407 ( .A1(n401), .A2(n427), .ZN(n426) );
  NAND2_X1 U408 ( .A1(n373), .A2(n372), .ZN(n364) );
  OR2_X1 U409 ( .A1(n682), .A2(KEYINPUT65), .ZN(n372) );
  NAND2_X1 U410 ( .A1(n682), .A2(KEYINPUT65), .ZN(n373) );
  XNOR2_X1 U411 ( .A(n486), .B(n550), .ZN(n485) );
  XNOR2_X1 U412 ( .A(n785), .B(n488), .ZN(n592) );
  XNOR2_X1 U413 ( .A(n544), .B(KEYINPUT16), .ZN(n489) );
  XNOR2_X1 U414 ( .A(n553), .B(n552), .ZN(n785) );
  XNOR2_X1 U415 ( .A(n555), .B(G902), .ZN(n628) );
  XNOR2_X1 U416 ( .A(n546), .B(n545), .ZN(n600) );
  INV_X1 U417 ( .A(n777), .ZN(n353) );
  XNOR2_X1 U418 ( .A(KEYINPUT90), .B(KEYINPUT15), .ZN(n555) );
  INV_X2 U419 ( .A(G953), .ZN(n795) );
  OR2_X1 U420 ( .A1(n390), .A2(n775), .ZN(n354) );
  NAND2_X1 U421 ( .A1(n358), .A2(n776), .ZN(n357) );
  INV_X1 U422 ( .A(n387), .ZN(n358) );
  XNOR2_X2 U423 ( .A(n685), .B(KEYINPUT75), .ZN(n371) );
  NAND2_X1 U424 ( .A1(n374), .A2(n366), .ZN(n365) );
  INV_X1 U425 ( .A(n372), .ZN(n367) );
  NAND2_X2 U426 ( .A1(n370), .A2(n368), .ZN(n387) );
  NAND2_X1 U427 ( .A1(n374), .A2(n369), .ZN(n368) );
  NOR2_X1 U428 ( .A1(n684), .A2(KEYINPUT65), .ZN(n369) );
  XNOR2_X2 U429 ( .A(n630), .B(n629), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n650), .B(KEYINPUT1), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n650), .B(KEYINPUT1), .ZN(n613) );
  NAND2_X2 U432 ( .A1(n426), .A2(n423), .ZN(n376) );
  NAND2_X1 U433 ( .A1(n426), .A2(n423), .ZN(n430) );
  BUF_X1 U434 ( .A(n657), .Z(n377) );
  XNOR2_X1 U435 ( .A(n557), .B(n431), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n557), .B(n431), .ZN(n380) );
  NOR2_X1 U437 ( .A1(n622), .A2(n432), .ZN(n604) );
  INV_X1 U438 ( .A(n352), .ZN(n432) );
  XNOR2_X1 U439 ( .A(n459), .B(n609), .ZN(n803) );
  BUF_X1 U440 ( .A(n586), .Z(n379) );
  NAND2_X1 U441 ( .A1(n489), .A2(n600), .ZN(n383) );
  NAND2_X1 U442 ( .A1(n381), .A2(n382), .ZN(n384) );
  NAND2_X1 U443 ( .A1(n384), .A2(n383), .ZN(n784) );
  INV_X1 U444 ( .A(n489), .ZN(n381) );
  INV_X1 U445 ( .A(n600), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n376), .B(KEYINPUT102), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n376), .B(KEYINPUT102), .ZN(n632) );
  XNOR2_X1 U448 ( .A(n412), .B(KEYINPUT101), .ZN(n411) );
  NAND2_X1 U449 ( .A1(n461), .A2(n460), .ZN(n412) );
  XNOR2_X1 U450 ( .A(n490), .B(KEYINPUT100), .ZN(n461) );
  XNOR2_X2 U451 ( .A(n603), .B(n602), .ZN(n701) );
  XNOR2_X1 U452 ( .A(n410), .B(n627), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n410), .B(n627), .ZN(n781) );
  XNOR2_X1 U454 ( .A(n784), .B(n592), .ZN(n487) );
  AND2_X1 U455 ( .A1(n638), .A2(n637), .ZN(n639) );
  OR2_X1 U456 ( .A1(n478), .A2(KEYINPUT85), .ZN(n472) );
  BUF_X1 U457 ( .A(n699), .Z(n388) );
  XNOR2_X1 U458 ( .A(n487), .B(n484), .ZN(n699) );
  XNOR2_X2 U459 ( .A(n565), .B(n394), .ZN(n437) );
  NOR2_X1 U460 ( .A1(G953), .A2(G237), .ZN(n595) );
  OR2_X1 U461 ( .A1(n646), .A2(n729), .ZN(n648) );
  NAND2_X1 U462 ( .A1(n425), .A2(n417), .ZN(n424) );
  NAND2_X1 U463 ( .A1(n422), .A2(n666), .ZN(n421) );
  NAND2_X1 U464 ( .A1(n672), .A2(n471), .ZN(n441) );
  XNOR2_X1 U465 ( .A(n663), .B(n662), .ZN(n471) );
  INV_X1 U466 ( .A(n729), .ZN(n500) );
  XNOR2_X1 U467 ( .A(G113), .B(G101), .ZN(n596) );
  INV_X1 U468 ( .A(G134), .ZN(n584) );
  INV_X1 U469 ( .A(G116), .ZN(n545) );
  OR2_X2 U470 ( .A1(n418), .A2(n415), .ZN(n650) );
  NAND2_X1 U471 ( .A1(n420), .A2(n419), .ZN(n418) );
  NAND2_X1 U472 ( .A1(n494), .A2(G902), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n399), .B(n398), .ZN(n612) );
  INV_X1 U474 ( .A(KEYINPUT77), .ZN(n398) );
  NAND2_X1 U475 ( .A1(n495), .A2(n400), .ZN(n399) );
  AND2_X1 U476 ( .A1(n375), .A2(n496), .ZN(n495) );
  INV_X1 U477 ( .A(KEYINPUT22), .ZN(n450) );
  NAND2_X1 U478 ( .A1(G237), .A2(G234), .ZN(n561) );
  XNOR2_X1 U479 ( .A(n649), .B(n483), .ZN(n482) );
  INV_X1 U480 ( .A(KEYINPUT28), .ZN(n483) );
  XNOR2_X1 U481 ( .A(n409), .B(n408), .ZN(n757) );
  INV_X1 U482 ( .A(KEYINPUT41), .ZN(n408) );
  XNOR2_X1 U483 ( .A(n498), .B(n497), .ZN(n680) );
  INV_X1 U484 ( .A(KEYINPUT39), .ZN(n497) );
  INV_X1 U485 ( .A(KEYINPUT36), .ZN(n513) );
  INV_X1 U486 ( .A(KEYINPUT34), .ZN(n605) );
  INV_X1 U487 ( .A(n702), .ZN(n460) );
  INV_X1 U488 ( .A(KEYINPUT44), .ZN(n462) );
  NAND2_X1 U489 ( .A1(n594), .A2(n417), .ZN(n416) );
  NAND2_X1 U490 ( .A1(n741), .A2(KEYINPUT105), .ZN(n407) );
  XNOR2_X1 U491 ( .A(n653), .B(KEYINPUT78), .ZN(n400) );
  INV_X1 U492 ( .A(G472), .ZN(n425) );
  NAND2_X1 U493 ( .A1(G902), .A2(G472), .ZN(n427) );
  XNOR2_X1 U494 ( .A(G143), .B(KEYINPUT95), .ZN(n519) );
  XNOR2_X1 U495 ( .A(G131), .B(G140), .ZN(n523) );
  XOR2_X1 U496 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n524) );
  XNOR2_X1 U497 ( .A(n501), .B(G146), .ZN(n574) );
  XNOR2_X1 U498 ( .A(KEYINPUT10), .B(G125), .ZN(n501) );
  XNOR2_X1 U499 ( .A(n549), .B(n551), .ZN(n486) );
  XOR2_X1 U500 ( .A(KEYINPUT17), .B(KEYINPUT76), .Z(n549) );
  XNOR2_X1 U501 ( .A(n548), .B(n547), .ZN(n550) );
  XNOR2_X1 U502 ( .A(G125), .B(G146), .ZN(n548) );
  INV_X1 U503 ( .A(KEYINPUT72), .ZN(n488) );
  XNOR2_X1 U504 ( .A(n439), .B(n438), .ZN(n478) );
  INV_X1 U505 ( .A(KEYINPUT48), .ZN(n438) );
  NOR2_X1 U506 ( .A1(n421), .A2(n441), .ZN(n440) );
  NAND2_X1 U507 ( .A1(n476), .A2(n475), .ZN(n474) );
  INV_X1 U508 ( .A(KEYINPUT85), .ZN(n475) );
  INV_X1 U509 ( .A(n726), .ZN(n476) );
  NOR2_X1 U510 ( .A1(G237), .A2(G902), .ZN(n556) );
  XNOR2_X1 U511 ( .A(KEYINPUT5), .B(G137), .ZN(n598) );
  XOR2_X1 U512 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n569) );
  INV_X1 U513 ( .A(KEYINPUT32), .ZN(n435) );
  INV_X1 U514 ( .A(KEYINPUT30), .ZN(n445) );
  NAND2_X1 U515 ( .A1(n482), .A2(n389), .ZN(n661) );
  XNOR2_X1 U516 ( .A(n577), .B(KEYINPUT25), .ZN(n578) );
  NOR2_X1 U517 ( .A1(n686), .A2(G902), .ZN(n579) );
  INV_X1 U518 ( .A(KEYINPUT42), .ZN(n402) );
  XNOR2_X1 U519 ( .A(n514), .B(n512), .ZN(n658) );
  XNOR2_X1 U520 ( .A(n513), .B(KEYINPUT87), .ZN(n512) );
  INV_X1 U521 ( .A(n686), .ZN(n509) );
  INV_X1 U522 ( .A(KEYINPUT60), .ZN(n464) );
  INV_X1 U523 ( .A(KEYINPUT56), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n652), .B(G137), .ZN(G39) );
  AND2_X1 U525 ( .A1(n481), .A2(n651), .ZN(n389) );
  NOR2_X1 U526 ( .A1(n729), .A2(n610), .ZN(n391) );
  AND2_X1 U527 ( .A1(n726), .A2(KEYINPUT85), .ZN(n392) );
  INV_X1 U528 ( .A(G902), .ZN(n417) );
  AND2_X1 U529 ( .A1(n692), .A2(n474), .ZN(n393) );
  INV_X1 U530 ( .A(n375), .ZN(n448) );
  XNOR2_X1 U531 ( .A(n564), .B(KEYINPUT0), .ZN(n394) );
  XOR2_X1 U532 ( .A(n694), .B(n693), .Z(n395) );
  XOR2_X1 U533 ( .A(n388), .B(n698), .Z(n396) );
  XOR2_X1 U534 ( .A(n701), .B(KEYINPUT62), .Z(n397) );
  NAND2_X1 U535 ( .A1(n701), .A2(G472), .ZN(n401) );
  XNOR2_X2 U536 ( .A(n793), .B(G146), .ZN(n603) );
  NAND2_X1 U537 ( .A1(n403), .A2(n407), .ZN(n406) );
  NAND2_X1 U538 ( .A1(n740), .A2(KEYINPUT105), .ZN(n403) );
  NOR2_X1 U539 ( .A1(n740), .A2(n405), .ZN(n404) );
  OR2_X1 U540 ( .A1(n741), .A2(KEYINPUT105), .ZN(n405) );
  NAND2_X1 U541 ( .A1(n744), .A2(n742), .ZN(n409) );
  NAND2_X1 U542 ( .A1(n413), .A2(n411), .ZN(n410) );
  XNOR2_X1 U543 ( .A(n414), .B(n462), .ZN(n413) );
  NAND2_X1 U544 ( .A1(n457), .A2(n458), .ZN(n414) );
  NOR2_X1 U545 ( .A1(n768), .A2(n416), .ZN(n415) );
  NAND2_X1 U546 ( .A1(n768), .A2(n494), .ZN(n420) );
  INV_X1 U547 ( .A(n723), .ZN(n422) );
  OR2_X1 U548 ( .A1(n701), .A2(n424), .ZN(n423) );
  NAND2_X1 U549 ( .A1(n482), .A2(n651), .ZN(n659) );
  INV_X1 U550 ( .A(n661), .ZN(n716) );
  INV_X1 U551 ( .A(n378), .ZN(n641) );
  BUF_X1 U552 ( .A(n793), .Z(n428) );
  INV_X1 U553 ( .A(n452), .ZN(n429) );
  XNOR2_X1 U554 ( .A(n436), .B(n435), .ZN(n806) );
  AND2_X1 U555 ( .A1(n558), .A2(G210), .ZN(n431) );
  INV_X1 U556 ( .A(n660), .ZN(n481) );
  XNOR2_X1 U557 ( .A(n657), .B(n559), .ZN(n660) );
  NAND2_X1 U558 ( .A1(n646), .A2(n500), .ZN(n499) );
  INV_X1 U559 ( .A(n646), .ZN(n496) );
  BUF_X1 U560 ( .A(n784), .Z(n433) );
  BUF_X1 U561 ( .A(n386), .Z(n434) );
  AND2_X1 U562 ( .A1(n456), .A2(n455), .ZN(n454) );
  NAND2_X1 U563 ( .A1(n449), .A2(n447), .ZN(n436) );
  NAND2_X1 U564 ( .A1(n454), .A2(n451), .ZN(n457) );
  NAND2_X1 U565 ( .A1(n437), .A2(n391), .ZN(n611) );
  NAND2_X2 U566 ( .A1(n473), .A2(n472), .ZN(n684) );
  INV_X1 U567 ( .A(n437), .ZN(n619) );
  NAND2_X1 U568 ( .A1(n437), .A2(n736), .ZN(n624) );
  NAND2_X1 U569 ( .A1(n442), .A2(n440), .ZN(n439) );
  XNOR2_X1 U570 ( .A(n444), .B(n443), .ZN(n442) );
  INV_X1 U571 ( .A(KEYINPUT46), .ZN(n443) );
  NAND2_X1 U572 ( .A1(n652), .A2(n690), .ZN(n444) );
  XNOR2_X1 U573 ( .A(n446), .B(n445), .ZN(n638) );
  NAND2_X1 U574 ( .A1(n632), .A2(n674), .ZN(n446) );
  INV_X1 U575 ( .A(n612), .ZN(n447) );
  XNOR2_X2 U576 ( .A(n611), .B(n450), .ZN(n449) );
  INV_X1 U577 ( .A(n803), .ZN(n458) );
  NAND2_X1 U578 ( .A1(n453), .A2(n452), .ZN(n451) );
  INV_X1 U579 ( .A(n806), .ZN(n452) );
  NOR2_X1 U580 ( .A1(n711), .A2(n463), .ZN(n453) );
  NAND2_X1 U581 ( .A1(n711), .A2(n463), .ZN(n455) );
  NAND2_X1 U582 ( .A1(n806), .A2(n463), .ZN(n456) );
  INV_X1 U583 ( .A(KEYINPUT86), .ZN(n463) );
  XNOR2_X1 U584 ( .A(n510), .B(n509), .ZN(n508) );
  XNOR2_X1 U585 ( .A(n505), .B(n397), .ZN(n504) );
  NAND2_X1 U586 ( .A1(n504), .A2(n353), .ZN(n503) );
  NAND2_X1 U587 ( .A1(n508), .A2(n353), .ZN(n507) );
  XNOR2_X1 U588 ( .A(n507), .B(KEYINPUT121), .ZN(G66) );
  XNOR2_X1 U589 ( .A(n503), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U590 ( .A(n465), .B(n464), .ZN(G60) );
  NAND2_X1 U591 ( .A1(n468), .A2(n353), .ZN(n465) );
  XNOR2_X1 U592 ( .A(n467), .B(n466), .ZN(G51) );
  NAND2_X1 U593 ( .A1(n469), .A2(n353), .ZN(n467) );
  XNOR2_X1 U594 ( .A(n695), .B(n395), .ZN(n468) );
  XNOR2_X1 U595 ( .A(n700), .B(n396), .ZN(n469) );
  NAND2_X1 U596 ( .A1(n470), .A2(n621), .ZN(n493) );
  XNOR2_X1 U597 ( .A(n620), .B(KEYINPUT92), .ZN(n470) );
  XNOR2_X2 U598 ( .A(n518), .B(G113), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n478), .A2(n392), .ZN(n477) );
  NAND2_X1 U600 ( .A1(n639), .A2(n479), .ZN(n498) );
  AND2_X1 U601 ( .A1(n640), .A2(n643), .ZN(n479) );
  AND2_X1 U602 ( .A1(n639), .A2(n640), .ZN(n480) );
  NAND2_X1 U603 ( .A1(n480), .A2(n668), .ZN(n689) );
  XNOR2_X1 U604 ( .A(n379), .B(n485), .ZN(n484) );
  INV_X1 U605 ( .A(n493), .ZN(n703) );
  NAND2_X1 U606 ( .A1(n491), .A2(n745), .ZN(n490) );
  NAND2_X1 U607 ( .A1(n493), .A2(n492), .ZN(n491) );
  INV_X1 U608 ( .A(n721), .ZN(n492) );
  INV_X1 U609 ( .A(n594), .ZN(n494) );
  NAND2_X1 U610 ( .A1(n650), .A2(n727), .ZN(n631) );
  AND2_X2 U611 ( .A1(n625), .A2(n502), .ZN(n711) );
  NOR2_X1 U612 ( .A1(n385), .A2(n646), .ZN(n502) );
  NAND2_X1 U613 ( .A1(n774), .A2(G472), .ZN(n505) );
  NAND2_X1 U614 ( .A1(n774), .A2(G217), .ZN(n510) );
  NAND2_X1 U615 ( .A1(n516), .A2(n515), .ZN(n514) );
  INV_X1 U616 ( .A(n377), .ZN(n515) );
  XNOR2_X1 U617 ( .A(n673), .B(n517), .ZN(n516) );
  INV_X1 U618 ( .A(KEYINPUT106), .ZN(n517) );
  NOR2_X2 U619 ( .A1(n684), .A2(n683), .ZN(n685) );
  INV_X1 U620 ( .A(KEYINPUT18), .ZN(n547) );
  XNOR2_X1 U621 ( .A(KEYINPUT23), .B(G119), .ZN(n566) );
  INV_X1 U622 ( .A(KEYINPUT82), .ZN(n629) );
  XNOR2_X1 U623 ( .A(n570), .B(n569), .ZN(n573) );
  XNOR2_X1 U624 ( .A(n573), .B(n572), .ZN(n575) );
  XNOR2_X1 U625 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U626 ( .A(n608), .B(KEYINPUT35), .ZN(n609) );
  INV_X1 U627 ( .A(KEYINPUT40), .ZN(n644) );
  XNOR2_X1 U628 ( .A(n645), .B(n644), .ZN(n690) );
  XNOR2_X2 U629 ( .A(G122), .B(G104), .ZN(n518) );
  XOR2_X1 U630 ( .A(n544), .B(n574), .Z(n528) );
  XOR2_X1 U631 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n520) );
  XNOR2_X1 U632 ( .A(n520), .B(n519), .ZN(n522) );
  NAND2_X1 U633 ( .A1(n595), .A2(G214), .ZN(n521) );
  XNOR2_X1 U634 ( .A(n522), .B(n521), .ZN(n526) );
  XNOR2_X1 U635 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U636 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U637 ( .A(n528), .B(n527), .ZN(n694) );
  NAND2_X1 U638 ( .A1(n694), .A2(n417), .ZN(n530) );
  XOR2_X1 U639 ( .A(KEYINPUT13), .B(G475), .Z(n529) );
  XNOR2_X1 U640 ( .A(n530), .B(n529), .ZN(n617) );
  XOR2_X1 U641 ( .A(KEYINPUT7), .B(G116), .Z(n532) );
  XNOR2_X1 U642 ( .A(G107), .B(G122), .ZN(n531) );
  XNOR2_X1 U643 ( .A(n532), .B(n531), .ZN(n536) );
  XOR2_X1 U644 ( .A(G134), .B(KEYINPUT98), .Z(n534) );
  XNOR2_X1 U645 ( .A(KEYINPUT97), .B(KEYINPUT9), .ZN(n533) );
  XNOR2_X1 U646 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U647 ( .A(n536), .B(n535), .Z(n540) );
  XOR2_X1 U648 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n538) );
  NAND2_X1 U649 ( .A1(G234), .A2(n795), .ZN(n537) );
  XNOR2_X1 U650 ( .A(n538), .B(n537), .ZN(n571) );
  NAND2_X1 U651 ( .A1(G217), .A2(n571), .ZN(n539) );
  XNOR2_X1 U652 ( .A(n540), .B(n539), .ZN(n542) );
  INV_X1 U653 ( .A(n554), .ZN(n541) );
  XNOR2_X1 U654 ( .A(n542), .B(n541), .ZN(n775) );
  NAND2_X1 U655 ( .A1(n775), .A2(n417), .ZN(n543) );
  XNOR2_X1 U656 ( .A(n543), .B(G478), .ZN(n616) );
  NAND2_X1 U657 ( .A1(n617), .A2(n616), .ZN(n667) );
  XNOR2_X1 U658 ( .A(KEYINPUT3), .B(G119), .ZN(n546) );
  NAND2_X1 U659 ( .A1(G224), .A2(n795), .ZN(n551) );
  XOR2_X1 U660 ( .A(G101), .B(G110), .Z(n553) );
  XNOR2_X1 U661 ( .A(G107), .B(KEYINPUT74), .ZN(n552) );
  XNOR2_X2 U662 ( .A(n554), .B(KEYINPUT4), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n699), .A2(n628), .ZN(n557) );
  XNOR2_X1 U664 ( .A(KEYINPUT73), .B(n556), .ZN(n558) );
  NAND2_X1 U665 ( .A1(n558), .A2(G214), .ZN(n674) );
  INV_X1 U666 ( .A(n674), .ZN(n741) );
  NAND2_X1 U667 ( .A1(n380), .A2(n674), .ZN(n657) );
  XOR2_X1 U668 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n559) );
  NOR2_X1 U669 ( .A1(G898), .A2(n795), .ZN(n787) );
  NAND2_X1 U670 ( .A1(n787), .A2(G902), .ZN(n560) );
  NAND2_X1 U671 ( .A1(G952), .A2(n795), .ZN(n634) );
  NAND2_X1 U672 ( .A1(n560), .A2(n634), .ZN(n562) );
  XNOR2_X1 U673 ( .A(n561), .B(KEYINPUT14), .ZN(n753) );
  NAND2_X1 U674 ( .A1(n562), .A2(n753), .ZN(n563) );
  NOR2_X2 U675 ( .A1(n660), .A2(n563), .ZN(n565) );
  INV_X1 U676 ( .A(KEYINPUT89), .ZN(n564) );
  INV_X1 U677 ( .A(n566), .ZN(n568) );
  XNOR2_X1 U678 ( .A(G128), .B(G110), .ZN(n567) );
  XNOR2_X1 U679 ( .A(n568), .B(n567), .ZN(n570) );
  NAND2_X1 U680 ( .A1(G221), .A2(n571), .ZN(n572) );
  XOR2_X1 U681 ( .A(G137), .B(G140), .Z(n588) );
  XNOR2_X1 U682 ( .A(n588), .B(n574), .ZN(n791) );
  XNOR2_X1 U683 ( .A(n575), .B(n791), .ZN(n686) );
  NAND2_X1 U684 ( .A1(n628), .A2(G234), .ZN(n576) );
  XNOR2_X1 U685 ( .A(n576), .B(KEYINPUT20), .ZN(n580) );
  NAND2_X1 U686 ( .A1(G217), .A2(n580), .ZN(n577) );
  NAND2_X1 U687 ( .A1(n580), .A2(G221), .ZN(n581) );
  XNOR2_X1 U688 ( .A(KEYINPUT21), .B(n581), .ZN(n729) );
  XOR2_X1 U689 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n583) );
  XNOR2_X1 U690 ( .A(KEYINPUT71), .B(G469), .ZN(n582) );
  XNOR2_X1 U691 ( .A(n583), .B(n582), .ZN(n594) );
  XNOR2_X1 U692 ( .A(n584), .B(G131), .ZN(n585) );
  XNOR2_X2 U693 ( .A(n586), .B(n585), .ZN(n793) );
  XOR2_X1 U694 ( .A(n587), .B(n588), .Z(n590) );
  NAND2_X1 U695 ( .A1(G227), .A2(n795), .ZN(n589) );
  XNOR2_X1 U696 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U697 ( .A(n592), .B(n591), .ZN(n593) );
  NAND2_X1 U698 ( .A1(n727), .A2(n613), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n595), .A2(G210), .ZN(n597) );
  XNOR2_X1 U700 ( .A(n597), .B(n596), .ZN(n599) );
  XNOR2_X1 U701 ( .A(n599), .B(n598), .ZN(n601) );
  XNOR2_X1 U702 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U703 ( .A(n604), .B(KEYINPUT33), .ZN(n748) );
  NOR2_X1 U704 ( .A1(n748), .A2(n619), .ZN(n606) );
  INV_X1 U705 ( .A(KEYINPUT84), .ZN(n608) );
  NOR2_X1 U706 ( .A1(n617), .A2(n616), .ZN(n742) );
  INV_X1 U707 ( .A(n742), .ZN(n610) );
  INV_X1 U708 ( .A(n617), .ZN(n614) );
  NAND2_X1 U709 ( .A1(n614), .A2(n616), .ZN(n615) );
  XNOR2_X1 U710 ( .A(n615), .B(KEYINPUT99), .ZN(n720) );
  INV_X1 U711 ( .A(n616), .ZN(n618) );
  AND2_X1 U712 ( .A1(n618), .A2(n617), .ZN(n718) );
  NOR2_X1 U713 ( .A1(n720), .A2(n718), .ZN(n669) );
  INV_X1 U714 ( .A(n376), .ZN(n621) );
  NOR2_X1 U715 ( .A1(n622), .A2(n621), .ZN(n736) );
  XOR2_X1 U716 ( .A(KEYINPUT31), .B(KEYINPUT93), .Z(n623) );
  NAND2_X1 U717 ( .A1(n625), .A2(n432), .ZN(n626) );
  XOR2_X1 U718 ( .A(KEYINPUT83), .B(KEYINPUT45), .Z(n627) );
  INV_X1 U719 ( .A(n628), .ZN(n681) );
  NAND2_X1 U720 ( .A1(n781), .A2(n681), .ZN(n630) );
  XNOR2_X1 U721 ( .A(n631), .B(KEYINPUT103), .ZN(n640) );
  NOR2_X1 U722 ( .A1(G900), .A2(n795), .ZN(n633) );
  NAND2_X1 U723 ( .A1(n633), .A2(G902), .ZN(n635) );
  NAND2_X1 U724 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U725 ( .A1(n753), .A2(n636), .ZN(n647) );
  INV_X1 U726 ( .A(n647), .ZN(n637) );
  INV_X1 U727 ( .A(KEYINPUT38), .ZN(n642) );
  INV_X1 U728 ( .A(n740), .ZN(n643) );
  INV_X1 U729 ( .A(n718), .ZN(n656) );
  NOR2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n385), .A2(n654), .ZN(n649) );
  XNOR2_X1 U732 ( .A(n650), .B(KEYINPUT104), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n352), .A2(n654), .ZN(n655) );
  NOR2_X1 U734 ( .A1(n658), .A2(n448), .ZN(n723) );
  NAND2_X1 U735 ( .A1(n661), .A2(KEYINPUT47), .ZN(n663) );
  INV_X1 U736 ( .A(KEYINPUT81), .ZN(n662) );
  INV_X1 U737 ( .A(n669), .ZN(n745) );
  AND2_X1 U738 ( .A1(n716), .A2(n745), .ZN(n665) );
  INV_X1 U739 ( .A(KEYINPUT47), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U741 ( .A1(n641), .A2(n667), .ZN(n668) );
  NAND2_X1 U742 ( .A1(n669), .A2(KEYINPUT47), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n689), .A2(n670), .ZN(n671) );
  XNOR2_X1 U744 ( .A(n671), .B(KEYINPUT79), .ZN(n672) );
  NOR2_X1 U745 ( .A1(n375), .A2(n673), .ZN(n675) );
  AND2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n677) );
  INV_X1 U747 ( .A(KEYINPUT43), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n678), .A2(n641), .ZN(n726) );
  INV_X1 U750 ( .A(n720), .ZN(n679) );
  OR2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n692) );
  NAND2_X1 U752 ( .A1(n681), .A2(KEYINPUT2), .ZN(n682) );
  NAND2_X1 U753 ( .A1(n386), .A2(KEYINPUT2), .ZN(n683) );
  INV_X1 U754 ( .A(G952), .ZN(n687) );
  AND2_X1 U755 ( .A1(n687), .A2(G953), .ZN(n777) );
  XNOR2_X1 U756 ( .A(G143), .B(KEYINPUT112), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n689), .B(n688), .ZN(G45) );
  XNOR2_X1 U758 ( .A(n690), .B(G131), .ZN(G33) );
  XNOR2_X1 U759 ( .A(G134), .B(KEYINPUT114), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n692), .B(n691), .ZN(G36) );
  NAND2_X1 U761 ( .A1(n774), .A2(G475), .ZN(n695) );
  XOR2_X1 U762 ( .A(KEYINPUT119), .B(KEYINPUT59), .Z(n693) );
  NAND2_X1 U763 ( .A1(n774), .A2(G210), .ZN(n700) );
  XNOR2_X1 U764 ( .A(KEYINPUT88), .B(KEYINPUT54), .ZN(n697) );
  XNOR2_X1 U765 ( .A(KEYINPUT55), .B(KEYINPUT80), .ZN(n696) );
  XNOR2_X1 U766 ( .A(n697), .B(n696), .ZN(n698) );
  XOR2_X1 U767 ( .A(G101), .B(n702), .Z(G3) );
  XOR2_X1 U768 ( .A(n587), .B(KEYINPUT107), .Z(n705) );
  NAND2_X1 U769 ( .A1(n703), .A2(n718), .ZN(n704) );
  XNOR2_X1 U770 ( .A(n705), .B(n704), .ZN(G6) );
  XOR2_X1 U771 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n707) );
  XNOR2_X1 U772 ( .A(G107), .B(KEYINPUT26), .ZN(n706) );
  XNOR2_X1 U773 ( .A(n707), .B(n706), .ZN(n708) );
  XOR2_X1 U774 ( .A(KEYINPUT108), .B(n708), .Z(n710) );
  NAND2_X1 U775 ( .A1(n703), .A2(n720), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n710), .B(n709), .ZN(G9) );
  XOR2_X1 U777 ( .A(G110), .B(n711), .Z(n712) );
  XNOR2_X1 U778 ( .A(KEYINPUT110), .B(n712), .ZN(G12) );
  XOR2_X1 U779 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n714) );
  NAND2_X1 U780 ( .A1(n716), .A2(n720), .ZN(n713) );
  XNOR2_X1 U781 ( .A(n714), .B(n713), .ZN(n715) );
  XOR2_X1 U782 ( .A(G128), .B(n715), .Z(G30) );
  NAND2_X1 U783 ( .A1(n716), .A2(n718), .ZN(n717) );
  XNOR2_X1 U784 ( .A(n717), .B(G146), .ZN(G48) );
  NAND2_X1 U785 ( .A1(n721), .A2(n718), .ZN(n719) );
  XNOR2_X1 U786 ( .A(n719), .B(G113), .ZN(G15) );
  NAND2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U788 ( .A(n722), .B(G116), .ZN(G18) );
  XOR2_X1 U789 ( .A(KEYINPUT37), .B(KEYINPUT113), .Z(n725) );
  XNOR2_X1 U790 ( .A(G125), .B(n723), .ZN(n724) );
  XNOR2_X1 U791 ( .A(n725), .B(n724), .ZN(G27) );
  XNOR2_X1 U792 ( .A(G140), .B(n726), .ZN(G42) );
  NOR2_X1 U793 ( .A1(n727), .A2(n375), .ZN(n728) );
  XNOR2_X1 U794 ( .A(KEYINPUT50), .B(n728), .ZN(n735) );
  XOR2_X1 U795 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n731) );
  NAND2_X1 U796 ( .A1(n496), .A2(n729), .ZN(n730) );
  XNOR2_X1 U797 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U798 ( .A1(n732), .A2(n376), .ZN(n733) );
  XOR2_X1 U799 ( .A(KEYINPUT116), .B(n733), .Z(n734) );
  NOR2_X1 U800 ( .A1(n735), .A2(n734), .ZN(n737) );
  NOR2_X1 U801 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U802 ( .A(KEYINPUT51), .B(n738), .Z(n739) );
  NOR2_X1 U803 ( .A1(n757), .A2(n739), .ZN(n751) );
  NAND2_X1 U804 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U805 ( .A1(n743), .A2(n742), .ZN(n747) );
  NAND2_X1 U806 ( .A1(n745), .A2(n744), .ZN(n746) );
  AND2_X1 U807 ( .A1(n747), .A2(n746), .ZN(n749) );
  BUF_X1 U808 ( .A(n748), .Z(n758) );
  NOR2_X1 U809 ( .A1(n749), .A2(n758), .ZN(n750) );
  NOR2_X1 U810 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U811 ( .A(KEYINPUT52), .B(n752), .ZN(n755) );
  NAND2_X1 U812 ( .A1(G952), .A2(n753), .ZN(n754) );
  NOR2_X1 U813 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U814 ( .A1(G953), .A2(n756), .ZN(n761) );
  NOR2_X1 U815 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U816 ( .A(n759), .B(KEYINPUT117), .ZN(n760) );
  NAND2_X1 U817 ( .A1(n761), .A2(n760), .ZN(n766) );
  INV_X1 U818 ( .A(n434), .ZN(n763) );
  NOR2_X1 U819 ( .A1(n684), .A2(n763), .ZN(n764) );
  NOR2_X1 U820 ( .A1(n766), .A2(n363), .ZN(n767) );
  XNOR2_X1 U821 ( .A(KEYINPUT53), .B(n767), .ZN(G75) );
  XNOR2_X1 U822 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n770) );
  XNOR2_X1 U823 ( .A(n768), .B(KEYINPUT57), .ZN(n769) );
  XNOR2_X1 U824 ( .A(n770), .B(n769), .ZN(n772) );
  NAND2_X1 U825 ( .A1(n774), .A2(G469), .ZN(n771) );
  XOR2_X1 U826 ( .A(n772), .B(n771), .Z(n773) );
  NOR2_X1 U827 ( .A1(n777), .A2(n773), .ZN(G54) );
  INV_X1 U828 ( .A(n775), .ZN(n776) );
  NAND2_X1 U829 ( .A1(G224), .A2(G953), .ZN(n778) );
  XNOR2_X1 U830 ( .A(n778), .B(KEYINPUT61), .ZN(n779) );
  XNOR2_X1 U831 ( .A(KEYINPUT122), .B(n779), .ZN(n780) );
  NAND2_X1 U832 ( .A1(G898), .A2(n780), .ZN(n783) );
  NAND2_X1 U833 ( .A1(n434), .A2(n795), .ZN(n782) );
  NAND2_X1 U834 ( .A1(n783), .A2(n782), .ZN(n790) );
  XNOR2_X1 U835 ( .A(n433), .B(n785), .ZN(n786) );
  NOR2_X1 U836 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U837 ( .A(KEYINPUT123), .B(n788), .Z(n789) );
  XNOR2_X1 U838 ( .A(n790), .B(n789), .ZN(G69) );
  XNOR2_X1 U839 ( .A(n791), .B(KEYINPUT124), .ZN(n792) );
  XOR2_X1 U840 ( .A(n428), .B(n792), .Z(n797) );
  XNOR2_X1 U841 ( .A(n797), .B(KEYINPUT125), .ZN(n794) );
  XNOR2_X1 U842 ( .A(n762), .B(n794), .ZN(n796) );
  NAND2_X1 U843 ( .A1(n796), .A2(n795), .ZN(n802) );
  XNOR2_X1 U844 ( .A(G227), .B(n797), .ZN(n798) );
  XNOR2_X1 U845 ( .A(n798), .B(KEYINPUT126), .ZN(n799) );
  NAND2_X1 U846 ( .A1(n799), .A2(G900), .ZN(n800) );
  NAND2_X1 U847 ( .A1(n800), .A2(G953), .ZN(n801) );
  NAND2_X1 U848 ( .A1(n802), .A2(n801), .ZN(G72) );
  XNOR2_X1 U849 ( .A(G122), .B(KEYINPUT127), .ZN(n805) );
  BUF_X1 U850 ( .A(n803), .Z(n804) );
  XNOR2_X1 U851 ( .A(n805), .B(n804), .ZN(G24) );
  XOR2_X1 U852 ( .A(n429), .B(G119), .Z(G21) );
endmodule

