//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n467), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(KEYINPUT3), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(G137), .A3(new_n466), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n478));
  OAI21_X1  g053(.A(G101), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n471), .B1(new_n480), .B2(new_n464), .ZN(G160));
  INV_X1    g056(.A(new_n466), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n477), .A2(new_n478), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(KEYINPUT3), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT71), .ZN(new_n488));
  INV_X1    g063(.A(G100), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n489), .A2(new_n464), .A3(KEYINPUT72), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT72), .B1(new_n489), .B2(new_n464), .ZN(new_n491));
  OAI221_X1 g066(.A(G2104), .B1(G112), .B2(new_n464), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n485), .A2(new_n464), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n488), .A2(new_n492), .A3(new_n494), .ZN(G162));
  AND2_X1   g070(.A1(new_n466), .A2(new_n468), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(new_n497), .A3(G138), .A4(new_n464), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n475), .A2(G138), .A3(new_n464), .A4(new_n466), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n497), .B1(new_n500), .B2(KEYINPUT75), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT75), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n484), .A2(new_n502), .A3(G138), .A4(new_n464), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n475), .A2(G126), .A3(new_n466), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(KEYINPUT73), .B2(G114), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT73), .A2(G114), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n464), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n464), .A2(G102), .A3(G2104), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n505), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n509), .B1(new_n484), .B2(G126), .ZN(new_n515));
  OAI211_X1 g090(.A(KEYINPUT74), .B(new_n512), .C1(new_n515), .C2(new_n464), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n504), .B1(new_n514), .B2(new_n516), .ZN(G164));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT76), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT6), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n518), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT77), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT78), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n521), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT5), .B(G543), .Z(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT5), .B(G543), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT76), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT76), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g109(.A(KEYINPUT78), .B(new_n530), .C1(new_n534), .C2(new_n521), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G88), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n530), .A2(G62), .ZN(new_n539));
  NAND2_X1  g114(.A1(G75), .A2(G543), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT79), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n519), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n525), .A2(new_n538), .A3(new_n542), .ZN(G303));
  INV_X1    g118(.A(G303), .ZN(G166));
  NAND2_X1  g119(.A1(new_n523), .A2(G51), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT80), .B(KEYINPUT7), .ZN(new_n546));
  AND3_X1   g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  AND2_X1   g124(.A1(G63), .A2(G651), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n548), .A2(new_n549), .B1(new_n530), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n529), .A2(G89), .A3(new_n535), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(G286));
  INV_X1    g129(.A(G286), .ZN(G168));
  NAND3_X1  g130(.A1(new_n529), .A2(G90), .A3(new_n535), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT81), .B(G52), .Z(new_n557));
  NAND2_X1  g132(.A1(G77), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G64), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n528), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n523), .A2(new_n557), .B1(new_n560), .B2(new_n519), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT82), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n556), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(G171));
  NAND3_X1  g141(.A1(new_n529), .A2(G81), .A3(new_n535), .ZN(new_n567));
  NAND2_X1  g142(.A1(G68), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G56), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n528), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n523), .A2(G43), .B1(new_n570), .B2(new_n519), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT83), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n567), .A2(new_n571), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT83), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G860), .ZN(G153));
  NAND4_X1  g154(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g155(.A1(G1), .A2(G3), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT8), .ZN(new_n582));
  NAND4_X1  g157(.A1(G319), .A2(G483), .A3(G661), .A4(new_n582), .ZN(G188));
  XNOR2_X1  g158(.A(new_n530), .B(KEYINPUT85), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  INV_X1    g160(.A(G78), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n584), .A2(new_n585), .B1(new_n586), .B2(new_n518), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT84), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(KEYINPUT9), .ZN(new_n589));
  INV_X1    g164(.A(G53), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n588), .B2(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n523), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n587), .A2(G651), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n529), .A2(G91), .A3(new_n535), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n523), .B(new_n591), .C1(new_n588), .C2(KEYINPUT9), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(G299));
  INV_X1    g172(.A(G171), .ZN(G301));
  NAND3_X1  g173(.A1(new_n529), .A2(G87), .A3(new_n535), .ZN(new_n599));
  INV_X1    g174(.A(G651), .ZN(new_n600));
  INV_X1    g175(.A(G74), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n528), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n523), .B2(G49), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G288));
  NAND3_X1  g179(.A1(new_n529), .A2(G86), .A3(new_n535), .ZN(new_n605));
  NAND2_X1  g180(.A1(G73), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G61), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n528), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n523), .A2(G48), .B1(new_n608), .B2(new_n519), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(G305));
  NAND2_X1  g185(.A1(G72), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G60), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n528), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n523), .A2(G47), .B1(new_n613), .B2(new_n519), .ZN(new_n614));
  INV_X1    g189(.A(G85), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n536), .B2(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n584), .B2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n600), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n528), .A2(KEYINPUT85), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n530), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n625), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(KEYINPUT86), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n621), .A2(new_n627), .B1(G54), .B2(new_n523), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n630));
  INV_X1    g205(.A(G92), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n536), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  MUX2_X1   g210(.A(G301), .B(new_n634), .S(new_n635), .Z(G284));
  MUX2_X1   g211(.A(G301), .B(new_n634), .S(new_n635), .Z(G321));
  NAND2_X1  g212(.A1(G286), .A2(G868), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n585), .B1(new_n622), .B2(new_n624), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n586), .A2(new_n518), .ZN(new_n640));
  OAI21_X1  g215(.A(G651), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n592), .A2(new_n589), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(new_n642), .A3(new_n596), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n643), .A2(new_n594), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n638), .B1(new_n644), .B2(G868), .ZN(G297));
  OAI21_X1  g220(.A(new_n638), .B1(new_n644), .B2(G868), .ZN(G280));
  INV_X1    g221(.A(new_n634), .ZN(new_n647));
  INV_X1    g222(.A(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n648), .B2(G860), .ZN(G148));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n648), .A3(G868), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n578), .A2(new_n635), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT11), .Z(G282));
  INV_X1    g228(.A(new_n652), .ZN(G323));
  NOR2_X1   g229(.A1(new_n483), .A2(G2105), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(new_n496), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT12), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT13), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n486), .A2(G135), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n493), .A2(G123), .ZN(new_n661));
  NOR2_X1   g236(.A1(G99), .A2(G2105), .ZN(new_n662));
  OAI21_X1  g237(.A(G2104), .B1(new_n464), .B2(G111), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n666), .ZN(G156));
  XOR2_X1   g242(.A(G2451), .B(G2454), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1341), .B(G1348), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2427), .B(G2438), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2430), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT15), .B(G2435), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n678), .A3(KEYINPUT14), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n673), .A2(new_n680), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n681), .A2(new_n682), .A3(G14), .ZN(G401));
  XOR2_X1   g258(.A(G2084), .B(G2090), .Z(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n684), .ZN(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(KEYINPUT87), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT17), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n684), .B2(new_n685), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(KEYINPUT17), .ZN(new_n693));
  OAI221_X1 g268(.A(new_n686), .B1(new_n685), .B2(new_n689), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n686), .A2(new_n688), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT18), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(new_n665), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G2100), .ZN(G227));
  XNOR2_X1  g274(.A(G1956), .B(G2474), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1961), .B(G1966), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G1971), .B(G1976), .Z(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT19), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(KEYINPUT19), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n700), .A2(new_n701), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n702), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n704), .A2(KEYINPUT89), .A3(new_n705), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n707), .A2(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n706), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT20), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(G1981), .B(G1986), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT91), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT90), .ZN(new_n721));
  XOR2_X1   g296(.A(G1991), .B(G1996), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n719), .B(new_n723), .ZN(G229));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G23), .ZN(new_n726));
  NAND2_X1  g301(.A1(G288), .A2(KEYINPUT94), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT94), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n599), .A2(new_n728), .A3(new_n603), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n726), .B1(new_n730), .B2(new_n725), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT33), .Z(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(G1976), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(G1976), .ZN(new_n734));
  NOR2_X1   g309(.A1(G6), .A2(G16), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n605), .A2(new_n609), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT32), .ZN(new_n738));
  INV_X1    g313(.A(G1981), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G16), .A2(G22), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G166), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1971), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n733), .A2(new_n734), .A3(new_n740), .A4(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(KEYINPUT34), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n486), .A2(G131), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT92), .ZN(new_n749));
  OR2_X1    g324(.A1(G95), .A2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G107), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n467), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n493), .A2(G119), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  MUX2_X1   g329(.A(G25), .B(new_n754), .S(G29), .Z(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT93), .Z(new_n756));
  XOR2_X1   g331(.A(KEYINPUT35), .B(G1991), .Z(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n756), .A2(new_n758), .ZN(new_n760));
  MUX2_X1   g335(.A(G24), .B(G290), .S(G16), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1986), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n746), .A2(new_n747), .A3(new_n759), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT36), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n725), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1956), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n647), .A2(new_n725), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G4), .B2(new_n725), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G29), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G35), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G162), .B2(new_n776), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT29), .Z(new_n779));
  INV_X1    g354(.A(G2090), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n725), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n725), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n771), .B(new_n781), .C1(G1961), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G164), .A2(new_n776), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G27), .B2(new_n776), .ZN(new_n786));
  INV_X1    g361(.A(G2078), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n773), .B2(new_n774), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n788), .B(new_n790), .C1(new_n780), .C2(new_n779), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n725), .A2(G19), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n578), .B2(new_n725), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT95), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1341), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n776), .A2(G32), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n486), .A2(G141), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n493), .A2(G129), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT26), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n655), .A2(G105), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n797), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT99), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n796), .B1(new_n805), .B2(new_n776), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G1961), .B2(new_n783), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n776), .A2(G33), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n496), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n464), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT97), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT25), .Z(new_n815));
  AOI211_X1 g390(.A(new_n812), .B(new_n815), .C1(G139), .C2(new_n486), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(new_n776), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT98), .B(G2072), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT100), .B(G28), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(KEYINPUT30), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT101), .ZN(new_n822));
  AOI21_X1  g397(.A(G29), .B1(new_n820), .B2(KEYINPUT30), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT31), .B(G11), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n824), .B(new_n825), .C1(new_n664), .C2(new_n776), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT102), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n725), .A2(G21), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G168), .B2(new_n725), .ZN(new_n829));
  INV_X1    g404(.A(G1966), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n819), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n776), .A2(G26), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT28), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n486), .A2(G140), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n493), .A2(G128), .ZN(new_n836));
  NOR2_X1   g411(.A1(G104), .A2(G2105), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n834), .B1(new_n839), .B2(G29), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT96), .B(G2067), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT24), .ZN(new_n843));
  INV_X1    g418(.A(G34), .ZN(new_n844));
  AOI21_X1  g419(.A(G29), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G160), .B2(new_n776), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G2084), .ZN(new_n848));
  NOR4_X1   g423(.A1(new_n809), .A2(new_n832), .A3(new_n842), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n784), .A2(new_n791), .A3(new_n795), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n766), .A2(new_n850), .ZN(G311));
  INV_X1    g426(.A(G311), .ZN(G150));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  INV_X1    g428(.A(G67), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n528), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n519), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n523), .A2(G55), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n856), .B(new_n857), .C1(new_n536), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n647), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n573), .A2(new_n576), .A3(new_n859), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n856), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n537), .B2(G93), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n867), .A3(new_n574), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT103), .B1(new_n572), .B2(new_n859), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n863), .B(new_n870), .Z(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  INV_X1    g448(.A(G860), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n872), .B2(KEYINPUT39), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n861), .B1(new_n873), .B2(new_n875), .ZN(G145));
  NAND2_X1  g451(.A1(new_n805), .A2(new_n816), .ZN(new_n877));
  INV_X1    g452(.A(new_n804), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n816), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n754), .B(new_n657), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n506), .A2(new_n510), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G2105), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n512), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n501), .A2(new_n503), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n498), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n839), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n486), .A2(G142), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n493), .A2(G130), .ZN(new_n891));
  NOR2_X1   g466(.A1(G106), .A2(G2105), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n890), .B(new_n891), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n889), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n881), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n664), .B(G160), .ZN(new_n897));
  XNOR2_X1  g472(.A(G162), .B(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n898), .B2(new_n896), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g476(.A1(new_n859), .A2(new_n635), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n647), .A2(new_n648), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n870), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n629), .A2(new_n632), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n523), .A2(G54), .ZN(new_n907));
  OAI21_X1  g482(.A(G651), .B1(new_n626), .B2(KEYINPUT86), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n619), .A2(new_n620), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(G299), .B(new_n905), .C1(new_n906), .C2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n905), .B1(new_n643), .B2(new_n594), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n593), .A2(new_n595), .A3(KEYINPUT104), .A4(new_n596), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n628), .A4(new_n633), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n911), .A2(new_n914), .A3(KEYINPUT41), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n904), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n915), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n904), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT42), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n924));
  XNOR2_X1  g499(.A(G305), .B(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(G303), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n730), .B(G290), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n926), .B(new_n927), .Z(new_n928));
  XNOR2_X1  g503(.A(new_n923), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n902), .B1(new_n929), .B2(new_n635), .ZN(G295));
  OAI21_X1  g505(.A(new_n902), .B1(new_n929), .B2(new_n635), .ZN(G331));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n868), .A2(new_n869), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n563), .A2(G286), .A3(KEYINPUT107), .A4(new_n565), .ZN(new_n935));
  NAND2_X1  g510(.A1(G286), .A2(KEYINPUT107), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n552), .A2(new_n937), .A3(new_n553), .ZN(new_n938));
  NAND3_X1  g513(.A1(G171), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n934), .A2(new_n864), .A3(new_n935), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n935), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n870), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n917), .A2(new_n918), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n921), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n928), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n926), .B(new_n927), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(new_n945), .A3(new_n943), .ZN(new_n950));
  AND4_X1   g525(.A1(new_n933), .A2(new_n947), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G37), .B1(new_n946), .B2(new_n928), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n933), .B1(new_n952), .B2(new_n950), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT106), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n951), .B2(new_n953), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n932), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT44), .B1(new_n954), .B2(KEYINPUT108), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT109), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n932), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n952), .A2(new_n950), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n952), .A2(new_n933), .A3(new_n950), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT108), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(KEYINPUT108), .B2(new_n954), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n961), .B(new_n962), .C1(new_n967), .C2(new_n932), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n960), .A2(new_n968), .ZN(G397));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n736), .A2(new_n970), .A3(new_n739), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT115), .B1(G305), .B2(G1981), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT118), .Z(new_n974));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(G160), .B2(G40), .ZN(new_n976));
  AOI21_X1  g551(.A(G2105), .B1(new_n476), .B2(new_n479), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR4_X1   g553(.A1(new_n977), .A2(KEYINPUT110), .A3(new_n978), .A4(new_n471), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n504), .B2(new_n884), .ZN(new_n982));
  OAI21_X1  g557(.A(G8), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n970), .B1(new_n736), .B2(new_n739), .ZN(new_n984));
  NOR3_X1   g559(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT116), .B1(G305), .B2(G1981), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n987), .B(new_n739), .C1(new_n605), .C2(new_n609), .ZN(new_n988));
  OAI22_X1  g563(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT49), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n973), .B(KEYINPUT49), .C1(new_n986), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT117), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n995), .A3(new_n992), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(G288), .A2(G1976), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n974), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n480), .A2(new_n464), .ZN(new_n1000));
  INV_X1    g575(.A(new_n471), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(G40), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT110), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G160), .A2(new_n975), .A3(G40), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT45), .B(new_n981), .C1(new_n504), .C2(new_n884), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n516), .A2(new_n514), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n1007), .B2(new_n887), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1005), .B(new_n1006), .C1(new_n1008), .C2(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n743), .ZN(new_n1010));
  AOI21_X1  g585(.A(G2090), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1012), .B(new_n981), .C1(new_n504), .C2(new_n884), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1011), .B(new_n1013), .C1(new_n1008), .C2(new_n1012), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT112), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n1013), .A4(new_n1011), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1010), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT113), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G303), .A2(G8), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n1021), .B(KEYINPUT55), .Z(new_n1022));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1010), .A2(new_n1015), .A3(new_n1023), .A4(new_n1018), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1020), .A2(G8), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  OAI221_X1 g600(.A(new_n981), .B1(new_n504), .B2(new_n884), .C1(new_n976), .C2(new_n979), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n727), .A2(G1976), .A3(new_n729), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1026), .A2(G8), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G8), .ZN(new_n1033));
  INV_X1    g608(.A(new_n982), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(new_n1005), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1035), .A2(KEYINPUT114), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1027), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1032), .A2(new_n1036), .B1(KEYINPUT52), .B2(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n991), .A2(new_n995), .A3(new_n992), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n995), .B1(new_n991), .B2(new_n992), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n999), .A2(new_n983), .B1(new_n1025), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n644), .B(KEYINPUT57), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(G164), .B2(G1384), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1005), .A3(new_n1006), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n980), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1956), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1045), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1005), .B(new_n1013), .C1(new_n1008), .C2(new_n1012), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n774), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1026), .A2(G2067), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n647), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT74), .B1(new_n883), .B2(new_n512), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n511), .A2(new_n505), .A3(new_n513), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n887), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n1012), .A3(new_n981), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(new_n1005), .A3(new_n1052), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n770), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1065), .A2(new_n1044), .A3(new_n1049), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1054), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1044), .A3(new_n1049), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1054), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1068), .B1(new_n1070), .B2(KEYINPUT120), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n1072));
  AOI211_X1 g647(.A(new_n1072), .B(KEYINPUT61), .C1(new_n1054), .C2(new_n1069), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1056), .A2(new_n634), .A3(new_n1057), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1059), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT60), .ZN(new_n1077));
  INV_X1    g652(.A(G1996), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1047), .A2(new_n1078), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1026), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT59), .B1(new_n1082), .B2(new_n578), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1084), .B(new_n577), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n634), .A2(KEYINPUT60), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1056), .A2(new_n1057), .A3(new_n1086), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1077), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1067), .B1(new_n1074), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1047), .A2(new_n787), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  AOI21_X1  g667(.A(G171), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1961), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1055), .A2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g670(.A1(G164), .A2(new_n1046), .A3(G1384), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n982), .A2(new_n1046), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1092), .A2(G2078), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1097), .A2(new_n1005), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1093), .A2(new_n1095), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(KEYINPUT53), .B(G40), .C1(KEYINPUT123), .C2(G2078), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1103), .B1(KEYINPUT123), .B2(G2078), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1001), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(KEYINPUT122), .B2(new_n977), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(KEYINPUT122), .B2(new_n977), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1046), .B2(new_n982), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1055), .A2(new_n1094), .B1(new_n1108), .B2(new_n1006), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1110));
  AOI21_X1  g685(.A(G301), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n1102), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n1100), .A3(new_n1095), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1093), .A2(new_n1109), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1010), .B1(G2090), .B2(new_n1064), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1022), .B1(G8), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1041), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1098), .A2(new_n1005), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n830), .B1(new_n1122), .B2(new_n1096), .ZN(new_n1123));
  INV_X1    g698(.A(G2084), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1016), .A2(new_n1124), .A3(new_n1005), .A4(new_n1013), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(G8), .ZN(new_n1127));
  NAND2_X1  g702(.A1(G286), .A2(G8), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT121), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(KEYINPUT51), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1129), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1126), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1033), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(new_n1131), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1118), .A2(new_n1025), .A3(new_n1121), .A4(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1043), .B1(new_n1090), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1134), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n997), .A2(new_n1139), .A3(new_n1038), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1025), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1033), .B1(new_n1019), .B2(KEYINPUT113), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1022), .B1(new_n1142), .B2(new_n1024), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1140), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1037), .A2(KEYINPUT52), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n994), .B2(new_n996), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1119), .A2(G8), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1022), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1127), .A2(G286), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1148), .A2(new_n1025), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n1153), .B2(KEYINPUT119), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1121), .A2(new_n1155), .A3(new_n1025), .A4(new_n1152), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1144), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT124), .B1(new_n1138), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(KEYINPUT119), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1144), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI221_X4 g738(.A(KEYINPUT54), .B1(new_n1093), .B2(new_n1109), .C1(new_n1113), .C2(G171), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(G171), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1115), .B1(new_n1166), .B2(new_n1101), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1136), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1148), .A2(new_n1025), .A3(new_n1151), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1044), .B1(new_n1065), .B2(new_n1049), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT120), .B1(new_n1066), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT61), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1070), .A2(KEYINPUT120), .A3(new_n1068), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1173), .A2(new_n1174), .A3(new_n1077), .A4(new_n1088), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1067), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1042), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1163), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1136), .A2(KEYINPUT62), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT125), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1169), .A2(new_n1114), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1182), .B(new_n1183), .C1(KEYINPUT62), .C2(new_n1136), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1158), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1098), .A2(new_n980), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n839), .B(G2067), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT111), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n878), .A2(new_n1078), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1189), .B1(new_n805), .B2(new_n1078), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n754), .B(new_n757), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(G290), .B(G1986), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1186), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1185), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1186), .A2(KEYINPUT46), .A3(new_n1078), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT46), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1186), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(G1996), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1188), .A2(new_n878), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1197), .B(new_n1200), .C1(new_n1201), .C2(new_n1199), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT126), .Z(new_n1203));
  OR2_X1    g778(.A1(new_n1203), .A2(KEYINPUT47), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1203), .A2(KEYINPUT47), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1191), .A2(new_n757), .A3(new_n749), .A4(new_n753), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n839), .A2(G2067), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1199), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(G290), .A2(G1986), .ZN(new_n1209));
  AOI21_X1  g784(.A(KEYINPUT48), .B1(new_n1186), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1210), .B1(new_n1193), .B2(new_n1186), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1186), .A2(KEYINPUT48), .A3(new_n1209), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1208), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AND3_X1   g788(.A1(new_n1204), .A2(new_n1205), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1196), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g790(.A1(G227), .A2(new_n462), .ZN(new_n1217));
  XNOR2_X1  g791(.A(new_n1217), .B(KEYINPUT127), .ZN(new_n1218));
  NOR3_X1   g792(.A1(new_n1218), .A2(G401), .A3(G229), .ZN(new_n1219));
  OAI211_X1 g793(.A(new_n1219), .B(new_n900), .C1(new_n953), .C2(new_n951), .ZN(G225));
  INV_X1    g794(.A(G225), .ZN(G308));
endmodule


