

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U551 ( .A(n536), .Z(n518) );
  NAND2_X1 U552 ( .A1(G8), .A2(n681), .ZN(n714) );
  NOR2_X1 U553 ( .A1(G2104), .A2(n521), .ZN(n536) );
  INV_X1 U554 ( .A(n681), .ZN(n661) );
  NAND2_X1 U555 ( .A1(n729), .A2(n727), .ZN(n681) );
  BUF_X1 U556 ( .A(n543), .Z(n527) );
  INV_X1 U557 ( .A(n990), .ZN(n647) );
  INV_X1 U558 ( .A(KEYINPUT96), .ZN(n613) );
  XNOR2_X1 U559 ( .A(n625), .B(n624), .ZN(n674) );
  INV_X1 U560 ( .A(n531), .ZN(n891) );
  XOR2_X1 U561 ( .A(KEYINPUT30), .B(n618), .Z(n519) );
  NOR2_X1 U562 ( .A1(n714), .A2(n700), .ZN(n520) );
  INV_X1 U563 ( .A(KEYINPUT31), .ZN(n624) );
  XNOR2_X1 U564 ( .A(n614), .B(n613), .ZN(n617) );
  INV_X1 U565 ( .A(KEYINPUT17), .ZN(n528) );
  XNOR2_X1 U566 ( .A(n528), .B(KEYINPUT68), .ZN(n529) );
  XNOR2_X1 U567 ( .A(n530), .B(n529), .ZN(n537) );
  AND2_X2 U568 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  INV_X1 U569 ( .A(KEYINPUT108), .ZN(n772) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n799) );
  XNOR2_X1 U571 ( .A(n772), .B(KEYINPUT40), .ZN(n773) );
  INV_X1 U572 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U573 ( .A1(n536), .A2(G126), .ZN(n522) );
  XOR2_X1 U574 ( .A(KEYINPUT87), .B(n522), .Z(n524) );
  NAND2_X1 U575 ( .A1(n895), .A2(G114), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U577 ( .A(KEYINPUT88), .B(n525), .ZN(n535) );
  NAND2_X1 U578 ( .A1(n521), .A2(G2104), .ZN(n526) );
  XNOR2_X1 U579 ( .A(n526), .B(KEYINPUT65), .ZN(n543) );
  NAND2_X1 U580 ( .A1(n527), .A2(G102), .ZN(n533) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  INV_X1 U582 ( .A(n537), .ZN(n531) );
  NAND2_X1 U583 ( .A1(G138), .A2(n891), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U585 ( .A1(n535), .A2(n534), .ZN(G164) );
  NAND2_X1 U586 ( .A1(G125), .A2(n518), .ZN(n539) );
  NAND2_X1 U587 ( .A1(G137), .A2(n537), .ZN(n538) );
  NAND2_X1 U588 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U589 ( .A1(G113), .A2(n895), .ZN(n540) );
  XNOR2_X1 U590 ( .A(KEYINPUT67), .B(n540), .ZN(n541) );
  NOR2_X1 U591 ( .A1(n542), .A2(n541), .ZN(n550) );
  XOR2_X1 U592 ( .A(KEYINPUT23), .B(KEYINPUT66), .Z(n545) );
  NAND2_X1 U593 ( .A1(G101), .A2(n543), .ZN(n544) );
  XNOR2_X1 U594 ( .A(n545), .B(n544), .ZN(n548) );
  NAND2_X1 U595 ( .A1(n550), .A2(n548), .ZN(n547) );
  INV_X1 U596 ( .A(KEYINPUT64), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n547), .A2(n546), .ZN(n552) );
  AND2_X1 U598 ( .A1(n548), .A2(KEYINPUT64), .ZN(n549) );
  NAND2_X1 U599 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U600 ( .A1(n552), .A2(n551), .ZN(G160) );
  XOR2_X1 U601 ( .A(KEYINPUT0), .B(G543), .Z(n594) );
  NOR2_X2 U602 ( .A1(G651), .A2(n594), .ZN(n803) );
  NAND2_X1 U603 ( .A1(n803), .A2(G51), .ZN(n553) );
  XNOR2_X1 U604 ( .A(n553), .B(KEYINPUT76), .ZN(n556) );
  INV_X1 U605 ( .A(G651), .ZN(n559) );
  NOR2_X1 U606 ( .A1(G543), .A2(n559), .ZN(n554) );
  XOR2_X1 U607 ( .A(KEYINPUT1), .B(n554), .Z(n800) );
  NAND2_X1 U608 ( .A1(G63), .A2(n800), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U610 ( .A(KEYINPUT6), .B(n557), .ZN(n565) );
  NAND2_X1 U611 ( .A1(n799), .A2(G89), .ZN(n558) );
  XNOR2_X1 U612 ( .A(n558), .B(KEYINPUT4), .ZN(n562) );
  OR2_X1 U613 ( .A1(n559), .A2(n594), .ZN(n560) );
  XNOR2_X1 U614 ( .A(KEYINPUT69), .B(n560), .ZN(n798) );
  NAND2_X1 U615 ( .A1(G76), .A2(n798), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U617 ( .A(n563), .B(KEYINPUT5), .Z(n564) );
  NOR2_X1 U618 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U619 ( .A(KEYINPUT77), .B(n566), .Z(n567) );
  XOR2_X1 U620 ( .A(KEYINPUT7), .B(n567), .Z(G168) );
  NAND2_X1 U621 ( .A1(G52), .A2(n803), .ZN(n569) );
  NAND2_X1 U622 ( .A1(G64), .A2(n800), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n569), .A2(n568), .ZN(n576) );
  XNOR2_X1 U624 ( .A(KEYINPUT72), .B(KEYINPUT9), .ZN(n574) );
  NAND2_X1 U625 ( .A1(n799), .A2(G90), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n798), .A2(G77), .ZN(n570) );
  XOR2_X1 U627 ( .A(KEYINPUT71), .B(n570), .Z(n571) );
  NAND2_X1 U628 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U629 ( .A(n574), .B(n573), .Z(n575) );
  NOR2_X1 U630 ( .A1(n576), .A2(n575), .ZN(G171) );
  NAND2_X1 U631 ( .A1(G91), .A2(n799), .ZN(n578) );
  NAND2_X1 U632 ( .A1(G78), .A2(n798), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U634 ( .A(KEYINPUT74), .B(n579), .Z(n583) );
  NAND2_X1 U635 ( .A1(n803), .A2(G53), .ZN(n581) );
  NAND2_X1 U636 ( .A1(G65), .A2(n800), .ZN(n580) );
  AND2_X1 U637 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n583), .A2(n582), .ZN(G299) );
  NAND2_X1 U639 ( .A1(G50), .A2(n803), .ZN(n585) );
  NAND2_X1 U640 ( .A1(G62), .A2(n800), .ZN(n584) );
  NAND2_X1 U641 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U642 ( .A(KEYINPUT83), .B(n586), .ZN(n590) );
  NAND2_X1 U643 ( .A1(G88), .A2(n799), .ZN(n588) );
  NAND2_X1 U644 ( .A1(G75), .A2(n798), .ZN(n587) );
  AND2_X1 U645 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U646 ( .A1(n590), .A2(n589), .ZN(G303) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U648 ( .A1(G49), .A2(n803), .ZN(n592) );
  NAND2_X1 U649 ( .A1(G74), .A2(G651), .ZN(n591) );
  NAND2_X1 U650 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U651 ( .A1(n800), .A2(n593), .ZN(n596) );
  NAND2_X1 U652 ( .A1(n594), .A2(G87), .ZN(n595) );
  NAND2_X1 U653 ( .A1(n596), .A2(n595), .ZN(G288) );
  NAND2_X1 U654 ( .A1(G61), .A2(n800), .ZN(n603) );
  NAND2_X1 U655 ( .A1(G86), .A2(n799), .ZN(n598) );
  NAND2_X1 U656 ( .A1(G48), .A2(n803), .ZN(n597) );
  NAND2_X1 U657 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U658 ( .A1(n798), .A2(G73), .ZN(n599) );
  XOR2_X1 U659 ( .A(KEYINPUT2), .B(n599), .Z(n600) );
  NOR2_X1 U660 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U661 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U662 ( .A(n604), .B(KEYINPUT82), .ZN(G305) );
  NAND2_X1 U663 ( .A1(G47), .A2(n803), .ZN(n606) );
  NAND2_X1 U664 ( .A1(G60), .A2(n800), .ZN(n605) );
  NAND2_X1 U665 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U666 ( .A1(G72), .A2(n798), .ZN(n607) );
  XOR2_X1 U667 ( .A(KEYINPUT70), .B(n607), .Z(n608) );
  NOR2_X1 U668 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U669 ( .A1(n799), .A2(G85), .ZN(n610) );
  NAND2_X1 U670 ( .A1(n611), .A2(n610), .ZN(G290) );
  NOR2_X1 U671 ( .A1(G164), .A2(G1384), .ZN(n729) );
  NAND2_X1 U672 ( .A1(G160), .A2(G40), .ZN(n612) );
  XNOR2_X1 U673 ( .A(n612), .B(KEYINPUT89), .ZN(n727) );
  NOR2_X1 U674 ( .A1(n714), .A2(G1966), .ZN(n614) );
  INV_X1 U675 ( .A(n617), .ZN(n676) );
  INV_X1 U676 ( .A(G8), .ZN(n615) );
  NOR2_X1 U677 ( .A1(G2084), .A2(n681), .ZN(n678) );
  NOR2_X1 U678 ( .A1(n615), .A2(n678), .ZN(n616) );
  AND2_X1 U679 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U680 ( .A1(G168), .A2(n519), .ZN(n623) );
  XOR2_X1 U681 ( .A(G2078), .B(KEYINPUT25), .Z(n1011) );
  NOR2_X1 U682 ( .A1(n1011), .A2(n681), .ZN(n619) );
  XNOR2_X1 U683 ( .A(n619), .B(KEYINPUT97), .ZN(n621) );
  OR2_X1 U684 ( .A1(G1961), .A2(n661), .ZN(n620) );
  NAND2_X1 U685 ( .A1(n621), .A2(n620), .ZN(n626) );
  NOR2_X1 U686 ( .A1(G171), .A2(n626), .ZN(n622) );
  NOR2_X1 U687 ( .A1(n623), .A2(n622), .ZN(n625) );
  AND2_X1 U688 ( .A1(n626), .A2(G171), .ZN(n672) );
  AND2_X1 U689 ( .A1(n661), .A2(G1996), .ZN(n627) );
  XOR2_X1 U690 ( .A(KEYINPUT26), .B(n627), .Z(n629) );
  NAND2_X1 U691 ( .A1(n681), .A2(G1341), .ZN(n628) );
  AND2_X1 U692 ( .A1(n629), .A2(n628), .ZN(n651) );
  NAND2_X1 U693 ( .A1(G56), .A2(n800), .ZN(n630) );
  XOR2_X1 U694 ( .A(KEYINPUT14), .B(n630), .Z(n636) );
  NAND2_X1 U695 ( .A1(n799), .A2(G81), .ZN(n631) );
  XNOR2_X1 U696 ( .A(n631), .B(KEYINPUT12), .ZN(n633) );
  NAND2_X1 U697 ( .A1(G68), .A2(n798), .ZN(n632) );
  NAND2_X1 U698 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U699 ( .A(KEYINPUT13), .B(n634), .Z(n635) );
  NOR2_X1 U700 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U701 ( .A1(n803), .A2(G43), .ZN(n637) );
  NAND2_X1 U702 ( .A1(n638), .A2(n637), .ZN(n995) );
  INV_X1 U703 ( .A(n995), .ZN(n649) );
  NAND2_X1 U704 ( .A1(n651), .A2(n649), .ZN(n648) );
  NAND2_X1 U705 ( .A1(G79), .A2(n798), .ZN(n645) );
  NAND2_X1 U706 ( .A1(G92), .A2(n799), .ZN(n640) );
  NAND2_X1 U707 ( .A1(G66), .A2(n800), .ZN(n639) );
  NAND2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U709 ( .A1(G54), .A2(n803), .ZN(n641) );
  XNOR2_X1 U710 ( .A(KEYINPUT75), .B(n641), .ZN(n642) );
  NOR2_X1 U711 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U712 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n646), .B(KEYINPUT15), .ZN(n990) );
  NAND2_X1 U714 ( .A1(n648), .A2(n647), .ZN(n659) );
  AND2_X1 U715 ( .A1(n649), .A2(n990), .ZN(n650) );
  NAND2_X1 U716 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U717 ( .A1(G2067), .A2(n661), .ZN(n652) );
  XOR2_X1 U718 ( .A(KEYINPUT99), .B(n652), .Z(n654) );
  NAND2_X1 U719 ( .A1(G1348), .A2(n681), .ZN(n653) );
  NAND2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U721 ( .A(KEYINPUT100), .B(n655), .ZN(n656) );
  NAND2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n665) );
  NAND2_X1 U724 ( .A1(n661), .A2(G2072), .ZN(n660) );
  XNOR2_X1 U725 ( .A(n660), .B(KEYINPUT27), .ZN(n663) );
  XOR2_X1 U726 ( .A(KEYINPUT98), .B(G1956), .Z(n927) );
  NOR2_X1 U727 ( .A1(n661), .A2(n927), .ZN(n662) );
  NOR2_X1 U728 ( .A1(n663), .A2(n662), .ZN(n666) );
  INV_X1 U729 ( .A(G299), .ZN(n989) );
  NAND2_X1 U730 ( .A1(n666), .A2(n989), .ZN(n664) );
  NAND2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n669) );
  NOR2_X1 U732 ( .A1(n666), .A2(n989), .ZN(n667) );
  XOR2_X1 U733 ( .A(n667), .B(KEYINPUT28), .Z(n668) );
  NAND2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U735 ( .A(KEYINPUT29), .B(n670), .ZN(n671) );
  OR2_X2 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n685) );
  XNOR2_X1 U738 ( .A(n685), .B(KEYINPUT101), .ZN(n675) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n677), .B(KEYINPUT102), .ZN(n680) );
  NAND2_X1 U741 ( .A1(n678), .A2(G8), .ZN(n679) );
  NAND2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n691) );
  NOR2_X1 U743 ( .A1(G1971), .A2(n714), .ZN(n683) );
  NOR2_X1 U744 ( .A1(G2090), .A2(n681), .ZN(n682) );
  NOR2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U746 ( .A1(n684), .A2(G303), .ZN(n687) );
  NAND2_X1 U747 ( .A1(G286), .A2(n685), .ZN(n686) );
  NAND2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U749 ( .A1(G8), .A2(n688), .ZN(n689) );
  XNOR2_X1 U750 ( .A(n689), .B(KEYINPUT32), .ZN(n690) );
  NAND2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n708) );
  NOR2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n693) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n692) );
  NOR2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n997) );
  XOR2_X1 U755 ( .A(G1981), .B(G305), .Z(n983) );
  INV_X1 U756 ( .A(n983), .ZN(n696) );
  NAND2_X1 U757 ( .A1(n693), .A2(KEYINPUT33), .ZN(n694) );
  NOR2_X1 U758 ( .A1(n714), .A2(n694), .ZN(n695) );
  OR2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n700) );
  INV_X1 U760 ( .A(n700), .ZN(n697) );
  AND2_X1 U761 ( .A1(n697), .A2(KEYINPUT33), .ZN(n703) );
  INV_X1 U762 ( .A(n703), .ZN(n698) );
  AND2_X1 U763 ( .A1(n997), .A2(n698), .ZN(n699) );
  NAND2_X1 U764 ( .A1(n708), .A2(n699), .ZN(n705) );
  NAND2_X1 U765 ( .A1(G288), .A2(G1976), .ZN(n701) );
  XOR2_X1 U766 ( .A(KEYINPUT103), .B(n701), .Z(n994) );
  AND2_X1 U767 ( .A1(n520), .A2(n994), .ZN(n702) );
  OR2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U769 ( .A1(n705), .A2(n704), .ZN(n711) );
  NOR2_X1 U770 ( .A1(G2090), .A2(G303), .ZN(n706) );
  NAND2_X1 U771 ( .A1(G8), .A2(n706), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n709), .A2(n714), .ZN(n710) );
  NAND2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n716) );
  NOR2_X1 U775 ( .A1(G1981), .A2(G305), .ZN(n712) );
  XOR2_X1 U776 ( .A(n712), .B(KEYINPUT24), .Z(n713) );
  NOR2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n752) );
  XOR2_X1 U779 ( .A(KEYINPUT37), .B(G2067), .Z(n756) );
  NAND2_X1 U780 ( .A1(G128), .A2(n518), .ZN(n718) );
  NAND2_X1 U781 ( .A1(G116), .A2(n895), .ZN(n717) );
  NAND2_X1 U782 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U783 ( .A(n719), .B(KEYINPUT35), .ZN(n724) );
  NAND2_X1 U784 ( .A1(n527), .A2(G104), .ZN(n721) );
  NAND2_X1 U785 ( .A1(G140), .A2(n891), .ZN(n720) );
  NAND2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U787 ( .A(KEYINPUT34), .B(n722), .Z(n723) );
  NAND2_X1 U788 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U789 ( .A(n725), .B(KEYINPUT36), .ZN(n913) );
  NAND2_X1 U790 ( .A1(n756), .A2(n913), .ZN(n726) );
  XNOR2_X1 U791 ( .A(n726), .B(KEYINPUT91), .ZN(n976) );
  INV_X1 U792 ( .A(n727), .ZN(n728) );
  NOR2_X1 U793 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U794 ( .A(KEYINPUT90), .B(n730), .Z(n768) );
  INV_X1 U795 ( .A(n768), .ZN(n750) );
  AND2_X1 U796 ( .A1(n976), .A2(n750), .ZN(n765) );
  NAND2_X1 U797 ( .A1(G119), .A2(n518), .ZN(n732) );
  NAND2_X1 U798 ( .A1(G107), .A2(n895), .ZN(n731) );
  NAND2_X1 U799 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U800 ( .A(KEYINPUT92), .B(n733), .Z(n737) );
  NAND2_X1 U801 ( .A1(n891), .A2(G131), .ZN(n735) );
  NAND2_X1 U802 ( .A1(n527), .A2(G95), .ZN(n734) );
  AND2_X1 U803 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U804 ( .A1(n737), .A2(n736), .ZN(n905) );
  NAND2_X1 U805 ( .A1(n905), .A2(G1991), .ZN(n748) );
  NAND2_X1 U806 ( .A1(n527), .A2(G105), .ZN(n739) );
  XNOR2_X1 U807 ( .A(KEYINPUT94), .B(KEYINPUT38), .ZN(n738) );
  XNOR2_X1 U808 ( .A(n739), .B(n738), .ZN(n746) );
  NAND2_X1 U809 ( .A1(G129), .A2(n518), .ZN(n741) );
  NAND2_X1 U810 ( .A1(G141), .A2(n891), .ZN(n740) );
  NAND2_X1 U811 ( .A1(n741), .A2(n740), .ZN(n744) );
  NAND2_X1 U812 ( .A1(G117), .A2(n895), .ZN(n742) );
  XNOR2_X1 U813 ( .A(KEYINPUT93), .B(n742), .ZN(n743) );
  NOR2_X1 U814 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U815 ( .A1(n746), .A2(n745), .ZN(n910) );
  NAND2_X1 U816 ( .A1(G1996), .A2(n910), .ZN(n747) );
  NAND2_X1 U817 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U818 ( .A(n749), .B(KEYINPUT95), .Z(n955) );
  AND2_X1 U819 ( .A1(n750), .A2(n955), .ZN(n760) );
  OR2_X1 U820 ( .A1(n765), .A2(n760), .ZN(n751) );
  OR2_X1 U821 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U822 ( .A(n753), .B(KEYINPUT104), .ZN(n755) );
  XOR2_X1 U823 ( .A(G1986), .B(G290), .Z(n1001) );
  NOR2_X1 U824 ( .A1(n1001), .A2(n768), .ZN(n754) );
  NOR2_X1 U825 ( .A1(n755), .A2(n754), .ZN(n771) );
  NOR2_X1 U826 ( .A1(n913), .A2(n756), .ZN(n956) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n910), .ZN(n963) );
  NOR2_X1 U828 ( .A1(G1986), .A2(G290), .ZN(n758) );
  NOR2_X1 U829 ( .A1(G1991), .A2(n905), .ZN(n757) );
  XOR2_X1 U830 ( .A(KEYINPUT105), .B(n757), .Z(n968) );
  NOR2_X1 U831 ( .A1(n758), .A2(n968), .ZN(n759) );
  NOR2_X1 U832 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U833 ( .A(n761), .B(KEYINPUT106), .ZN(n762) );
  NOR2_X1 U834 ( .A1(n963), .A2(n762), .ZN(n763) );
  XOR2_X1 U835 ( .A(KEYINPUT39), .B(n763), .Z(n764) );
  NOR2_X1 U836 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U837 ( .A1(n956), .A2(n766), .ZN(n767) );
  NOR2_X1 U838 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U839 ( .A(KEYINPUT107), .B(n769), .Z(n770) );
  NOR2_X1 U840 ( .A1(n771), .A2(n770), .ZN(n774) );
  XNOR2_X1 U841 ( .A(n774), .B(n773), .ZN(G329) );
  INV_X1 U842 ( .A(G132), .ZN(G219) );
  INV_X1 U843 ( .A(G82), .ZN(G220) );
  INV_X1 U844 ( .A(G120), .ZN(G236) );
  NAND2_X1 U845 ( .A1(G94), .A2(G452), .ZN(n775) );
  XNOR2_X1 U846 ( .A(n775), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n776) );
  XNOR2_X1 U848 ( .A(n776), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U849 ( .A(G223), .ZN(n845) );
  NAND2_X1 U850 ( .A1(n845), .A2(G567), .ZN(n777) );
  XOR2_X1 U851 ( .A(KEYINPUT11), .B(n777), .Z(G234) );
  INV_X1 U852 ( .A(G860), .ZN(n853) );
  OR2_X1 U853 ( .A1(n995), .A2(n853), .ZN(G153) );
  INV_X1 U854 ( .A(G171), .ZN(G301) );
  NAND2_X1 U855 ( .A1(G868), .A2(G301), .ZN(n779) );
  OR2_X1 U856 ( .A1(n990), .A2(G868), .ZN(n778) );
  NAND2_X1 U857 ( .A1(n779), .A2(n778), .ZN(G284) );
  INV_X1 U858 ( .A(G868), .ZN(n817) );
  NOR2_X1 U859 ( .A1(G286), .A2(n817), .ZN(n781) );
  NOR2_X1 U860 ( .A1(G868), .A2(G299), .ZN(n780) );
  NOR2_X1 U861 ( .A1(n781), .A2(n780), .ZN(G297) );
  NAND2_X1 U862 ( .A1(n853), .A2(G559), .ZN(n782) );
  NAND2_X1 U863 ( .A1(n782), .A2(n990), .ZN(n783) );
  XNOR2_X1 U864 ( .A(n783), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U865 ( .A1(n990), .A2(G868), .ZN(n784) );
  NOR2_X1 U866 ( .A1(G559), .A2(n784), .ZN(n785) );
  XNOR2_X1 U867 ( .A(n785), .B(KEYINPUT78), .ZN(n787) );
  NOR2_X1 U868 ( .A1(n995), .A2(G868), .ZN(n786) );
  NOR2_X1 U869 ( .A1(n787), .A2(n786), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G111), .A2(n895), .ZN(n789) );
  NAND2_X1 U871 ( .A1(G135), .A2(n891), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U873 ( .A1(n518), .A2(G123), .ZN(n790) );
  XOR2_X1 U874 ( .A(KEYINPUT18), .B(n790), .Z(n791) );
  NOR2_X1 U875 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U876 ( .A1(n527), .A2(G99), .ZN(n793) );
  NAND2_X1 U877 ( .A1(n794), .A2(n793), .ZN(n969) );
  XOR2_X1 U878 ( .A(n969), .B(G2096), .Z(n796) );
  XNOR2_X1 U879 ( .A(G2100), .B(KEYINPUT79), .ZN(n795) );
  NAND2_X1 U880 ( .A1(n796), .A2(n795), .ZN(G156) );
  INV_X1 U881 ( .A(G303), .ZN(G166) );
  NAND2_X1 U882 ( .A1(G559), .A2(n990), .ZN(n797) );
  XOR2_X1 U883 ( .A(n995), .B(n797), .Z(n852) );
  XNOR2_X1 U884 ( .A(n989), .B(G305), .ZN(n815) );
  NAND2_X1 U885 ( .A1(G80), .A2(n798), .ZN(n808) );
  NAND2_X1 U886 ( .A1(G93), .A2(n799), .ZN(n802) );
  NAND2_X1 U887 ( .A1(G67), .A2(n800), .ZN(n801) );
  NAND2_X1 U888 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U889 ( .A1(n803), .A2(G55), .ZN(n804) );
  XOR2_X1 U890 ( .A(KEYINPUT80), .B(n804), .Z(n805) );
  NOR2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n807) );
  NAND2_X1 U892 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U893 ( .A(n809), .B(KEYINPUT81), .Z(n854) );
  XOR2_X1 U894 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n810) );
  XNOR2_X1 U895 ( .A(G288), .B(n810), .ZN(n811) );
  XOR2_X1 U896 ( .A(n854), .B(n811), .Z(n813) );
  XNOR2_X1 U897 ( .A(G290), .B(G166), .ZN(n812) );
  XNOR2_X1 U898 ( .A(n813), .B(n812), .ZN(n814) );
  XNOR2_X1 U899 ( .A(n815), .B(n814), .ZN(n916) );
  XNOR2_X1 U900 ( .A(n852), .B(n916), .ZN(n816) );
  NAND2_X1 U901 ( .A1(n816), .A2(G868), .ZN(n819) );
  NAND2_X1 U902 ( .A1(n817), .A2(n854), .ZN(n818) );
  NAND2_X1 U903 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U904 ( .A1(G2084), .A2(G2078), .ZN(n820) );
  XOR2_X1 U905 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U906 ( .A1(G2090), .A2(n821), .ZN(n822) );
  XNOR2_X1 U907 ( .A(KEYINPUT21), .B(n822), .ZN(n823) );
  NAND2_X1 U908 ( .A1(n823), .A2(G2072), .ZN(n824) );
  XOR2_X1 U909 ( .A(KEYINPUT85), .B(n824), .Z(G158) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U911 ( .A1(G69), .A2(G57), .ZN(n825) );
  NOR2_X1 U912 ( .A1(G236), .A2(n825), .ZN(n826) );
  XNOR2_X1 U913 ( .A(KEYINPUT86), .B(n826), .ZN(n827) );
  NAND2_X1 U914 ( .A1(n827), .A2(G108), .ZN(n850) );
  NAND2_X1 U915 ( .A1(n850), .A2(G567), .ZN(n832) );
  NOR2_X1 U916 ( .A1(G220), .A2(G219), .ZN(n828) );
  XOR2_X1 U917 ( .A(KEYINPUT22), .B(n828), .Z(n829) );
  NOR2_X1 U918 ( .A1(G218), .A2(n829), .ZN(n830) );
  NAND2_X1 U919 ( .A1(G96), .A2(n830), .ZN(n851) );
  NAND2_X1 U920 ( .A1(n851), .A2(G2106), .ZN(n831) );
  NAND2_X1 U921 ( .A1(n832), .A2(n831), .ZN(n856) );
  NAND2_X1 U922 ( .A1(G483), .A2(G661), .ZN(n833) );
  NOR2_X1 U923 ( .A1(n856), .A2(n833), .ZN(n849) );
  NAND2_X1 U924 ( .A1(n849), .A2(G36), .ZN(G176) );
  XNOR2_X1 U925 ( .A(G2446), .B(G2451), .ZN(n843) );
  XOR2_X1 U926 ( .A(G2430), .B(KEYINPUT110), .Z(n835) );
  XNOR2_X1 U927 ( .A(G2454), .B(G2435), .ZN(n834) );
  XNOR2_X1 U928 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U929 ( .A(G2438), .B(KEYINPUT109), .Z(n837) );
  XNOR2_X1 U930 ( .A(G1341), .B(G1348), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U932 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U933 ( .A(G2427), .B(G2443), .ZN(n840) );
  XNOR2_X1 U934 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U935 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U936 ( .A1(n844), .A2(G14), .ZN(n921) );
  XNOR2_X1 U937 ( .A(KEYINPUT111), .B(n921), .ZN(G401) );
  NAND2_X1 U938 ( .A1(n845), .A2(G2106), .ZN(n846) );
  XNOR2_X1 U939 ( .A(n846), .B(KEYINPUT112), .ZN(G217) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U941 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U943 ( .A1(n849), .A2(n848), .ZN(G188) );
  XNOR2_X1 U944 ( .A(G69), .B(KEYINPUT113), .ZN(G235) );
  INV_X1 U946 ( .A(G108), .ZN(G238) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  INV_X1 U948 ( .A(G57), .ZN(G237) );
  NOR2_X1 U949 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U950 ( .A(G325), .ZN(G261) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(G145) );
  INV_X1 U953 ( .A(n856), .ZN(G319) );
  XOR2_X1 U954 ( .A(G2096), .B(KEYINPUT43), .Z(n858) );
  XNOR2_X1 U955 ( .A(G2090), .B(KEYINPUT42), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n859), .B(G2678), .Z(n861) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U960 ( .A(KEYINPUT114), .B(G2100), .Z(n863) );
  XNOR2_X1 U961 ( .A(G2084), .B(G2078), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(G227) );
  XOR2_X1 U964 ( .A(G1976), .B(G1971), .Z(n867) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1966), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U967 ( .A(n868), .B(KEYINPUT41), .Z(n870) );
  XNOR2_X1 U968 ( .A(G1991), .B(G1996), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U970 ( .A(G2474), .B(G1981), .Z(n872) );
  XNOR2_X1 U971 ( .A(G1961), .B(G1956), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(G229) );
  NAND2_X1 U974 ( .A1(G124), .A2(n518), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n875), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G112), .A2(n895), .ZN(n876) );
  XOR2_X1 U977 ( .A(KEYINPUT115), .B(n876), .Z(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n527), .A2(G100), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G136), .A2(n891), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(G162) );
  NAND2_X1 U983 ( .A1(n527), .A2(G103), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G139), .A2(n891), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G127), .A2(n518), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G115), .A2(n895), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n957) );
  XNOR2_X1 U991 ( .A(n957), .B(G160), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n890), .B(n969), .ZN(n903) );
  NAND2_X1 U993 ( .A1(n527), .A2(G106), .ZN(n893) );
  NAND2_X1 U994 ( .A1(G142), .A2(n891), .ZN(n892) );
  NAND2_X1 U995 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n894), .B(KEYINPUT45), .ZN(n900) );
  NAND2_X1 U997 ( .A1(G130), .A2(n518), .ZN(n897) );
  NAND2_X1 U998 ( .A1(G118), .A2(n895), .ZN(n896) );
  NAND2_X1 U999 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U1000 ( .A(KEYINPUT116), .B(n898), .Z(n899) );
  NAND2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n901), .B(G162), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n912) );
  XOR2_X1 U1004 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n904) );
  XNOR2_X1 U1005 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1006 ( .A(n906), .B(KEYINPUT48), .Z(n908) );
  XNOR2_X1 U1007 ( .A(G164), .B(KEYINPUT46), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n915), .ZN(G395) );
  XNOR2_X1 U1013 ( .A(n995), .B(n916), .ZN(n918) );
  XNOR2_X1 U1014 ( .A(G171), .B(n990), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n919), .B(G286), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n920), .ZN(G397) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n921), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1025 ( .A(G1966), .B(G21), .ZN(n939) );
  XNOR2_X1 U1026 ( .A(n927), .B(G20), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(KEYINPUT59), .B(G1348), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n928), .B(G4), .ZN(n930) );
  XOR2_X1 U1029 ( .A(G1341), .B(G19), .Z(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1031 ( .A(KEYINPUT125), .B(G1981), .Z(n931) );
  XNOR2_X1 U1032 ( .A(G6), .B(n931), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(n936), .B(KEYINPUT60), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(KEYINPUT126), .B(n937), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n949) );
  XNOR2_X1 U1038 ( .A(G1961), .B(KEYINPUT124), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(n940), .B(G5), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(G1971), .B(G22), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G23), .B(G1976), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n944) );
  XOR2_X1 U1043 ( .A(G1986), .B(G24), .Z(n943) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(KEYINPUT58), .B(n945), .ZN(n946) );
  NOR2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(n950), .B(KEYINPUT61), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(KEYINPUT127), .B(n951), .ZN(n953) );
  INV_X1 U1050 ( .A(G16), .ZN(n952) );
  NAND2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n954), .A2(G11), .ZN(n982) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n974) );
  XNOR2_X1 U1054 ( .A(G164), .B(G2078), .ZN(n960) );
  XOR2_X1 U1055 ( .A(G2072), .B(n957), .Z(n958) );
  XNOR2_X1 U1056 ( .A(KEYINPUT119), .B(n958), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(n961), .B(KEYINPUT50), .ZN(n972) );
  XNOR2_X1 U1059 ( .A(G2084), .B(G160), .ZN(n966) );
  XOR2_X1 U1060 ( .A(G2090), .B(G162), .Z(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1062 ( .A(KEYINPUT51), .B(n964), .Z(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT52), .B(n977), .Z(n978) );
  NOR2_X1 U1070 ( .A1(KEYINPUT55), .A2(n978), .ZN(n980) );
  INV_X1 U1071 ( .A(G29), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n1009) );
  XNOR2_X1 U1074 ( .A(G16), .B(KEYINPUT56), .ZN(n1007) );
  XNOR2_X1 U1075 ( .A(G301), .B(G1961), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n985), .B(KEYINPUT123), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT57), .B(n986), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n1005) );
  XNOR2_X1 U1081 ( .A(n989), .B(G1956), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n990), .B(G1348), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n1003) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n999) );
  XOR2_X1 U1086 ( .A(G1341), .B(n995), .Z(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1093 ( .A1(n1009), .A2(n1008), .ZN(n1032) );
  XOR2_X1 U1094 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n1028) );
  XNOR2_X1 U1095 ( .A(G2090), .B(G35), .ZN(n1023) );
  XOR2_X1 U1096 ( .A(G1991), .B(G25), .Z(n1010) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(G28), .ZN(n1020) );
  XNOR2_X1 U1098 ( .A(G1996), .B(G32), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1011), .B(G27), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT120), .B(n1014), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(G2067), .B(G26), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G33), .B(G2072), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(KEYINPUT53), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(G2084), .B(G34), .Z(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT54), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1028), .B(n1027), .ZN(n1030) );
  XNOR2_X1 U1113 ( .A(KEYINPUT122), .B(G29), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(n1033), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

