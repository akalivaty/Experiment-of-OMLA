//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993, new_n994, new_n995;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G227gat), .ZN(new_n205));
  INV_X1    g004(.A(G233gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G113gat), .B(G120gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  XNOR2_X1  g009(.A(G127gat), .B(G134gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G113gat), .B(G120gat), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(G134gat), .ZN(new_n215));
  INV_X1    g014(.A(G134gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G127gat), .ZN(new_n217));
  OAI22_X1  g016(.A1(new_n213), .A2(KEYINPUT1), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT27), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G183gat), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n221), .B(KEYINPUT67), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT28), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT27), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n221), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n227), .A2(new_n228), .B1(new_n220), .B2(G183gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n234), .A2(new_n224), .A3(new_n225), .A4(new_n231), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  INV_X1    g038(.A(G169gat), .ZN(new_n240));
  INV_X1    g039(.A(G176gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n238), .A2(new_n242), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n233), .A2(new_n235), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT23), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n245), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n247), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n249));
  NAND2_X1  g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G190gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n230), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT64), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n246), .B(new_n248), .C1(new_n254), .C2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n260));
  AND3_X1   g059(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(new_n257), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n230), .B1(new_n222), .B2(new_n223), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n247), .A2(KEYINPUT23), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n265), .A2(new_n246), .A3(new_n237), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n259), .A2(new_n260), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n219), .B1(new_n244), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n266), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n265), .A2(new_n246), .A3(new_n237), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT64), .B1(new_n261), .B2(new_n257), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n252), .A2(new_n249), .B1(new_n230), .B2(new_n255), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n269), .B1(new_n273), .B2(KEYINPUT25), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n212), .A2(new_n218), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n233), .A2(new_n235), .A3(new_n243), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n208), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n204), .B1(new_n278), .B2(KEYINPUT33), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n268), .A2(new_n277), .ZN(new_n283));
  AOI221_X4 g082(.A(new_n280), .B1(KEYINPUT33), .B2(new_n204), .C1(new_n283), .C2(new_n207), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT68), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n244), .A2(new_n267), .A3(new_n219), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n275), .B1(new_n274), .B2(new_n276), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n207), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT33), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n291), .A3(new_n204), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n279), .A2(new_n281), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n286), .B2(new_n287), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n268), .A2(KEYINPUT69), .A3(new_n277), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n208), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT70), .B1(new_n299), .B2(KEYINPUT34), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n283), .A2(KEYINPUT34), .A3(new_n207), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n285), .B(new_n295), .C1(new_n300), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT34), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n207), .B1(new_n283), .B2(new_n296), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(new_n298), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n302), .B1(new_n308), .B2(KEYINPUT70), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n282), .A2(new_n284), .ZN(new_n310));
  INV_X1    g109(.A(new_n300), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G8gat), .B(G36gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G197gat), .B(G204gat), .Z(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT72), .B(G211gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G218gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n318), .B1(new_n323), .B2(KEYINPUT73), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT22), .B1(new_n320), .B2(G218gat), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n325), .B(new_n317), .C1(new_n326), .C2(new_n319), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n244), .B2(new_n267), .ZN(new_n332));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n262), .A2(new_n263), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n272), .A2(new_n271), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT25), .B1(new_n337), .B2(new_n266), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n276), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n333), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n330), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT74), .B1(new_n332), .B2(new_n333), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n329), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n334), .A2(new_n328), .A3(new_n341), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n316), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT30), .B1(new_n346), .B2(KEYINPUT75), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n340), .B1(new_n339), .B2(new_n331), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n333), .B1(new_n274), .B2(new_n276), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT74), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n330), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n328), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n345), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n348), .B(new_n349), .C1(new_n356), .C2(new_n316), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n316), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n347), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(G228gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(G148gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G141gat), .ZN(new_n362));
  INV_X1    g161(.A(G141gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G148gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G155gat), .ZN(new_n366));
  INV_X1    g165(.A(G162gat), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT2), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G155gat), .B(G162gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G155gat), .B(G162gat), .Z(new_n374));
  OAI211_X1 g173(.A(new_n368), .B(new_n365), .C1(new_n374), .C2(new_n370), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n323), .A2(new_n318), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n317), .B1(new_n326), .B2(new_n319), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n331), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n380), .A2(new_n381), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n377), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n376), .A2(new_n383), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n331), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n328), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n360), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n324), .A2(new_n331), .A3(new_n327), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n376), .B1(new_n391), .B2(new_n383), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT79), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n389), .B(new_n360), .C1(new_n392), .C2(KEYINPUT79), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT80), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n392), .A2(KEYINPUT79), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n389), .A2(new_n360), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .A4(new_n393), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n390), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G78gat), .B(G106gat), .Z(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(G22gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  NOR2_X1   g204(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n405), .ZN(new_n407));
  AOI211_X1 g206(.A(new_n407), .B(new_n390), .C1(new_n396), .C2(new_n400), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n373), .A2(KEYINPUT3), .A3(new_n375), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n387), .A2(new_n219), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n376), .B2(new_n275), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n376), .A2(new_n275), .A3(new_n413), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n411), .B(new_n412), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n376), .A2(new_n275), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n219), .A2(new_n375), .A3(new_n373), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n412), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n417), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT77), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n416), .A2(new_n425), .A3(new_n422), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(G85gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT0), .B(G57gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT6), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n432), .B2(new_n428), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n313), .A2(new_n359), .A3(new_n409), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT35), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT35), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n406), .B2(new_n408), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(KEYINPUT82), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n428), .A2(new_n442), .A3(KEYINPUT6), .A4(new_n432), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n440), .B1(new_n434), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n347), .A2(new_n357), .A3(new_n358), .ZN(new_n446));
  OAI22_X1  g245(.A1(new_n304), .A2(new_n300), .B1(new_n284), .B2(new_n282), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n312), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n438), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n285), .A2(new_n295), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n304), .A2(new_n300), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n312), .B(KEYINPUT36), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT71), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT71), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n305), .A2(new_n456), .A3(KEYINPUT36), .A4(new_n312), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT36), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n316), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT29), .B1(new_n274), .B2(new_n276), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n341), .B1(new_n462), .B2(new_n340), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n343), .B1(new_n463), .B2(KEYINPUT74), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n345), .B1(new_n464), .B2(new_n328), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n328), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n463), .B2(new_n329), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT38), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n346), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n466), .B1(new_n354), .B2(new_n355), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT37), .B(new_n345), .C1(new_n464), .C2(new_n328), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n316), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT38), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n444), .A2(new_n471), .A3(new_n434), .A4(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n415), .A2(new_n414), .ZN(new_n477));
  INV_X1    g276(.A(new_n411), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n421), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n479), .B(KEYINPUT39), .C1(new_n421), .C2(new_n420), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(new_n421), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT40), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n432), .B1(KEYINPUT81), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n483), .A2(KEYINPUT81), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n428), .A2(new_n432), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n480), .A2(new_n486), .A3(new_n482), .A4(new_n484), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n446), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n409), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n406), .A2(new_n408), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n434), .A2(new_n435), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(new_n446), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n460), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n451), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT13), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT84), .B(G36gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G29gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n506));
  NOR2_X1   g305(.A1(G29gat), .A2(G36gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT14), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n503), .A2(new_n505), .A3(new_n506), .A4(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G29gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n507), .B(KEYINPUT14), .ZN(new_n513));
  OAI211_X1 g312(.A(KEYINPUT15), .B(new_n504), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT85), .ZN(new_n517));
  INV_X1    g316(.A(G1gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(KEYINPUT85), .A3(G1gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G8gat), .ZN(new_n524));
  INV_X1    g323(.A(G8gat), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n519), .A2(new_n525), .A3(new_n520), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(KEYINPUT87), .A3(new_n526), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n515), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n515), .A3(new_n530), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n500), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n510), .A2(new_n514), .A3(KEYINPUT17), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n535), .B1(new_n539), .B2(new_n527), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n524), .A2(new_n526), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n541), .A2(KEYINPUT86), .A3(new_n538), .A4(new_n537), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n540), .A2(new_n499), .A3(new_n542), .A4(new_n533), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n534), .B1(new_n544), .B2(KEYINPUT18), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G169gat), .B(G197gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT12), .Z(new_n555));
  NAND3_X1  g354(.A1(new_n543), .A2(KEYINPUT88), .A3(new_n546), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n545), .A2(new_n549), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n555), .ZN(new_n558));
  INV_X1    g357(.A(new_n547), .ZN(new_n559));
  INV_X1    g358(.A(new_n500), .ZN(new_n560));
  INV_X1    g359(.A(new_n533), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(new_n531), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n543), .B2(new_n546), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n558), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n498), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n566), .A2(KEYINPUT89), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(KEYINPUT89), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G71gat), .B(G78gat), .Z(new_n570));
  XOR2_X1   g369(.A(G57gat), .B(G64gat), .Z(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT90), .ZN(new_n572));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT9), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n570), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  INV_X1    g376(.A(G71gat), .ZN(new_n578));
  INV_X1    g377(.A(G78gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT9), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n573), .A2(KEYINPUT91), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT91), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n571), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n583), .A3(KEYINPUT92), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT92), .B1(new_n581), .B2(new_n583), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n576), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(new_n214), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(G155gat), .ZN(new_n591));
  XOR2_X1   g390(.A(G183gat), .B(G211gat), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT94), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n591), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n586), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n572), .A2(new_n575), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n597), .A2(new_n584), .B1(new_n598), .B2(new_n570), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n529), .A2(new_n530), .B1(KEYINPUT21), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n596), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT7), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n610));
  NOR2_X1   g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  AOI211_X1 g411(.A(new_n610), .B(new_n611), .C1(KEYINPUT8), .C2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G85gat), .ZN(new_n614));
  INV_X1    g413(.A(G92gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT8), .A2(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(KEYINPUT98), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n609), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G99gat), .B(G106gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n609), .B(new_n619), .C1(new_n613), .C2(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n537), .A2(new_n623), .A3(new_n538), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n626));
  INV_X1    g425(.A(new_n515), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(new_n623), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT99), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n537), .A2(new_n623), .A3(new_n538), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n621), .A2(new_n622), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n515), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n630), .A2(new_n631), .A3(new_n633), .A4(new_n626), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n629), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n629), .B2(new_n634), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n606), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n629), .A2(new_n634), .ZN(new_n639));
  INV_X1    g438(.A(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n629), .A2(new_n634), .A3(new_n635), .ZN(new_n642));
  INV_X1    g441(.A(new_n606), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(G190gat), .B(G218gat), .Z(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  AND3_X1   g446(.A1(new_n638), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n638), .B2(new_n644), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n605), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n620), .A2(KEYINPUT100), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n632), .A2(new_n599), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n623), .B1(new_n587), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n632), .A2(new_n599), .A3(new_n660), .A4(KEYINPUT10), .ZN(new_n661));
  OAI211_X1 g460(.A(KEYINPUT10), .B(new_n576), .C1(new_n585), .C2(new_n586), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT101), .B1(new_n662), .B2(new_n623), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n653), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n653), .B1(new_n655), .B2(new_n657), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n665), .B(new_n671), .C1(new_n670), .C2(new_n669), .ZN(new_n672));
  INV_X1    g471(.A(new_n653), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n661), .A2(new_n663), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n655), .A2(new_n657), .A3(new_n658), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n668), .B1(new_n676), .B2(new_n669), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n652), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n569), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n495), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g482(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n684));
  OAI211_X1 g483(.A(new_n446), .B(new_n679), .C1(new_n567), .C2(new_n568), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n684), .B1(new_n687), .B2(new_n525), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT16), .B(G8gat), .Z(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n681), .A2(KEYINPUT42), .A3(new_n446), .A4(new_n689), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1325gat));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n460), .A2(new_n694), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n454), .A2(KEYINPUT71), .B1(new_n448), .B2(new_n458), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(KEYINPUT105), .A3(new_n457), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(G15gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT106), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n681), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n680), .B2(new_n448), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1326gat));
  NAND2_X1  g505(.A1(new_n681), .A2(new_n494), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  INV_X1    g508(.A(new_n605), .ZN(new_n710));
  INV_X1    g509(.A(new_n678), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n651), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n569), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n495), .A2(new_n511), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT45), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n437), .A2(KEYINPUT35), .B1(new_n445), .B2(new_n449), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n493), .A2(new_n496), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n698), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n648), .B2(new_n649), .ZN(new_n723));
  INV_X1    g522(.A(new_n647), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n636), .A2(new_n637), .A3(new_n606), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n643), .B1(new_n641), .B2(new_n642), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n638), .A2(new_n644), .A3(new_n647), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(KEYINPUT108), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n718), .B1(new_n721), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n498), .A2(KEYINPUT44), .A3(new_n650), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n565), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n712), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n436), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n717), .A2(new_n738), .ZN(G1328gat));
  NAND2_X1  g538(.A1(new_n446), .A2(new_n501), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n714), .A2(KEYINPUT46), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n502), .B1(new_n737), .B2(new_n359), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT46), .B1(new_n714), .B2(new_n740), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n741), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(G1329gat));
  INV_X1    g546(.A(new_n737), .ZN(new_n748));
  INV_X1    g547(.A(new_n698), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n748), .A2(G43gat), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(G43gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n714), .B2(new_n448), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1330gat));
  NAND3_X1  g554(.A1(new_n748), .A2(G50gat), .A3(new_n494), .ZN(new_n756));
  INV_X1    g555(.A(G50gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n714), .B2(new_n409), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g559(.A1(new_n721), .A2(new_n565), .A3(new_n652), .A4(new_n711), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n495), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n446), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT49), .B(G64gat), .Z(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(G1333gat));
  NAND3_X1  g570(.A1(new_n765), .A2(G71gat), .A3(new_n749), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n578), .B1(new_n764), .B2(new_n448), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1334gat));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n409), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(new_n579), .ZN(G1335gat));
  NOR3_X1   g580(.A1(new_n605), .A2(new_n565), .A3(new_n711), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT105), .B1(new_n696), .B2(new_n457), .ZN(new_n783));
  AND4_X1   g582(.A1(KEYINPUT105), .A2(new_n455), .A3(new_n457), .A4(new_n459), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n720), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n731), .B1(new_n785), .B2(new_n451), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n733), .B(new_n782), .C1(new_n786), .C2(KEYINPUT44), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n732), .A2(KEYINPUT113), .A3(new_n733), .A4(new_n782), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n436), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT114), .B1(new_n721), .B2(new_n651), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n605), .A2(new_n565), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n493), .A2(new_n496), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n695), .B2(new_n697), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n795), .B(new_n650), .C1(new_n797), .C2(new_n719), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n793), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT51), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n793), .A2(new_n801), .A3(new_n794), .A4(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n678), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n495), .A2(new_n614), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n792), .B1(new_n803), .B2(new_n804), .ZN(G1336gat));
  NOR2_X1   g604(.A1(new_n359), .A2(G92gat), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n800), .A2(new_n678), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  OAI21_X1  g607(.A(G92gat), .B1(new_n787), .B2(new_n359), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n359), .B1(new_n789), .B2(new_n790), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n615), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n812), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT115), .B1(new_n812), .B2(KEYINPUT52), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(G1337gat));
  OAI21_X1  g614(.A(G99gat), .B1(new_n791), .B2(new_n698), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n448), .A2(G99gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n803), .B2(new_n817), .ZN(G1338gat));
  AOI21_X1  g617(.A(new_n409), .B1(new_n789), .B2(new_n790), .ZN(new_n819));
  XNOR2_X1  g618(.A(KEYINPUT116), .B(G106gat), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n409), .A2(G106gat), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n819), .A2(new_n821), .B1(new_n803), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT53), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n803), .A2(new_n825), .A3(new_n822), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n803), .B2(new_n822), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n734), .A2(new_n494), .A3(new_n782), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT53), .B1(new_n828), .B2(new_n820), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n824), .B1(new_n826), .B2(new_n830), .ZN(G1339gat));
  NOR3_X1   g630(.A1(new_n652), .A2(new_n565), .A3(new_n678), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n540), .A2(new_n542), .A3(new_n533), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(G229gat), .A3(G233gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n532), .A2(new_n533), .A3(new_n500), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n554), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n557), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n668), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n676), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n674), .A2(new_n673), .A3(new_n675), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n843), .A3(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n672), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT55), .B1(new_n841), .B2(new_n843), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n838), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n730), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n557), .A2(new_n678), .A3(new_n837), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n845), .A2(new_n846), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n565), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n730), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n605), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n848), .B(KEYINPUT118), .C1(new_n730), .C2(new_n851), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n832), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n436), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n313), .A2(new_n409), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n446), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(G113gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n565), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n857), .A2(new_n409), .A3(new_n449), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n565), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(new_n862), .ZN(G1340gat));
  AND2_X1   g665(.A1(new_n864), .A2(new_n678), .ZN(new_n867));
  INV_X1    g666(.A(G120gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n678), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT119), .Z(new_n870));
  OAI22_X1  g669(.A1(new_n867), .A2(new_n868), .B1(new_n860), .B2(new_n870), .ZN(G1341gat));
  AOI21_X1  g670(.A(G127gat), .B1(new_n861), .B2(new_n605), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n710), .A2(new_n214), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n864), .B2(new_n873), .ZN(G1342gat));
  NAND3_X1  g673(.A1(new_n861), .A2(new_n216), .A3(new_n650), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n216), .B1(new_n864), .B2(new_n650), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n875), .A2(KEYINPUT56), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n879), .A2(KEYINPUT120), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(KEYINPUT120), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(G1343gat));
  NOR2_X1   g681(.A1(new_n851), .A2(new_n730), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n844), .A2(new_n672), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n841), .A2(new_n843), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT55), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n884), .A2(new_n557), .A3(new_n887), .A4(new_n837), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n729), .B2(new_n723), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n853), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n710), .A3(new_n855), .ZN(new_n891));
  INV_X1    g690(.A(new_n832), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n409), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n698), .A2(new_n495), .A3(new_n359), .ZN(new_n895));
  NOR4_X1   g694(.A1(new_n894), .A2(G141gat), .A3(new_n735), .A4(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(KEYINPUT58), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n846), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n898), .A2(new_n884), .A3(new_n565), .A4(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n849), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n650), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n889), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n904), .A2(new_n605), .ZN(new_n905));
  OAI211_X1 g704(.A(KEYINPUT57), .B(new_n494), .C1(new_n905), .C2(new_n832), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n907));
  INV_X1    g706(.A(new_n895), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G141gat), .B1(new_n909), .B2(new_n735), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n897), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT57), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n912), .B1(new_n856), .B2(new_n409), .ZN(new_n913));
  AOI211_X1 g712(.A(KEYINPUT122), .B(new_n895), .C1(new_n913), .C2(new_n906), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n915), .B1(new_n907), .B2(new_n908), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n565), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n896), .B1(new_n917), .B2(G141gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n911), .B1(new_n918), .B2(new_n919), .ZN(G1344gat));
  NOR2_X1   g719(.A1(new_n894), .A2(new_n895), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n361), .A3(new_n678), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G148gat), .ZN(new_n924));
  INV_X1    g723(.A(new_n916), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n915), .A3(new_n908), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n924), .B1(new_n927), .B2(new_n678), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT57), .B1(new_n856), .B2(new_n409), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n888), .A2(new_n651), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n903), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n710), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n903), .A2(new_n931), .A3(new_n930), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n892), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n912), .A3(new_n494), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n678), .A3(new_n908), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n923), .B1(new_n938), .B2(G148gat), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n922), .B1(new_n928), .B2(new_n939), .ZN(G1345gat));
  AOI21_X1  g739(.A(G155gat), .B1(new_n921), .B2(new_n605), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n710), .A2(new_n366), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n927), .B2(new_n942), .ZN(G1346gat));
  NAND3_X1  g742(.A1(new_n921), .A2(new_n367), .A3(new_n650), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n731), .B1(new_n925), .B2(new_n926), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n367), .ZN(G1347gat));
  NOR3_X1   g745(.A1(new_n856), .A2(new_n495), .A3(new_n359), .ZN(new_n947));
  INV_X1    g746(.A(new_n858), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n240), .A3(new_n565), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n436), .A2(new_n446), .ZN(new_n952));
  NOR4_X1   g751(.A1(new_n856), .A2(new_n448), .A3(new_n494), .A4(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(new_n565), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n240), .B2(new_n954), .ZN(G1348gat));
  AOI21_X1  g754(.A(G176gat), .B1(new_n950), .B2(new_n678), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n711), .A2(new_n241), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n953), .B2(new_n957), .ZN(G1349gat));
  AND2_X1   g757(.A1(new_n953), .A2(new_n605), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n605), .A2(new_n221), .A3(new_n231), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n959), .A2(new_n230), .B1(new_n949), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g761(.A(new_n255), .B1(new_n953), .B2(new_n650), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT61), .Z(new_n964));
  NAND3_X1  g763(.A1(new_n950), .A2(new_n229), .A3(new_n730), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1351gat));
  NOR2_X1   g765(.A1(new_n749), .A2(new_n952), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n893), .A2(new_n967), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n968), .A2(G197gat), .A3(new_n735), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT124), .Z(new_n970));
  NAND2_X1  g769(.A1(new_n937), .A2(new_n967), .ZN(new_n971));
  OAI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n735), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1352gat));
  NOR2_X1   g772(.A1(new_n711), .A2(G204gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n893), .A2(new_n967), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n975), .B(KEYINPUT62), .Z(new_n976));
  NAND4_X1  g775(.A1(new_n929), .A2(new_n936), .A3(new_n678), .A4(new_n967), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(G204gat), .B1(new_n977), .B2(new_n978), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n976), .B(new_n983), .C1(new_n979), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1353gat));
  OR3_X1    g784(.A1(new_n968), .A2(new_n320), .A3(new_n710), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n937), .A2(new_n605), .A3(new_n967), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n987), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  AOI21_X1  g787(.A(KEYINPUT63), .B1(new_n987), .B2(G211gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(G1354gat));
  INV_X1    g789(.A(G218gat), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n971), .A2(new_n991), .A3(new_n651), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n991), .B1(new_n968), .B2(new_n731), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n993), .A2(KEYINPUT127), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n993), .A2(KEYINPUT127), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(G1355gat));
endmodule


