//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT16), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n189), .A3(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(G146), .A3(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT24), .B(G110), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT76), .ZN(new_n202));
  XNOR2_X1  g016(.A(new_n201), .B(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G128), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n205), .B(KEYINPUT75), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n204), .B2(G128), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n213), .A2(new_n205), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n210), .B1(new_n215), .B2(G110), .ZN(new_n216));
  INV_X1    g030(.A(G110), .ZN(new_n217));
  AOI211_X1 g031(.A(KEYINPUT77), .B(new_n217), .C1(new_n211), .C2(new_n214), .ZN(new_n218));
  OAI221_X1 g032(.A(new_n200), .B1(new_n203), .B2(new_n209), .C1(new_n216), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n199), .A2(KEYINPUT78), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n193), .A2(new_n221), .A3(G146), .A4(new_n195), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n190), .A2(new_n192), .A3(new_n197), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n203), .A2(new_n209), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n215), .A2(G110), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n223), .B(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n219), .A2(new_n227), .A3(KEYINPUT79), .ZN(new_n231));
  INV_X1    g045(.A(G953), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(G221), .A3(G234), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n233), .B(KEYINPUT22), .ZN(new_n234));
  INV_X1    g048(.A(G137), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n228), .A2(new_n236), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n188), .B1(new_n240), .B2(KEYINPUT25), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n237), .A2(new_n242), .A3(new_n238), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n237), .A2(new_n239), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n188), .A2(new_n238), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n197), .A2(G143), .ZN(new_n248));
  INV_X1    g062(.A(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(G143), .B2(new_n197), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n207), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  AND4_X1   g073(.A1(new_n255), .A2(new_n258), .A3(new_n248), .A4(new_n250), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n254), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G137), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n235), .A2(KEYINPUT11), .A3(G134), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(G137), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n264), .A2(new_n265), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n263), .A2(G137), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n235), .A2(G134), .ZN(new_n270));
  OAI21_X1  g084(.A(G131), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n248), .A2(new_n250), .A3(KEYINPUT0), .A4(G128), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT0), .B(G128), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n256), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G131), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n268), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n273), .A2(KEYINPUT30), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n258), .A2(new_n248), .A3(new_n250), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT65), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n256), .A2(new_n255), .A3(new_n258), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT1), .B1(new_n249), .B2(G146), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n286), .A2(new_n287), .B1(new_n291), .B2(new_n251), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n268), .A2(new_n271), .A3(KEYINPUT64), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT64), .B1(new_n268), .B2(new_n271), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n281), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G116), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(G119), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT67), .B1(new_n204), .B2(G116), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n298), .A3(G119), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT2), .B(G113), .Z(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n273), .A2(new_n306), .A3(new_n281), .A4(KEYINPUT30), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n283), .A2(new_n297), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n305), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n273), .A3(new_n281), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT26), .B(G101), .ZN(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G210), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n311), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT31), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT31), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n308), .A2(new_n322), .A3(new_n317), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n310), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n305), .B1(new_n295), .B2(new_n296), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n309), .A2(new_n273), .A3(KEYINPUT28), .A4(new_n281), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n316), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n322), .B1(new_n308), .B2(new_n317), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n321), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(G472), .A2(G902), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT71), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  AOI211_X1 g151(.A(KEYINPUT72), .B(KEYINPUT32), .C1(new_n334), .C2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n330), .B(new_n323), .C1(new_n332), .C2(KEYINPUT70), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT32), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n336), .A2(new_n343), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n340), .B2(new_n341), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT74), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n346), .C1(new_n340), .C2(new_n341), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n328), .A2(new_n329), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n308), .A2(new_n310), .ZN(new_n352));
  AOI211_X1 g166(.A(KEYINPUT29), .B(new_n351), .C1(new_n329), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n273), .A2(new_n281), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n305), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT73), .A3(new_n310), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n357), .A3(new_n305), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(KEYINPUT28), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n325), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n316), .A2(KEYINPUT29), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n238), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G472), .B1(new_n353), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n350), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n247), .B1(new_n345), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(G234), .A2(G237), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n367), .A2(G952), .A3(new_n232), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n367), .A2(G902), .A3(G953), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT21), .B(G898), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n373), .A2(KEYINPUT3), .A3(G107), .ZN(new_n374));
  AND2_X1   g188(.A1(KEYINPUT81), .A2(G104), .ZN(new_n375));
  NOR2_X1   g189(.A1(KEYINPUT81), .A2(G104), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n374), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(new_n375), .B2(new_n376), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n300), .A2(new_n302), .ZN(new_n384));
  INV_X1    g198(.A(new_n299), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(KEYINPUT5), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G113), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT5), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n387), .B1(new_n299), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n380), .B1(G104), .B2(new_n379), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G101), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n303), .A2(new_n304), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n383), .A2(new_n390), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n374), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(G104), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(new_n379), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n396), .B2(new_n379), .ZN(new_n399));
  OAI21_X1  g213(.A(G101), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n402), .B(G101), .C1(new_n397), .C2(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n305), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n394), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(G110), .B(G122), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n406), .B(new_n394), .C1(new_n401), .C2(new_n404), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(KEYINPUT6), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n276), .A2(G125), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n261), .B2(G125), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n232), .A2(G224), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n412), .B(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n405), .A2(new_n416), .A3(new_n407), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n410), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT7), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  OAI221_X1 g235(.A(new_n411), .B1(new_n419), .B2(new_n414), .C1(new_n261), .C2(G125), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n406), .B(KEYINPUT8), .ZN(new_n424));
  AND4_X1   g238(.A1(new_n393), .A2(new_n383), .A3(new_n390), .A4(new_n392), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n383), .A2(new_n392), .B1(new_n390), .B2(new_n393), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n409), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n238), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT84), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n431), .A3(new_n238), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n418), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G210), .B1(G237), .B2(G902), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n418), .A2(new_n430), .A3(new_n434), .A4(new_n432), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  OR2_X1    g253(.A1(KEYINPUT91), .A2(G122), .ZN(new_n440));
  NAND2_X1  g254(.A1(KEYINPUT91), .A2(G122), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n298), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n298), .A2(G122), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n379), .A3(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n298), .A2(G122), .ZN(new_n446));
  OAI21_X1  g260(.A(G107), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n207), .A2(G143), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n249), .A2(G128), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT13), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n263), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n452), .A2(new_n454), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n448), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n444), .B(KEYINPUT14), .ZN(new_n458));
  OAI21_X1  g272(.A(G107), .B1(new_n458), .B2(new_n442), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(G134), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n451), .A2(new_n263), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n445), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n457), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT9), .B(G234), .ZN(new_n466));
  INV_X1    g280(.A(G217), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n466), .A2(new_n467), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n463), .A2(new_n445), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n459), .A2(KEYINPUT92), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n460), .B(G107), .C1(new_n458), .C2(new_n442), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n471), .B(new_n462), .C1(new_n472), .C2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n468), .A3(new_n457), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G478), .B1(KEYINPUT93), .B2(KEYINPUT15), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(KEYINPUT93), .B2(KEYINPUT15), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT94), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT94), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AND4_X1   g300(.A1(new_n372), .A2(new_n438), .A3(new_n439), .A4(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT95), .ZN(new_n488));
  OAI21_X1  g302(.A(G221), .B1(new_n466), .B2(G902), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G469), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(new_n238), .ZN(new_n492));
  XNOR2_X1  g306(.A(G110), .B(G140), .ZN(new_n493));
  INV_X1    g307(.A(G227), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(G953), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n493), .B(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n279), .A2(new_n268), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT82), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n403), .A2(new_n277), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n401), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n382), .B1(new_n378), .B2(new_n381), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n276), .B1(new_n501), .B2(new_n402), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT82), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n383), .A2(new_n392), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT10), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n292), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n251), .B1(new_n253), .B2(new_n257), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n259), .B2(new_n260), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n383), .A3(new_n392), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n507), .A2(new_n509), .B1(new_n512), .B2(new_n508), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n497), .B1(new_n505), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT82), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT82), .B1(new_n502), .B2(new_n503), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n497), .B(new_n513), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n496), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n512), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n261), .B1(new_n383), .B2(new_n392), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n280), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT12), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n506), .A2(new_n292), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n512), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT12), .A3(new_n280), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n496), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n517), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(G902), .B1(new_n519), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n492), .B1(new_n531), .B2(new_n491), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n517), .A2(new_n529), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(new_n514), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n496), .B(KEYINPUT80), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(new_n528), .B2(new_n517), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT83), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n535), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT12), .B1(new_n526), .B2(new_n280), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n523), .B(new_n497), .C1(new_n525), .C2(new_n512), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n538), .B1(new_n518), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT83), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n280), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n517), .A3(new_n529), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n537), .A2(G469), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n490), .B1(new_n532), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n191), .A2(G140), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n189), .A2(G125), .ZN(new_n551));
  OAI21_X1  g365(.A(G146), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n224), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n312), .A2(G214), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n249), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n312), .A2(G143), .A3(G214), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(KEYINPUT18), .A2(G131), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n557), .A2(KEYINPUT86), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT86), .B1(new_n557), .B2(new_n559), .ZN(new_n561));
  OAI221_X1 g375(.A(new_n553), .B1(new_n557), .B2(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n198), .A2(new_n199), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n557), .A2(KEYINPUT17), .A3(G131), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n557), .A2(G131), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n555), .A2(new_n266), .A3(new_n556), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n563), .B(new_n564), .C1(new_n567), .C2(KEYINPUT17), .ZN(new_n568));
  XNOR2_X1  g382(.A(G113), .B(G122), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n373), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n562), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n562), .B2(new_n568), .ZN(new_n573));
  OAI211_X1 g387(.A(KEYINPUT90), .B(new_n238), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G475), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n562), .A2(new_n568), .ZN(new_n576));
  INV_X1    g390(.A(new_n570), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(G902), .B1(new_n578), .B2(new_n571), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(KEYINPUT90), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n582));
  OR2_X1    g396(.A1(KEYINPUT87), .A2(KEYINPUT19), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n582), .B(new_n583), .C1(new_n550), .C2(new_n551), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT87), .A4(KEYINPUT19), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n220), .A2(new_n222), .B1(new_n586), .B2(new_n197), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT88), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n567), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n197), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n223), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n562), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT89), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(KEYINPUT89), .B(new_n562), .C1(new_n589), .C2(new_n591), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n577), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n571), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT20), .ZN(new_n598));
  NOR2_X1   g412(.A1(G475), .A2(G902), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n570), .B1(new_n592), .B2(new_n593), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n572), .B1(new_n603), .B2(new_n595), .ZN(new_n604));
  INV_X1    g418(.A(new_n599), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n581), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n487), .A2(new_n488), .A3(new_n549), .A4(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n439), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n436), .B2(new_n437), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(new_n607), .A3(new_n372), .A4(new_n486), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n537), .A2(G469), .A3(new_n547), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n529), .B1(new_n545), .B2(new_n517), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n533), .A2(new_n541), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n491), .B(new_n238), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n492), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n489), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT95), .B1(new_n611), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n366), .A2(new_n608), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  NAND2_X1  g435(.A1(new_n610), .A2(new_n372), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n247), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n334), .A2(new_n238), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n624), .A2(G472), .B1(new_n337), .B2(new_n334), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n549), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  INV_X1    g441(.A(new_n470), .ZN(new_n628));
  INV_X1    g442(.A(new_n476), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n470), .A2(KEYINPUT33), .A3(new_n476), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n630), .A2(G478), .A3(new_n238), .A4(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n477), .A2(G478), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n633), .A2(KEYINPUT96), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(KEYINPUT96), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n600), .A2(new_n606), .ZN(new_n637));
  INV_X1    g451(.A(G475), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n579), .B2(KEYINPUT90), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(KEYINPUT90), .B2(new_n579), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n626), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT97), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n643), .B(new_n645), .ZN(G6));
  AND2_X1   g460(.A1(new_n640), .A2(new_n485), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n597), .A2(new_n599), .A3(new_n601), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n648), .A2(new_n606), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n648), .B2(new_n606), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n626), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND2_X1  g469(.A1(new_n230), .A2(new_n231), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g472(.A(new_n246), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n244), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n625), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n608), .A2(new_n619), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  XNOR2_X1  g479(.A(new_n368), .B(KEYINPUT99), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n668), .B2(new_n369), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n647), .B(new_n670), .C1(new_n650), .C2(new_n651), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n601), .B1(new_n597), .B2(new_n599), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n604), .A2(new_n605), .A3(new_n602), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT98), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n648), .A2(new_n606), .A3(new_n649), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n678), .A2(KEYINPUT100), .A3(new_n647), .A4(new_n670), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n673), .A2(new_n610), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT101), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n673), .A2(new_n679), .A3(new_n682), .A4(new_n610), .ZN(new_n683));
  INV_X1    g497(.A(new_n661), .ZN(new_n684));
  AOI211_X1 g498(.A(new_n684), .B(new_n618), .C1(new_n345), .C2(new_n365), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  XOR2_X1   g501(.A(new_n669), .B(KEYINPUT39), .Z(new_n688));
  NAND2_X1  g502(.A1(new_n549), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT40), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n438), .B(KEYINPUT102), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT38), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n342), .A2(new_n343), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT72), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n342), .A2(new_n339), .A3(new_n343), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n356), .A2(new_n358), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n238), .B1(new_n697), .B2(new_n316), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n329), .B1(new_n308), .B2(new_n310), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n348), .A2(new_n700), .A3(new_n350), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n684), .A2(new_n641), .A3(new_n439), .A4(new_n485), .ZN(new_n703));
  OR4_X1    g517(.A1(new_n690), .A2(new_n692), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT103), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  INV_X1    g520(.A(new_n350), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n349), .B1(new_n334), .B2(new_n346), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n694), .A3(new_n695), .A4(new_n363), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n641), .A2(new_n610), .A3(new_n636), .A4(new_n670), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n710), .A2(new_n549), .A3(new_n661), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  INV_X1    g527(.A(new_n247), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n642), .A2(new_n622), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n613), .A2(new_n614), .ZN(new_n716));
  OAI21_X1  g530(.A(G469), .B1(new_n716), .B2(G902), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n489), .A3(new_n615), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n710), .A2(new_n714), .A3(new_n715), .A4(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT41), .B(G113), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT104), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(G15));
  NOR2_X1   g537(.A1(new_n652), .A2(new_n622), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n710), .A2(new_n714), .A3(new_n724), .A4(new_n719), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NOR2_X1   g540(.A1(new_n611), .A2(new_n718), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n710), .A2(new_n727), .A3(new_n661), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NAND2_X1  g543(.A1(new_n624), .A2(G472), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n316), .B1(new_n359), .B2(new_n325), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT105), .B1(new_n731), .B2(new_n332), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n323), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n731), .A2(KEYINPUT105), .A3(new_n332), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n337), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n247), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n438), .A2(new_n439), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n738), .A2(new_n607), .A3(new_n486), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n372), .A3(new_n719), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  NOR2_X1   g555(.A1(new_n736), .A2(new_n684), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n642), .A2(new_n669), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n718), .A2(new_n738), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT106), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n191), .ZN(G27));
  AOI211_X1 g561(.A(G469), .B(G902), .C1(new_n519), .C2(new_n530), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n542), .A2(G469), .A3(new_n546), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n616), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n489), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n436), .A2(new_n439), .A3(new_n437), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT107), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n752), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n615), .A2(new_n616), .A3(new_n749), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .A4(new_n489), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n363), .A2(new_n347), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n247), .B1(new_n759), .B2(new_n693), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n758), .A2(KEYINPUT42), .A3(new_n743), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n758), .A2(new_n710), .A3(new_n714), .A4(new_n743), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT42), .B1(new_n763), .B2(KEYINPUT108), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n366), .A2(new_n765), .A3(new_n758), .A4(new_n743), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n762), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n266), .ZN(G33));
  AND2_X1   g582(.A1(new_n366), .A2(new_n758), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT109), .B1(new_n673), .B2(new_n679), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n673), .A2(KEYINPUT109), .A3(new_n679), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(KEYINPUT110), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n366), .A3(new_n758), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n775), .B2(new_n770), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NAND2_X1  g592(.A1(new_n636), .A2(new_n607), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT43), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n625), .A3(new_n684), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n752), .B1(new_n781), .B2(KEYINPUT44), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT45), .B1(new_n537), .B2(new_n547), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n542), .A2(KEYINPUT45), .A3(new_n546), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(G469), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n616), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n748), .B1(new_n786), .B2(new_n787), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n490), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(new_n688), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n782), .B(new_n791), .C1(KEYINPUT44), .C2(new_n781), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(KEYINPUT47), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n796), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n364), .A2(new_n338), .A3(new_n344), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n800), .A2(new_n247), .A3(new_n743), .A4(new_n754), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  NAND2_X1  g617(.A1(new_n717), .A2(new_n615), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT49), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n714), .A2(new_n489), .A3(new_n439), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n805), .A2(new_n806), .A3(new_n779), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n692), .A2(new_n807), .A3(new_n702), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n692), .A2(new_n609), .A3(new_n719), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n780), .A2(new_n666), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(new_n737), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n804), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(KEYINPUT114), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(KEYINPUT114), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n816), .A2(new_n817), .A3(new_n489), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n754), .B(new_n811), .C1(new_n799), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n719), .A2(new_n754), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT115), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n821), .A2(new_n810), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n742), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n714), .A2(new_n368), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n702), .A3(new_n824), .ZN(new_n825));
  OR3_X1    g639(.A1(new_n825), .A2(new_n641), .A3(new_n636), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n814), .A2(new_n819), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n763), .A2(KEYINPUT108), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT42), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n766), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n761), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n642), .B1(new_n641), .B2(new_n486), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n623), .A3(new_n549), .A4(new_n625), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n620), .A2(new_n728), .A3(new_n740), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n663), .A2(new_n720), .A3(new_n725), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n752), .A2(new_n581), .A3(new_n485), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n549), .A3(new_n678), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n800), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n730), .A2(new_n735), .A3(new_n641), .A4(new_n636), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n753), .B2(new_n757), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n661), .B(new_n670), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n837), .A2(new_n777), .A3(new_n842), .A4(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n751), .A2(new_n661), .A3(new_n669), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n850), .B(new_n739), .C1(new_n696), .C2(new_n701), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n712), .A2(new_n745), .A3(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n852), .A2(new_n686), .A3(KEYINPUT52), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(new_n852), .B2(new_n686), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n833), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n686), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n852), .A2(new_n686), .A3(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n663), .A2(new_n720), .A3(new_n725), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n728), .A2(new_n740), .A3(new_n839), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n862), .A2(new_n863), .A3(new_n620), .A4(new_n848), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n767), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n861), .A2(new_n865), .A3(new_n866), .A4(new_n777), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT54), .B1(new_n856), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n849), .B2(new_n855), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT112), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT112), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n871), .B(new_n866), .C1(new_n849), .C2(new_n855), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n861), .A2(new_n865), .A3(new_n777), .A4(new_n833), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n868), .B1(new_n874), .B2(KEYINPUT54), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n232), .A2(G952), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n811), .B2(new_n744), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n822), .A2(new_n760), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n878), .A2(KEYINPUT48), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(KEYINPUT48), .ZN(new_n880));
  OAI221_X1 g694(.A(new_n877), .B1(new_n642), .B2(new_n825), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n827), .B2(new_n828), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n831), .A2(new_n875), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n808), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n232), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n856), .A2(new_n867), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n238), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G210), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n410), .A2(new_n417), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n415), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT55), .Z(new_n895));
  OAI21_X1  g709(.A(new_n887), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n895), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n892), .A2(KEYINPUT117), .A3(new_n895), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(G51));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n856), .A2(new_n867), .A3(KEYINPUT54), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n492), .B(KEYINPUT57), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n716), .B(KEYINPUT118), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n783), .A2(new_n785), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n889), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n886), .B1(new_n909), .B2(new_n911), .ZN(G54));
  NAND2_X1  g726(.A1(KEYINPUT58), .A2(G475), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n889), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n604), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n889), .A2(new_n597), .A3(new_n914), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n887), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT119), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n916), .A2(new_n920), .A3(new_n887), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(G60));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n630), .A2(new_n631), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT120), .Z(new_n925));
  XOR2_X1   g739(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n926));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n923), .B1(new_n905), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n856), .A2(KEYINPUT54), .A3(new_n867), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n923), .B(new_n929), .C1(new_n931), .C2(new_n868), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n887), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n925), .B1(new_n875), .B2(new_n928), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT123), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n925), .C1(new_n875), .C2(new_n928), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n934), .B1(new_n936), .B2(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n888), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n658), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n245), .B(KEYINPUT124), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n888), .B2(new_n941), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n887), .A3(new_n945), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT61), .Z(G66));
  INV_X1    g761(.A(new_n842), .ZN(new_n948));
  NAND2_X1  g762(.A1(G224), .A2(G953), .ZN(new_n949));
  OAI22_X1  g763(.A1(new_n948), .A2(G953), .B1(new_n370), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n893), .B1(G898), .B2(new_n232), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT125), .Z(new_n952));
  XNOR2_X1  g766(.A(new_n950), .B(new_n952), .ZN(G69));
  OAI21_X1  g767(.A(G953), .B1(new_n494), .B2(new_n668), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(KEYINPUT126), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n791), .A2(new_n739), .A3(new_n760), .ZN(new_n956));
  AND4_X1   g770(.A1(new_n837), .A2(new_n792), .A3(new_n802), .A4(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n712), .A2(new_n745), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n957), .A2(new_n686), .A3(new_n777), .A4(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(G953), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n283), .A2(new_n297), .A3(new_n307), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n586), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n955), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n954), .A2(KEYINPUT126), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n704), .A2(new_n686), .A3(new_n958), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n689), .A2(new_n752), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n366), .A2(new_n969), .A3(new_n838), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n792), .A2(new_n802), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n232), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n962), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n964), .A2(new_n965), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n965), .B1(new_n964), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G72));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT63), .Z(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n959), .B2(new_n948), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n352), .A2(new_n316), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n983), .B(new_n979), .C1(new_n959), .C2(new_n948), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n979), .B1(new_n972), .B2(new_n948), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n886), .B1(new_n986), .B2(new_n699), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n979), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n982), .A2(new_n699), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n988), .B1(new_n874), .B2(new_n990), .ZN(G57));
endmodule


