

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U567 ( .A(n682), .ZN(n667) );
  NOR2_X4 U568 ( .A1(G651), .A2(n580), .ZN(n819) );
  BUF_X1 U569 ( .A(n733), .Z(n734) );
  XNOR2_X1 U570 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n675) );
  INV_X1 U571 ( .A(KEYINPUT28), .ZN(n661) );
  XNOR2_X1 U572 ( .A(n676), .B(n675), .ZN(n677) );
  AND2_X1 U573 ( .A1(G160), .A2(G40), .ZN(n607) );
  NAND2_X1 U574 ( .A1(G8), .A2(n682), .ZN(n730) );
  AND2_X2 U575 ( .A1(n533), .A2(G2104), .ZN(n912) );
  NOR2_X2 U576 ( .A1(G2104), .A2(n536), .ZN(n909) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n553), .Z(n818) );
  OR2_X1 U578 ( .A1(n786), .A2(n785), .ZN(n787) );
  INV_X1 U579 ( .A(KEYINPUT23), .ZN(n535) );
  INV_X1 U580 ( .A(G2105), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n912), .A2(G101), .ZN(n534) );
  XNOR2_X1 U582 ( .A(n535), .B(n534), .ZN(n538) );
  INV_X1 U583 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U584 ( .A1(n909), .A2(G125), .ZN(n537) );
  NAND2_X1 U585 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U586 ( .A(n539), .B(KEYINPUT64), .ZN(n545) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n540) );
  XOR2_X1 U588 ( .A(KEYINPUT17), .B(n540), .Z(n736) );
  NAND2_X1 U589 ( .A1(G137), .A2(n736), .ZN(n543) );
  NAND2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n541) );
  XNOR2_X1 U591 ( .A(n541), .B(KEYINPUT65), .ZN(n733) );
  NAND2_X1 U592 ( .A1(G113), .A2(n733), .ZN(n542) );
  NAND2_X1 U593 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X2 U594 ( .A1(n545), .A2(n544), .ZN(G160) );
  XOR2_X1 U595 ( .A(KEYINPUT0), .B(G543), .Z(n580) );
  NAND2_X1 U596 ( .A1(G52), .A2(n819), .ZN(n546) );
  XNOR2_X1 U597 ( .A(n546), .B(KEYINPUT67), .ZN(n551) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n822) );
  NAND2_X1 U599 ( .A1(G90), .A2(n822), .ZN(n548) );
  INV_X1 U600 ( .A(G651), .ZN(n552) );
  NOR2_X1 U601 ( .A1(n580), .A2(n552), .ZN(n823) );
  NAND2_X1 U602 ( .A1(G77), .A2(n823), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n555) );
  NOR2_X1 U606 ( .A1(G543), .A2(n552), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n818), .A2(G64), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n555), .A2(n554), .ZN(G301) );
  INV_X1 U609 ( .A(G301), .ZN(G171) );
  NAND2_X1 U610 ( .A1(G63), .A2(n818), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G51), .A2(n819), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U613 ( .A(KEYINPUT6), .B(n558), .ZN(n566) );
  XNOR2_X1 U614 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n564) );
  NAND2_X1 U615 ( .A1(n822), .A2(G89), .ZN(n559) );
  XNOR2_X1 U616 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G76), .A2(n823), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n562), .B(KEYINPUT5), .ZN(n563) );
  XNOR2_X1 U620 ( .A(n564), .B(n563), .ZN(n565) );
  NOR2_X1 U621 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U622 ( .A(KEYINPUT7), .B(KEYINPUT74), .Z(n567) );
  XNOR2_X1 U623 ( .A(n568), .B(n567), .ZN(G168) );
  NAND2_X1 U624 ( .A1(G88), .A2(n822), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G75), .A2(n823), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n576) );
  NAND2_X1 U627 ( .A1(n819), .A2(G50), .ZN(n571) );
  XNOR2_X1 U628 ( .A(n571), .B(KEYINPUT84), .ZN(n573) );
  NAND2_X1 U629 ( .A1(G62), .A2(n818), .ZN(n572) );
  NAND2_X1 U630 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U631 ( .A(KEYINPUT85), .B(n574), .Z(n575) );
  NOR2_X1 U632 ( .A1(n576), .A2(n575), .ZN(G166) );
  XNOR2_X1 U633 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  XOR2_X1 U634 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U635 ( .A1(G49), .A2(n819), .ZN(n578) );
  NAND2_X1 U636 ( .A1(G74), .A2(G651), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U638 ( .A1(n818), .A2(n579), .ZN(n582) );
  NAND2_X1 U639 ( .A1(n580), .A2(G87), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n582), .A2(n581), .ZN(G288) );
  NAND2_X1 U641 ( .A1(n822), .A2(G86), .ZN(n583) );
  XOR2_X1 U642 ( .A(KEYINPUT81), .B(n583), .Z(n585) );
  NAND2_X1 U643 ( .A1(n818), .A2(G61), .ZN(n584) );
  NAND2_X1 U644 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U645 ( .A(KEYINPUT82), .B(n586), .ZN(n590) );
  XOR2_X1 U646 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n588) );
  NAND2_X1 U647 ( .A1(n823), .A2(G73), .ZN(n587) );
  XOR2_X1 U648 ( .A(n588), .B(n587), .Z(n589) );
  NOR2_X1 U649 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U650 ( .A1(n819), .A2(G48), .ZN(n591) );
  NAND2_X1 U651 ( .A1(n592), .A2(n591), .ZN(G305) );
  NAND2_X1 U652 ( .A1(G85), .A2(n822), .ZN(n594) );
  NAND2_X1 U653 ( .A1(G72), .A2(n823), .ZN(n593) );
  NAND2_X1 U654 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U655 ( .A1(G60), .A2(n818), .ZN(n596) );
  NAND2_X1 U656 ( .A1(G47), .A2(n819), .ZN(n595) );
  NAND2_X1 U657 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U658 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U659 ( .A(KEYINPUT66), .B(n599), .Z(G290) );
  NAND2_X1 U660 ( .A1(G102), .A2(n912), .ZN(n601) );
  NAND2_X1 U661 ( .A1(G126), .A2(n909), .ZN(n600) );
  NAND2_X1 U662 ( .A1(n601), .A2(n600), .ZN(n606) );
  NAND2_X1 U663 ( .A1(G114), .A2(n733), .ZN(n602) );
  XNOR2_X1 U664 ( .A(n602), .B(KEYINPUT88), .ZN(n604) );
  NAND2_X1 U665 ( .A1(n736), .A2(G138), .ZN(n603) );
  NAND2_X1 U666 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U667 ( .A1(n606), .A2(n605), .ZN(G164) );
  NOR2_X1 U668 ( .A1(G164), .A2(G1384), .ZN(n755) );
  NAND2_X2 U669 ( .A1(n607), .A2(n755), .ZN(n682) );
  NAND2_X1 U670 ( .A1(G65), .A2(n818), .ZN(n609) );
  NAND2_X1 U671 ( .A1(G53), .A2(n819), .ZN(n608) );
  NAND2_X1 U672 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U673 ( .A1(G91), .A2(n822), .ZN(n611) );
  NAND2_X1 U674 ( .A1(G78), .A2(n823), .ZN(n610) );
  NAND2_X1 U675 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U676 ( .A1(n613), .A2(n612), .ZN(n956) );
  NAND2_X1 U677 ( .A1(G1956), .A2(n682), .ZN(n616) );
  NAND2_X1 U678 ( .A1(n667), .A2(G2072), .ZN(n614) );
  XOR2_X1 U679 ( .A(KEYINPUT27), .B(n614), .Z(n615) );
  NAND2_X1 U680 ( .A1(n616), .A2(n615), .ZN(n618) );
  INV_X1 U681 ( .A(KEYINPUT98), .ZN(n617) );
  XNOR2_X1 U682 ( .A(n618), .B(n617), .ZN(n660) );
  NAND2_X1 U683 ( .A1(n956), .A2(n660), .ZN(n659) );
  NAND2_X1 U684 ( .A1(G92), .A2(n822), .ZN(n620) );
  NAND2_X1 U685 ( .A1(G66), .A2(n818), .ZN(n619) );
  NAND2_X1 U686 ( .A1(n620), .A2(n619), .ZN(n626) );
  NAND2_X1 U687 ( .A1(n819), .A2(G54), .ZN(n621) );
  XNOR2_X1 U688 ( .A(n621), .B(KEYINPUT70), .ZN(n623) );
  NAND2_X1 U689 ( .A1(G79), .A2(n823), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U691 ( .A(KEYINPUT71), .B(n624), .Z(n625) );
  NOR2_X1 U692 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U693 ( .A(KEYINPUT15), .B(n627), .Z(n944) );
  NAND2_X1 U694 ( .A1(G1348), .A2(n682), .ZN(n628) );
  XNOR2_X1 U695 ( .A(KEYINPUT101), .B(n628), .ZN(n631) );
  NAND2_X1 U696 ( .A1(n667), .A2(G2067), .ZN(n629) );
  XOR2_X1 U697 ( .A(KEYINPUT102), .B(n629), .Z(n630) );
  NOR2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  OR2_X1 U699 ( .A1(n944), .A2(n632), .ZN(n657) );
  NAND2_X1 U700 ( .A1(n944), .A2(n632), .ZN(n655) );
  NAND2_X1 U701 ( .A1(n823), .A2(G68), .ZN(n633) );
  XNOR2_X1 U702 ( .A(KEYINPUT68), .B(n633), .ZN(n636) );
  NAND2_X1 U703 ( .A1(n822), .A2(G81), .ZN(n634) );
  XNOR2_X1 U704 ( .A(KEYINPUT12), .B(n634), .ZN(n635) );
  NAND2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n637), .B(KEYINPUT13), .ZN(n639) );
  NAND2_X1 U707 ( .A1(G43), .A2(n819), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U709 ( .A1(n818), .A2(G56), .ZN(n640) );
  XOR2_X1 U710 ( .A(KEYINPUT14), .B(n640), .Z(n641) );
  NOR2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n953) );
  XNOR2_X1 U712 ( .A(KEYINPUT99), .B(G1341), .ZN(n644) );
  AND2_X1 U713 ( .A1(n682), .A2(KEYINPUT26), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n649) );
  INV_X1 U715 ( .A(KEYINPUT99), .ZN(n647) );
  NAND2_X1 U716 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n645) );
  AND2_X1 U717 ( .A1(n645), .A2(n667), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n651) );
  OR2_X1 U720 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U722 ( .A(KEYINPUT100), .B(n652), .Z(n653) );
  NAND2_X1 U723 ( .A1(n953), .A2(n653), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n664) );
  NOR2_X1 U727 ( .A1(n956), .A2(n660), .ZN(n662) );
  XNOR2_X1 U728 ( .A(n662), .B(n661), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U730 ( .A(n665), .B(KEYINPUT29), .ZN(n671) );
  XOR2_X1 U731 ( .A(G2078), .B(KEYINPUT25), .Z(n666) );
  XNOR2_X1 U732 ( .A(KEYINPUT97), .B(n666), .ZN(n1000) );
  NOR2_X1 U733 ( .A1(n682), .A2(n1000), .ZN(n669) );
  XOR2_X1 U734 ( .A(KEYINPUT96), .B(G1961), .Z(n970) );
  NOR2_X1 U735 ( .A1(n667), .A2(n970), .ZN(n668) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n673) );
  AND2_X1 U737 ( .A1(G171), .A2(n673), .ZN(n670) );
  NOR2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(KEYINPUT103), .ZN(n693) );
  NOR2_X1 U740 ( .A1(G171), .A2(n673), .ZN(n679) );
  NOR2_X1 U741 ( .A1(G1966), .A2(n730), .ZN(n696) );
  NOR2_X1 U742 ( .A1(G2084), .A2(n682), .ZN(n695) );
  NOR2_X1 U743 ( .A1(n696), .A2(n695), .ZN(n674) );
  NAND2_X1 U744 ( .A1(G8), .A2(n674), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(G168), .ZN(n678) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n680), .B(KEYINPUT31), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(KEYINPUT105), .ZN(n694) );
  NOR2_X1 U749 ( .A1(G1971), .A2(n730), .ZN(n684) );
  NOR2_X1 U750 ( .A1(G2090), .A2(n682), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n685), .A2(G303), .ZN(n687) );
  AND2_X1 U753 ( .A1(n694), .A2(n687), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n693), .A2(n686), .ZN(n691) );
  INV_X1 U755 ( .A(n687), .ZN(n688) );
  OR2_X1 U756 ( .A1(n688), .A2(G286), .ZN(n689) );
  AND2_X1 U757 ( .A1(G8), .A2(n689), .ZN(n690) );
  NAND2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(KEYINPUT32), .ZN(n701) );
  AND2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n699) );
  AND2_X1 U761 ( .A1(G8), .A2(n695), .ZN(n697) );
  OR2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  OR2_X1 U763 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n716) );
  NOR2_X1 U765 ( .A1(G1976), .A2(G288), .ZN(n705) );
  NOR2_X1 U766 ( .A1(G1971), .A2(G303), .ZN(n702) );
  NOR2_X1 U767 ( .A1(n705), .A2(n702), .ZN(n945) );
  NAND2_X1 U768 ( .A1(n716), .A2(n945), .ZN(n703) );
  XOR2_X1 U769 ( .A(KEYINPUT106), .B(n703), .Z(n704) );
  NOR2_X1 U770 ( .A1(n730), .A2(n704), .ZN(n711) );
  NAND2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n957) );
  INV_X1 U772 ( .A(KEYINPUT33), .ZN(n713) );
  INV_X1 U773 ( .A(n730), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n722), .A2(n705), .ZN(n706) );
  NOR2_X1 U775 ( .A1(n713), .A2(n706), .ZN(n707) );
  XNOR2_X1 U776 ( .A(n707), .B(KEYINPUT107), .ZN(n712) );
  AND2_X1 U777 ( .A1(n957), .A2(n712), .ZN(n709) );
  XNOR2_X1 U778 ( .A(G1981), .B(G305), .ZN(n948) );
  INV_X1 U779 ( .A(n948), .ZN(n708) );
  AND2_X1 U780 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U781 ( .A1(n711), .A2(n710), .ZN(n726) );
  INV_X1 U782 ( .A(n712), .ZN(n714) );
  OR2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U784 ( .A1(n948), .A2(n715), .ZN(n724) );
  INV_X1 U785 ( .A(n716), .ZN(n720) );
  INV_X1 U786 ( .A(G2090), .ZN(n717) );
  NAND2_X1 U787 ( .A1(G8), .A2(n717), .ZN(n718) );
  NOR2_X1 U788 ( .A1(G303), .A2(n718), .ZN(n719) );
  NOR2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U791 ( .A1(n724), .A2(n723), .ZN(n725) );
  AND2_X1 U792 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U793 ( .A(n727), .B(KEYINPUT108), .ZN(n732) );
  NOR2_X1 U794 ( .A1(G1981), .A2(G305), .ZN(n728) );
  XOR2_X1 U795 ( .A(n728), .B(KEYINPUT24), .Z(n729) );
  OR2_X1 U796 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U797 ( .A1(n732), .A2(n731), .ZN(n771) );
  XOR2_X1 U798 ( .A(G1986), .B(G290), .Z(n963) );
  NAND2_X1 U799 ( .A1(G117), .A2(n734), .ZN(n735) );
  XNOR2_X1 U800 ( .A(n735), .B(KEYINPUT94), .ZN(n743) );
  NAND2_X1 U801 ( .A1(G129), .A2(n909), .ZN(n738) );
  BUF_X1 U802 ( .A(n736), .Z(n913) );
  NAND2_X1 U803 ( .A1(G141), .A2(n913), .ZN(n737) );
  NAND2_X1 U804 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U805 ( .A1(n912), .A2(G105), .ZN(n739) );
  XOR2_X1 U806 ( .A(KEYINPUT38), .B(n739), .Z(n740) );
  NOR2_X1 U807 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U808 ( .A1(n743), .A2(n742), .ZN(n894) );
  NAND2_X1 U809 ( .A1(G1996), .A2(n894), .ZN(n744) );
  XOR2_X1 U810 ( .A(KEYINPUT95), .B(n744), .Z(n753) );
  NAND2_X1 U811 ( .A1(G119), .A2(n909), .ZN(n746) );
  NAND2_X1 U812 ( .A1(G107), .A2(n734), .ZN(n745) );
  NAND2_X1 U813 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U814 ( .A(KEYINPUT93), .B(n747), .ZN(n751) );
  NAND2_X1 U815 ( .A1(n912), .A2(G95), .ZN(n749) );
  NAND2_X1 U816 ( .A1(G131), .A2(n913), .ZN(n748) );
  AND2_X1 U817 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U818 ( .A1(n751), .A2(n750), .ZN(n890) );
  NAND2_X1 U819 ( .A1(G1991), .A2(n890), .ZN(n752) );
  NAND2_X1 U820 ( .A1(n753), .A2(n752), .ZN(n775) );
  INV_X1 U821 ( .A(n775), .ZN(n1020) );
  NAND2_X1 U822 ( .A1(n963), .A2(n1020), .ZN(n756) );
  NAND2_X1 U823 ( .A1(G160), .A2(G40), .ZN(n754) );
  NOR2_X1 U824 ( .A1(n755), .A2(n754), .ZN(n783) );
  NAND2_X1 U825 ( .A1(n756), .A2(n783), .ZN(n769) );
  XNOR2_X1 U826 ( .A(KEYINPUT36), .B(KEYINPUT91), .ZN(n767) );
  NAND2_X1 U827 ( .A1(G104), .A2(n912), .ZN(n758) );
  NAND2_X1 U828 ( .A1(G140), .A2(n913), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U830 ( .A(KEYINPUT34), .B(n759), .ZN(n764) );
  NAND2_X1 U831 ( .A1(G128), .A2(n909), .ZN(n761) );
  NAND2_X1 U832 ( .A1(G116), .A2(n734), .ZN(n760) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U834 ( .A(n762), .B(KEYINPUT35), .Z(n763) );
  NOR2_X1 U835 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U836 ( .A(KEYINPUT90), .B(n765), .Z(n766) );
  XNOR2_X1 U837 ( .A(n767), .B(n766), .ZN(n888) );
  XNOR2_X1 U838 ( .A(G2067), .B(KEYINPUT37), .ZN(n780) );
  NOR2_X1 U839 ( .A1(n888), .A2(n780), .ZN(n1022) );
  NAND2_X1 U840 ( .A1(n1022), .A2(n783), .ZN(n768) );
  XNOR2_X1 U841 ( .A(KEYINPUT92), .B(n768), .ZN(n778) );
  NAND2_X1 U842 ( .A1(n769), .A2(n778), .ZN(n770) );
  NOR2_X1 U843 ( .A1(n771), .A2(n770), .ZN(n786) );
  NOR2_X1 U844 ( .A1(G1996), .A2(n894), .ZN(n1031) );
  NOR2_X1 U845 ( .A1(G1986), .A2(G290), .ZN(n772) );
  NOR2_X1 U846 ( .A1(G1991), .A2(n890), .ZN(n1026) );
  NOR2_X1 U847 ( .A1(n772), .A2(n1026), .ZN(n773) );
  XOR2_X1 U848 ( .A(KEYINPUT109), .B(n773), .Z(n774) );
  NOR2_X1 U849 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U850 ( .A1(n1031), .A2(n776), .ZN(n777) );
  XNOR2_X1 U851 ( .A(n777), .B(KEYINPUT39), .ZN(n779) );
  NAND2_X1 U852 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U853 ( .A1(n888), .A2(n780), .ZN(n1019) );
  NAND2_X1 U854 ( .A1(n781), .A2(n1019), .ZN(n782) );
  NAND2_X1 U855 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U856 ( .A(KEYINPUT110), .B(n784), .Z(n785) );
  XNOR2_X1 U857 ( .A(n787), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U858 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U859 ( .A1(G123), .A2(n909), .ZN(n788) );
  XNOR2_X1 U860 ( .A(n788), .B(KEYINPUT18), .ZN(n795) );
  NAND2_X1 U861 ( .A1(G135), .A2(n913), .ZN(n790) );
  NAND2_X1 U862 ( .A1(G111), .A2(n734), .ZN(n789) );
  NAND2_X1 U863 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U864 ( .A1(G99), .A2(n912), .ZN(n791) );
  XNOR2_X1 U865 ( .A(KEYINPUT77), .B(n791), .ZN(n792) );
  NOR2_X1 U866 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U867 ( .A1(n795), .A2(n794), .ZN(n1023) );
  XNOR2_X1 U868 ( .A(G2096), .B(n1023), .ZN(n796) );
  OR2_X1 U869 ( .A1(G2100), .A2(n796), .ZN(G156) );
  INV_X1 U870 ( .A(G57), .ZN(G237) );
  INV_X1 U871 ( .A(G132), .ZN(G219) );
  INV_X1 U872 ( .A(G82), .ZN(G220) );
  NAND2_X1 U873 ( .A1(G7), .A2(G661), .ZN(n798) );
  XNOR2_X1 U874 ( .A(n798), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U875 ( .A(G223), .ZN(n854) );
  NAND2_X1 U876 ( .A1(n854), .A2(G567), .ZN(n799) );
  XOR2_X1 U877 ( .A(KEYINPUT11), .B(n799), .Z(G234) );
  NAND2_X1 U878 ( .A1(G860), .A2(n953), .ZN(n800) );
  XOR2_X1 U879 ( .A(KEYINPUT69), .B(n800), .Z(G153) );
  NAND2_X1 U880 ( .A1(G868), .A2(G301), .ZN(n802) );
  INV_X1 U881 ( .A(n944), .ZN(n923) );
  INV_X1 U882 ( .A(G868), .ZN(n810) );
  NAND2_X1 U883 ( .A1(n923), .A2(n810), .ZN(n801) );
  NAND2_X1 U884 ( .A1(n802), .A2(n801), .ZN(G284) );
  INV_X1 U885 ( .A(n956), .ZN(G299) );
  NAND2_X1 U886 ( .A1(G868), .A2(G286), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G299), .A2(n810), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(G297) );
  INV_X1 U889 ( .A(G860), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n805), .A2(G559), .ZN(n806) );
  NAND2_X1 U891 ( .A1(n806), .A2(n944), .ZN(n807) );
  XNOR2_X1 U892 ( .A(n807), .B(KEYINPUT16), .ZN(n808) );
  XOR2_X1 U893 ( .A(KEYINPUT75), .B(n808), .Z(G148) );
  NOR2_X1 U894 ( .A1(G559), .A2(n810), .ZN(n809) );
  NAND2_X1 U895 ( .A1(n944), .A2(n809), .ZN(n812) );
  NAND2_X1 U896 ( .A1(n953), .A2(n810), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U898 ( .A(KEYINPUT76), .B(n813), .Z(G282) );
  XNOR2_X1 U899 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n817) );
  XOR2_X1 U900 ( .A(n953), .B(KEYINPUT78), .Z(n815) );
  NAND2_X1 U901 ( .A1(G559), .A2(n944), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n815), .B(n814), .ZN(n834) );
  NOR2_X1 U903 ( .A1(n834), .A2(G860), .ZN(n816) );
  XNOR2_X1 U904 ( .A(n817), .B(n816), .ZN(n828) );
  NAND2_X1 U905 ( .A1(G67), .A2(n818), .ZN(n821) );
  NAND2_X1 U906 ( .A1(G55), .A2(n819), .ZN(n820) );
  NAND2_X1 U907 ( .A1(n821), .A2(n820), .ZN(n827) );
  NAND2_X1 U908 ( .A1(G93), .A2(n822), .ZN(n825) );
  NAND2_X1 U909 ( .A1(G80), .A2(n823), .ZN(n824) );
  NAND2_X1 U910 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U911 ( .A1(n827), .A2(n826), .ZN(n836) );
  XOR2_X1 U912 ( .A(n828), .B(n836), .Z(G145) );
  XNOR2_X1 U913 ( .A(G290), .B(KEYINPUT19), .ZN(n830) );
  XNOR2_X1 U914 ( .A(G288), .B(G166), .ZN(n829) );
  XNOR2_X1 U915 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U916 ( .A(n836), .B(n831), .ZN(n833) );
  XNOR2_X1 U917 ( .A(G305), .B(n956), .ZN(n832) );
  XNOR2_X1 U918 ( .A(n833), .B(n832), .ZN(n924) );
  XNOR2_X1 U919 ( .A(n834), .B(n924), .ZN(n835) );
  NAND2_X1 U920 ( .A1(n835), .A2(G868), .ZN(n838) );
  OR2_X1 U921 ( .A1(G868), .A2(n836), .ZN(n837) );
  NAND2_X1 U922 ( .A1(n838), .A2(n837), .ZN(G295) );
  NAND2_X1 U923 ( .A1(G2084), .A2(G2078), .ZN(n839) );
  XOR2_X1 U924 ( .A(KEYINPUT20), .B(n839), .Z(n840) );
  NAND2_X1 U925 ( .A1(G2090), .A2(n840), .ZN(n841) );
  XNOR2_X1 U926 ( .A(KEYINPUT21), .B(n841), .ZN(n842) );
  NAND2_X1 U927 ( .A1(n842), .A2(G2072), .ZN(n843) );
  XNOR2_X1 U928 ( .A(KEYINPUT86), .B(n843), .ZN(G158) );
  XNOR2_X1 U929 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U930 ( .A1(G220), .A2(G219), .ZN(n844) );
  XOR2_X1 U931 ( .A(KEYINPUT22), .B(n844), .Z(n845) );
  NOR2_X1 U932 ( .A1(G218), .A2(n845), .ZN(n846) );
  NAND2_X1 U933 ( .A1(G96), .A2(n846), .ZN(n859) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n859), .ZN(n850) );
  NAND2_X1 U935 ( .A1(G69), .A2(G120), .ZN(n847) );
  NOR2_X1 U936 ( .A1(G237), .A2(n847), .ZN(n848) );
  NAND2_X1 U937 ( .A1(G108), .A2(n848), .ZN(n860) );
  NAND2_X1 U938 ( .A1(G567), .A2(n860), .ZN(n849) );
  NAND2_X1 U939 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U940 ( .A(KEYINPUT87), .B(n851), .ZN(G319) );
  INV_X1 U941 ( .A(G319), .ZN(n853) );
  NAND2_X1 U942 ( .A1(G661), .A2(G483), .ZN(n852) );
  NOR2_X1 U943 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U944 ( .A1(n858), .A2(G36), .ZN(G176) );
  NAND2_X1 U945 ( .A1(n854), .A2(G2106), .ZN(n855) );
  XOR2_X1 U946 ( .A(KEYINPUT111), .B(n855), .Z(G217) );
  AND2_X1 U947 ( .A1(G15), .A2(G2), .ZN(n856) );
  NAND2_X1 U948 ( .A1(G661), .A2(n856), .ZN(G259) );
  NAND2_X1 U949 ( .A1(G3), .A2(G1), .ZN(n857) );
  NAND2_X1 U950 ( .A1(n858), .A2(n857), .ZN(G188) );
  XOR2_X1 U951 ( .A(G96), .B(KEYINPUT112), .Z(G221) );
  INV_X1 U953 ( .A(G120), .ZN(G236) );
  INV_X1 U954 ( .A(G69), .ZN(G235) );
  NOR2_X1 U955 ( .A1(n860), .A2(n859), .ZN(G325) );
  INV_X1 U956 ( .A(G325), .ZN(G261) );
  XOR2_X1 U957 ( .A(G2100), .B(G2096), .Z(n862) );
  XNOR2_X1 U958 ( .A(KEYINPUT42), .B(G2678), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U960 ( .A(KEYINPUT43), .B(G2090), .Z(n864) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2072), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U963 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U964 ( .A(G2084), .B(G2078), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(G227) );
  XOR2_X1 U966 ( .A(G1986), .B(G1956), .Z(n870) );
  XNOR2_X1 U967 ( .A(G1976), .B(G1971), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U969 ( .A(G1991), .B(G1996), .Z(n872) );
  XNOR2_X1 U970 ( .A(G1966), .B(G1961), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U973 ( .A(KEYINPUT113), .B(G2474), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n878) );
  XOR2_X1 U975 ( .A(G1981), .B(KEYINPUT41), .Z(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(G229) );
  XOR2_X1 U977 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n880) );
  NAND2_X1 U978 ( .A1(G124), .A2(n909), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n880), .B(n879), .ZN(n887) );
  NAND2_X1 U980 ( .A1(G100), .A2(n912), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G112), .A2(n734), .ZN(n881) );
  NAND2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n883), .B(KEYINPUT115), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G136), .A2(n913), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  NOR2_X1 U986 ( .A1(n887), .A2(n886), .ZN(G162) );
  XOR2_X1 U987 ( .A(n888), .B(G162), .Z(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n898) );
  XNOR2_X1 U989 ( .A(KEYINPUT119), .B(KEYINPUT48), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n1023), .B(KEYINPUT116), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U992 ( .A(KEYINPUT46), .B(n893), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n894), .B(KEYINPUT118), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(n898), .B(n897), .Z(n908) );
  NAND2_X1 U996 ( .A1(G103), .A2(n912), .ZN(n900) );
  NAND2_X1 U997 ( .A1(G139), .A2(n913), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n906) );
  NAND2_X1 U999 ( .A1(G127), .A2(n909), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n734), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(KEYINPUT117), .B(n903), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(KEYINPUT47), .B(n904), .ZN(n905) );
  NOR2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n1015) );
  XNOR2_X1 U1005 ( .A(G164), .B(n1015), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n921) );
  NAND2_X1 U1007 ( .A1(G130), .A2(n909), .ZN(n911) );
  NAND2_X1 U1008 ( .A1(G118), .A2(n734), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n918) );
  NAND2_X1 U1010 ( .A1(G106), .A2(n912), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(G142), .A2(n913), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1013 ( .A(KEYINPUT45), .B(n916), .Z(n917) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(G160), .B(n919), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n922), .ZN(G395) );
  XNOR2_X1 U1018 ( .A(n924), .B(n923), .ZN(n925) );
  XNOR2_X1 U1019 ( .A(n925), .B(G286), .ZN(n927) );
  XOR2_X1 U1020 ( .A(n953), .B(G171), .Z(n926) );
  XNOR2_X1 U1021 ( .A(n927), .B(n926), .ZN(n928) );
  NOR2_X1 U1022 ( .A1(G37), .A2(n928), .ZN(G397) );
  XOR2_X1 U1023 ( .A(G2451), .B(G2430), .Z(n930) );
  XNOR2_X1 U1024 ( .A(G2438), .B(G2443), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(n930), .B(n929), .ZN(n936) );
  XOR2_X1 U1026 ( .A(G2435), .B(G2454), .Z(n932) );
  XNOR2_X1 U1027 ( .A(G1348), .B(G1341), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n932), .B(n931), .ZN(n934) );
  XOR2_X1 U1029 ( .A(G2446), .B(G2427), .Z(n933) );
  XNOR2_X1 U1030 ( .A(n934), .B(n933), .ZN(n935) );
  XOR2_X1 U1031 ( .A(n936), .B(n935), .Z(n937) );
  NAND2_X1 U1032 ( .A1(G14), .A2(n937), .ZN(n943) );
  NAND2_X1 U1033 ( .A1(G319), .A2(n943), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(G227), .A2(G229), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(KEYINPUT49), .B(n938), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(G395), .A2(G397), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(G225) );
  INV_X1 U1039 ( .A(G225), .ZN(G308) );
  INV_X1 U1040 ( .A(G108), .ZN(G238) );
  INV_X1 U1041 ( .A(n943), .ZN(G401) );
  XNOR2_X1 U1042 ( .A(KEYINPUT56), .B(G16), .ZN(n969) );
  XNOR2_X1 U1043 ( .A(n944), .B(G1348), .ZN(n946) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n952) );
  XOR2_X1 U1045 ( .A(G1966), .B(G168), .Z(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(KEYINPUT57), .B(n949), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(KEYINPUT122), .B(n950), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n967) );
  XNOR2_X1 U1050 ( .A(G1341), .B(n953), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(G1971), .A2(G303), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n965) );
  XNOR2_X1 U1053 ( .A(G1956), .B(n956), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1055 ( .A(G1961), .B(G301), .Z(n959) );
  XNOR2_X1 U1056 ( .A(KEYINPUT123), .B(n959), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n1045) );
  XOR2_X1 U1062 ( .A(G16), .B(KEYINPUT124), .Z(n995) );
  XNOR2_X1 U1063 ( .A(n970), .B(G5), .ZN(n989) );
  XNOR2_X1 U1064 ( .A(KEYINPUT59), .B(G4), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(n971), .B(KEYINPUT125), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G1348), .B(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(G1341), .B(G19), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G1981), .B(G6), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(G20), .B(G1956), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(n979), .B(KEYINPUT60), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G22), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(G24), .B(G1986), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(G1976), .B(KEYINPUT127), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(n982), .B(G23), .ZN(n983) );
  NAND2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(n985), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT126), .B(G1966), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(G21), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n993), .B(KEYINPUT61), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(G11), .A2(n996), .ZN(n1043) );
  XOR2_X1 U1089 ( .A(G1991), .B(G25), .Z(n997) );
  NAND2_X1 U1090 ( .A1(n997), .A2(G28), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G1996), .B(G32), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(G33), .B(G2072), .ZN(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1004) );
  XOR2_X1 U1094 ( .A(n1000), .B(G27), .Z(n1002) );
  XNOR2_X1 U1095 ( .A(G2067), .B(G26), .ZN(n1001) );
  NOR2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1099 ( .A(KEYINPUT53), .B(n1007), .Z(n1010) );
  XOR2_X1 U1100 ( .A(KEYINPUT54), .B(G34), .Z(n1008) );
  XNOR2_X1 U1101 ( .A(G2084), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(G35), .B(G2090), .ZN(n1011) );
  NOR2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1105 ( .A1(G29), .A2(n1013), .ZN(n1014) );
  XNOR2_X1 U1106 ( .A(n1014), .B(KEYINPUT55), .ZN(n1041) );
  XOR2_X1 U1107 ( .A(G2072), .B(n1015), .Z(n1017) );
  XOR2_X1 U1108 ( .A(G164), .B(G2078), .Z(n1016) );
  NOR2_X1 U1109 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1110 ( .A(KEYINPUT50), .B(n1018), .ZN(n1037) );
  NAND2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(G160), .B(G2084), .ZN(n1024) );
  NAND2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1116 ( .A(n1027), .B(KEYINPUT120), .ZN(n1028) );
  NAND2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1035) );
  XNOR2_X1 U1118 ( .A(G2090), .B(G162), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(n1030), .B(KEYINPUT121), .ZN(n1032) );
  NOR2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1121 ( .A(KEYINPUT51), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1124 ( .A(KEYINPUT52), .B(n1038), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(G29), .A2(n1039), .ZN(n1040) );
  NAND2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NOR2_X1 U1127 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NAND2_X1 U1128 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  XOR2_X1 U1129 ( .A(KEYINPUT62), .B(n1046), .Z(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

