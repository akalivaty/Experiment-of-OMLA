//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n468), .B1(new_n465), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n465), .A2(new_n467), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n463), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n473), .A2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n463), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n475), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT4), .A4(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n463), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n465), .A2(new_n467), .A3(G126), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n463), .A2(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n466), .A2(G2104), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT67), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n492), .B(new_n496), .C1(new_n502), .C2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n513), .A2(G50), .A3(G543), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT68), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n514), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT6), .B(G651), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT70), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n513), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(G543), .A3(new_n527), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n520), .B(new_n522), .C1(new_n523), .C2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n509), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n506), .A2(new_n508), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT69), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n529), .A2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n511), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n525), .A2(G543), .A3(new_n527), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G52), .B1(G90), .B2(new_n519), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(KEYINPUT71), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(KEYINPUT71), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(G651), .A3(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT72), .B(G81), .Z(new_n548));
  AOI22_X1  g123(.A1(new_n540), .A2(G43), .B1(new_n519), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n540), .A2(new_n558), .A3(KEYINPUT9), .A4(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n532), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n519), .A2(G91), .B1(G651), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n528), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n559), .A2(new_n563), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  OR2_X1    g143(.A1(new_n515), .A2(new_n517), .ZN(G303));
  NAND3_X1  g144(.A1(new_n540), .A2(KEYINPUT74), .A3(G49), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n531), .A2(new_n571), .A3(new_n533), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n519), .B2(G87), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  INV_X1    g149(.A(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n528), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n570), .A2(new_n573), .A3(new_n576), .ZN(G288));
  INV_X1    g152(.A(G73), .ZN(new_n578));
  OR3_X1    g153(.A1(new_n578), .A2(new_n505), .A3(KEYINPUT75), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT75), .B1(new_n578), .B2(new_n505), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n532), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(G48), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n532), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(new_n513), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  AND2_X1   g163(.A1(new_n534), .A2(G60), .ZN(new_n589));
  AND2_X1   g164(.A1(G72), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n540), .A2(G47), .B1(G85), .B2(new_n519), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G290));
  AND3_X1   g168(.A1(new_n509), .A2(G92), .A3(new_n513), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n540), .A2(G54), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n511), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G284));
  OAI21_X1  g177(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G321));
  NOR2_X1   g178(.A1(G168), .A2(new_n600), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n559), .A2(new_n563), .A3(new_n566), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(G868), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(KEYINPUT76), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(KEYINPUT76), .B2(new_n604), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(KEYINPUT76), .B2(new_n604), .ZN(G280));
  INV_X1    g185(.A(new_n599), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n550), .A2(new_n600), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n599), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n600), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n500), .A2(new_n501), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n464), .A2(G2105), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n481), .A2(G123), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n483), .A2(G135), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n623), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2435), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2438), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  AND2_X1   g217(.A1(new_n642), .A2(G14), .ZN(G401));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT78), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT17), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT77), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NOR3_X1   g225(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT79), .ZN(new_n652));
  INV_X1    g227(.A(new_n649), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n647), .B2(new_n650), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n644), .B2(new_n650), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n644), .A3(new_n650), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2096), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(G2100), .Z(G227));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT80), .B(KEYINPUT20), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n670), .A2(new_n662), .A3(new_n665), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n668), .B(new_n671), .C1(new_n662), .C2(new_n670), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(G1986), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT22), .B(G1981), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G229));
  XOR2_X1   g254(.A(KEYINPUT31), .B(G11), .Z(new_n680));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(G28), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(G28), .ZN(new_n683));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  AND3_X1   g259(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(G5), .A2(G16), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G171), .B2(G16), .ZN(new_n687));
  AOI211_X1 g262(.A(new_n680), .B(new_n685), .C1(new_n687), .C2(G1961), .ZN(new_n688));
  NOR2_X1   g263(.A1(G16), .A2(G21), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G168), .B2(G16), .ZN(new_n690));
  INV_X1    g265(.A(G1966), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n688), .B(new_n692), .C1(new_n684), .C2(new_n628), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT91), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G29), .A2(G35), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G162), .B2(G29), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT29), .ZN(new_n698));
  INV_X1    g273(.A(G2090), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n693), .A2(new_n694), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G4), .B2(G16), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n702), .A2(G4), .A3(G16), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n703), .B(new_n704), .C1(new_n599), .C2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT86), .B(G1348), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n695), .A2(new_n700), .A3(new_n701), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n684), .A2(G26), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n481), .A2(G128), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n483), .A2(G140), .ZN(new_n712));
  OR2_X1    g287(.A1(G104), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n710), .B1(new_n716), .B2(new_n684), .ZN(new_n717));
  MUX2_X1   g292(.A(new_n710), .B(new_n717), .S(KEYINPUT28), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G2067), .ZN(new_n719));
  NOR2_X1   g294(.A1(G29), .A2(G32), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n481), .A2(G129), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n619), .A2(G105), .ZN(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT26), .ZN(new_n726));
  AOI211_X1 g301(.A(new_n724), .B(new_n726), .C1(G141), .C2(new_n483), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n720), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT27), .B(G1996), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n551), .A2(G16), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G16), .B2(G19), .ZN(new_n734));
  INV_X1    g309(.A(G1341), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT24), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G34), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G160), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n687), .B2(G1961), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n734), .B2(new_n735), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n483), .A2(G139), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n619), .A2(G103), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n618), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n747), .B(new_n750), .C1(new_n751), .C2(new_n463), .ZN(new_n752));
  MUX2_X1   g327(.A(G33), .B(new_n752), .S(G29), .Z(new_n753));
  XOR2_X1   g328(.A(KEYINPUT88), .B(G2072), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n705), .A2(KEYINPUT23), .A3(G20), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT23), .ZN(new_n757));
  INV_X1    g332(.A(G20), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G16), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n759), .C1(new_n606), .C2(new_n705), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G1956), .Z(new_n761));
  NAND4_X1  g336(.A1(new_n736), .A2(new_n746), .A3(new_n755), .A4(new_n761), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n709), .A2(new_n719), .A3(new_n732), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n742), .A2(new_n743), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT89), .Z(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G23), .ZN(new_n766));
  AND3_X1   g341(.A1(new_n570), .A2(new_n573), .A3(new_n576), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT33), .B(G1976), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n705), .A2(G22), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G166), .B2(new_n705), .ZN(new_n772));
  INV_X1    g347(.A(G1971), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n705), .A2(G6), .ZN(new_n775));
  INV_X1    g350(.A(G305), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n705), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT32), .B(G1981), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n770), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT83), .B(KEYINPUT34), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT84), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n780), .B2(new_n781), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n684), .A2(G25), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n483), .A2(G131), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT81), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT82), .ZN(new_n788));
  OR3_X1    g363(.A1(new_n788), .A2(G95), .A3(G2105), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n463), .A2(G107), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n788), .B1(G95), .B2(G2105), .ZN(new_n791));
  AND4_X1   g366(.A1(G2104), .A2(new_n789), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G119), .B2(new_n481), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n786), .A2(KEYINPUT81), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n787), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n785), .B1(new_n796), .B2(new_n684), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT35), .B(G1991), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n797), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G16), .A2(G24), .ZN(new_n801));
  INV_X1    g376(.A(G290), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1986), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n782), .A2(new_n784), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n763), .A2(new_n765), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n684), .A2(G27), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G164), .B2(new_n684), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G2078), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n810), .A2(new_n813), .ZN(G311));
  INV_X1    g389(.A(G311), .ZN(G150));
  NAND2_X1  g390(.A1(new_n534), .A2(G67), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n511), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G55), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n528), .A2(new_n819), .B1(new_n820), .B2(new_n514), .ZN(new_n821));
  OAI21_X1  g396(.A(G860), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n611), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT39), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n818), .A2(new_n821), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(new_n550), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n550), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n826), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n823), .B1(new_n833), .B2(G860), .ZN(G145));
  INV_X1    g409(.A(KEYINPUT93), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n752), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n481), .A2(G130), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n483), .A2(G142), .ZN(new_n838));
  NOR2_X1   g413(.A1(G106), .A2(G2105), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n836), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n795), .B(new_n621), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n728), .A2(G164), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n728), .A2(G164), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n848), .A2(new_n716), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n716), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n752), .A2(new_n835), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n844), .A3(new_n845), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n628), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n854), .A2(new_n855), .A3(new_n857), .A4(new_n628), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G160), .B(G162), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n860), .A2(new_n863), .A3(new_n861), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT95), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n865), .A2(new_n870), .A3(new_n866), .A4(new_n867), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n869), .A2(KEYINPUT40), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT40), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(G395));
  AOI21_X1  g449(.A(new_n599), .B1(new_n606), .B2(KEYINPUT96), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(KEYINPUT96), .B2(new_n606), .ZN(new_n876));
  OR3_X1    g451(.A1(new_n611), .A2(new_n606), .A3(KEYINPUT96), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT41), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n830), .A2(new_n831), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n615), .ZN(new_n882));
  MUX2_X1   g457(.A(new_n878), .B(new_n880), .S(new_n882), .Z(new_n883));
  XNOR2_X1  g458(.A(G290), .B(G305), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G303), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n767), .B(KEYINPUT97), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(KEYINPUT98), .B(KEYINPUT42), .Z(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n883), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(G868), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(G868), .B2(new_n827), .ZN(G295));
  OAI21_X1  g467(.A(new_n891), .B1(G868), .B2(new_n827), .ZN(G331));
  XNOR2_X1  g468(.A(G286), .B(G301), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n832), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n881), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n879), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n881), .B(new_n894), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n898), .B(new_n887), .C1(new_n899), .C2(new_n878), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n866), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n895), .A2(new_n897), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n877), .A3(new_n876), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n887), .B1(new_n904), .B2(new_n898), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT43), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n878), .A2(KEYINPUT99), .A3(KEYINPUT41), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n899), .B(new_n908), .C1(KEYINPUT99), .C2(new_n879), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n887), .B1(new_n909), .B2(new_n904), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n901), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT44), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n901), .B2(new_n905), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n910), .A2(new_n901), .A3(KEYINPUT43), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n913), .B1(new_n917), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g493(.A(G1384), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n492), .A2(new_n496), .ZN(new_n920));
  INV_X1    g495(.A(new_n497), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT4), .B1(new_n618), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g500(.A(KEYINPUT100), .B(G40), .Z(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n472), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n618), .B2(G125), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n478), .B(new_n927), .C1(new_n929), .C2(new_n463), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT102), .ZN(new_n932));
  INV_X1    g507(.A(G1996), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT101), .Z(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n729), .ZN(new_n936));
  INV_X1    g511(.A(G2067), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n715), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n729), .B2(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  AND4_X1   g515(.A1(new_n799), .A2(new_n936), .A3(new_n796), .A4(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n715), .A2(G2067), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n932), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT127), .ZN(new_n944));
  INV_X1    g519(.A(new_n938), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n932), .B1(new_n728), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n935), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n935), .A2(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  XNOR2_X1  g526(.A(new_n795), .B(new_n798), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n952), .A2(KEYINPUT103), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(KEYINPUT103), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n932), .A3(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n936), .A2(new_n940), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(G290), .A2(G1986), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n931), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT48), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n944), .A2(new_n951), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT63), .ZN(new_n962));
  NAND3_X1  g537(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT108), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  NOR2_X1   g540(.A1(G166), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(KEYINPUT55), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(KEYINPUT109), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n966), .A2(new_n969), .A3(KEYINPUT55), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n964), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT110), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n964), .B(new_n973), .C1(new_n968), .C2(new_n970), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n921), .B1(new_n469), .B2(new_n470), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT4), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n463), .B1(new_n493), .B2(new_n494), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n984));
  OAI211_X1 g559(.A(G160), .B(new_n927), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n923), .A2(KEYINPUT105), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n985), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n976), .B1(new_n992), .B2(new_n699), .ZN(new_n993));
  AOI211_X1 g568(.A(KEYINPUT105), .B(G1384), .C1(new_n979), .C2(new_n982), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n987), .B1(new_n503), .B2(new_n919), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n991), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n930), .B1(KEYINPUT50), .B2(new_n923), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n976), .A3(new_n699), .A4(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n925), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n473), .A2(new_n479), .A3(new_n926), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n773), .B1(new_n999), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(G8), .B1(new_n993), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n962), .B1(new_n975), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n996), .A2(KEYINPUT112), .A3(new_n743), .A4(new_n997), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n994), .A2(new_n995), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1002), .B1(new_n1009), .B2(new_n924), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1008), .B1(new_n1010), .B2(G1966), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT112), .B1(new_n992), .B2(new_n743), .ZN(new_n1012));
  OAI21_X1  g587(.A(G8), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(G286), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n968), .A2(new_n970), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n963), .B(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1005), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1000), .B1(new_n994), .B2(new_n995), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n767), .A2(G1976), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(G8), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT52), .ZN(new_n1024));
  OR2_X1    g599(.A1(G305), .A2(G1981), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1025), .A2(KEYINPUT49), .A3(new_n1026), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1029), .A2(new_n1021), .A3(G8), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1021), .A2(new_n1022), .A3(new_n1033), .A4(G8), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1024), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1015), .B1(new_n1020), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT113), .B(new_n1035), .C1(new_n1005), .C2(new_n1019), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1007), .B(new_n1014), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT114), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n996), .A2(new_n997), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT107), .B1(new_n1041), .B2(G2090), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n998), .A3(new_n1003), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n971), .B1(new_n1043), .B2(G8), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT113), .B1(new_n1044), .B2(new_n1035), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1020), .A2(new_n1015), .A3(new_n1036), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n1014), .A4(new_n1007), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n975), .A2(new_n1006), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n999), .A2(new_n1002), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(G1971), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1000), .B1(KEYINPUT50), .B2(new_n923), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n1009), .B2(new_n990), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n699), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1019), .B1(new_n1055), .B2(new_n965), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT111), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1035), .B(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1050), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1014), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n962), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1040), .A2(new_n1049), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n930), .B1(new_n986), .B2(new_n988), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1031), .A2(new_n1032), .A3(new_n767), .ZN(new_n1064));
  AOI211_X1 g639(.A(new_n965), .B(new_n1063), .C1(new_n1064), .C2(new_n1025), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1050), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n1036), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G286), .A2(G8), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT51), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1013), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n996), .A2(new_n743), .A3(new_n997), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n930), .B1(KEYINPUT45), .B2(new_n983), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n989), .B2(KEYINPUT45), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n691), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1080), .A3(new_n1008), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1081), .A2(G8), .A3(G286), .ZN(new_n1082));
  OAI211_X1 g657(.A(G8), .B(new_n1072), .C1(new_n1081), .C2(G286), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1074), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1074), .A2(KEYINPUT121), .A3(new_n1083), .A4(new_n1082), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT62), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1090), .A3(new_n1087), .ZN(new_n1091));
  INV_X1    g666(.A(G2078), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1051), .A2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1094));
  INV_X1    g669(.A(G1961), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1093), .A2(new_n1094), .B1(new_n1041), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1010), .A2(new_n1097), .A3(new_n1092), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT53), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1097), .B1(new_n1010), .B2(new_n1092), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G171), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1089), .A2(new_n1091), .A3(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n925), .A2(new_n1000), .A3(new_n1001), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1078), .A2(KEYINPUT115), .A3(new_n925), .A4(new_n1105), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n930), .B1(new_n984), .B2(new_n983), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1956), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G299), .B(KEYINPUT57), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(KEYINPUT117), .ZN(new_n1116));
  NOR4_X1   g691(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1116), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1108), .B(new_n1109), .C1(new_n1054), .C2(G1956), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1119), .B2(new_n1114), .ZN(new_n1120));
  OR3_X1    g695(.A1(new_n1110), .A2(new_n1114), .A3(new_n1113), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1117), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1114), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1119), .A2(KEYINPUT116), .A3(new_n1114), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1115), .A3(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT58), .B(G1341), .Z(new_n1128));
  AOI22_X1  g703(.A1(new_n1051), .A2(new_n933), .B1(new_n1021), .B2(new_n1128), .ZN(new_n1129));
  OR3_X1    g704(.A1(new_n1129), .A2(KEYINPUT59), .A3(new_n550), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT59), .B1(new_n1129), .B2(new_n550), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n599), .A2(KEYINPUT118), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n992), .A2(new_n707), .B1(G2067), .B2(new_n1021), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n707), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1041), .A2(new_n1138), .B1(new_n937), .B2(new_n1063), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n599), .A2(KEYINPUT118), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1139), .A2(KEYINPUT60), .A3(new_n1133), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1122), .A2(new_n1127), .A3(new_n1132), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1123), .B1(new_n599), .B2(new_n1139), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1121), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT119), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1092), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n925), .A2(G160), .A3(new_n1001), .A4(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT125), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1096), .A2(G301), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1149), .B1(new_n1102), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1096), .A2(new_n1152), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(G171), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1157), .B(KEYINPUT54), .C1(new_n1101), .C2(G171), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1144), .A2(new_n1159), .A3(new_n1146), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1148), .A2(new_n1155), .A3(new_n1158), .A4(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1104), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1059), .B(KEYINPUT126), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1068), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n802), .A2(new_n804), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n931), .B1(new_n1165), .B2(new_n957), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n956), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT104), .Z(new_n1168));
  OAI21_X1  g743(.A(new_n961), .B1(new_n1164), .B2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g744(.A(G319), .B1(new_n915), .B2(new_n916), .ZN(new_n1171));
  NOR2_X1   g745(.A1(G227), .A2(G401), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n1172), .A2(new_n868), .ZN(new_n1173));
  NOR3_X1   g747(.A1(new_n1171), .A2(G229), .A3(new_n1173), .ZN(G308));
  OR3_X1    g748(.A1(new_n910), .A2(new_n901), .A3(KEYINPUT43), .ZN(new_n1175));
  AOI21_X1  g749(.A(new_n461), .B1(new_n1175), .B2(new_n914), .ZN(new_n1176));
  NAND4_X1  g750(.A1(new_n1176), .A2(new_n678), .A3(new_n868), .A4(new_n1172), .ZN(G225));
endmodule


