//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n209), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  INV_X1    g0020(.A(new_n201), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(new_n218), .A2(KEYINPUT0), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n224), .B1(KEYINPUT0), .B2(new_n218), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT64), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT66), .ZN(new_n229));
  AND2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n227), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n232), .A2(KEYINPUT67), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(KEYINPUT67), .ZN(new_n235));
  AOI22_X1  g0035(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  AOI22_X1  g0037(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n238));
  NAND3_X1  g0038(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g0039(.A(new_n213), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g0040(.A(new_n226), .B1(KEYINPUT1), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g0041(.A(new_n241), .B1(KEYINPUT1), .B2(new_n240), .ZN(G361));
  XOR2_X1   g0042(.A(G238), .B(G244), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G264), .B(G270), .Z(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n202), .A2(G68), .ZN(new_n254));
  INV_X1    g0054(.A(G68), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(G58), .B(G77), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n253), .B(new_n259), .ZN(G351));
  NAND3_X1  g0060(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n255), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT12), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n265), .A2(G50), .B1(G20), .B2(new_n255), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G77), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n219), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(KEYINPUT11), .A3(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n262), .A2(new_n273), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n211), .A2(G1), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G68), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n264), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT11), .B1(new_n271), .B2(new_n273), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n284), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(G238), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n289), .A2(new_n291), .A3(G226), .A4(new_n292), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n289), .A2(new_n291), .A3(G232), .A4(G1698), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n293), .B(new_n294), .C1(new_n267), .C2(new_n205), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n282), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT13), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n288), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n298), .A2(G190), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n288), .A2(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n281), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(KEYINPUT72), .A3(new_n298), .ZN(new_n303));
  OR3_X1    g0103(.A1(new_n300), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(G200), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n289), .A2(new_n291), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(G232), .A3(new_n292), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(G238), .A3(G1698), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n310), .B(new_n311), .C1(new_n206), .C2(new_n309), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n282), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n285), .B1(G244), .B2(new_n287), .ZN(new_n314));
  AOI21_X1  g0114(.A(G169), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n314), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n315), .A2(new_n316), .B1(new_n317), .B2(G179), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n313), .A2(KEYINPUT70), .A3(new_n319), .A4(new_n314), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n269), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n273), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n276), .A2(new_n270), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n275), .A2(new_n327), .B1(new_n270), .B2(new_n262), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n317), .B2(G200), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n313), .A2(G190), .A3(new_n314), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n318), .A2(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n309), .A2(G222), .A3(new_n292), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n309), .A2(G223), .A3(G1698), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n334), .B(new_n335), .C1(new_n270), .C2(new_n309), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n282), .ZN(new_n337));
  XOR2_X1   g0137(.A(KEYINPUT68), .B(G226), .Z(new_n338));
  AOI21_X1  g0138(.A(new_n285), .B1(new_n287), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(G190), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT9), .ZN(new_n341));
  INV_X1    g0141(.A(new_n273), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n322), .A2(new_n268), .B1(G150), .B2(new_n265), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n203), .A2(G20), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n277), .A2(KEYINPUT69), .A3(G50), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT69), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n276), .B2(new_n202), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n275), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n262), .A2(new_n202), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n341), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n343), .A2(new_n344), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n273), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n354), .A2(KEYINPUT9), .A3(new_n350), .A4(new_n349), .ZN(new_n355));
  AND3_X1   g0155(.A1(new_n340), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n337), .A2(new_n339), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G200), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n356), .B(new_n358), .C1(KEYINPUT71), .C2(KEYINPUT10), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n345), .A2(new_n351), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(G179), .B2(new_n357), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT10), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n340), .A2(new_n355), .A3(KEYINPUT71), .A4(new_n352), .ZN(new_n366));
  INV_X1    g0166(.A(new_n358), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n340), .A2(new_n355), .A3(new_n352), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n365), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n333), .A2(new_n359), .A3(new_n364), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n303), .A2(new_n304), .A3(G169), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n298), .A2(G179), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n371), .A2(KEYINPUT14), .B1(new_n301), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n303), .A2(new_n304), .A3(new_n374), .A4(G169), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n375), .A2(new_n376), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI211_X1 g0179(.A(new_n307), .B(new_n370), .C1(new_n379), .C2(new_n281), .ZN(new_n380));
  AND2_X1   g0180(.A1(G58), .A2(G68), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(new_n201), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G20), .B1(G159), .B2(new_n265), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT76), .ZN(new_n384));
  NAND2_X1  g0184(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n290), .A2(KEYINPUT74), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n388), .A3(G33), .ZN(new_n389));
  AOI21_X1  g0189(.A(G20), .B1(new_n389), .B2(new_n289), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n385), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n289), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(G33), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n396), .A2(G20), .A3(new_n391), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n384), .B(G68), .C1(new_n393), .C2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n391), .B1(new_n396), .B2(G20), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n389), .A2(new_n289), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(new_n211), .A3(new_n392), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n402), .A3(new_n385), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n384), .B1(new_n403), .B2(G68), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT16), .B(new_n383), .C1(new_n399), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n309), .B2(G20), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n407), .A2(G20), .ZN(new_n409));
  AOI21_X1  g0209(.A(G33), .B1(new_n386), .B2(new_n388), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n255), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n383), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n406), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n405), .A2(new_n415), .A3(new_n273), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n321), .A2(new_n276), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n275), .B1(new_n262), .B2(new_n321), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n285), .B1(G232), .B2(new_n287), .ZN(new_n419));
  INV_X1    g0219(.A(new_n282), .ZN(new_n420));
  MUX2_X1   g0220(.A(G223), .B(G226), .S(G1698), .Z(new_n421));
  AOI22_X1  g0221(.A1(new_n396), .A2(new_n421), .B1(G33), .B2(G87), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G200), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G190), .B2(new_n423), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n416), .A2(new_n418), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(KEYINPUT77), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT77), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n416), .A2(new_n431), .A3(new_n426), .A4(new_n418), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n429), .B1(new_n433), .B2(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n416), .A2(new_n418), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n423), .A2(G169), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n319), .B2(new_n423), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(KEYINPUT18), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n440), .B1(new_n435), .B2(new_n437), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n380), .A2(new_n434), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n262), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT25), .B1(new_n262), .B2(new_n206), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n210), .A2(G33), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n342), .A2(new_n261), .A3(new_n447), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n445), .A2(new_n446), .B1(new_n448), .B2(new_n206), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n396), .A2(KEYINPUT22), .A3(new_n211), .A4(G87), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT22), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n211), .A2(G87), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n308), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G116), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G20), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n211), .B2(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n450), .A2(new_n453), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT24), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT24), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n450), .A2(new_n453), .A3(new_n462), .A4(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n449), .B1(new_n464), .B2(new_n273), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT85), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G250), .A2(G1698), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n216), .B2(G1698), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n396), .A2(new_n468), .B1(G33), .B2(G294), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n466), .B1(new_n469), .B2(new_n420), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  INV_X1    g0273(.A(G41), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT5), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT79), .B1(new_n476), .B2(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(G41), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n472), .B(new_n475), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n479), .A2(G264), .A3(new_n420), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n479), .A2(new_n283), .A3(new_n282), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n470), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n468), .A2(new_n389), .A3(new_n289), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G294), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n420), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT85), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n362), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT86), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n479), .A2(G264), .A3(new_n420), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n490), .B(new_n491), .C1(new_n469), .C2(new_n420), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT86), .B1(new_n486), .B2(new_n480), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n481), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G179), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n465), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G190), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n470), .A2(new_n487), .A3(new_n482), .A4(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n494), .B2(G200), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n465), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n465), .A3(KEYINPUT87), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n496), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n324), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n261), .ZN(new_n506));
  INV_X1    g0306(.A(G87), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n448), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  XOR2_X1   g0309(.A(KEYINPUT78), .B(G97), .Z(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n269), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n389), .A2(new_n211), .A3(G68), .A4(new_n289), .ZN(new_n512));
  OR2_X1    g0312(.A1(KEYINPUT78), .A2(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(KEYINPUT78), .A2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n515), .A2(G87), .A3(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n267), .A2(new_n205), .ZN(new_n517));
  AOI21_X1  g0317(.A(G20), .B1(new_n517), .B2(KEYINPUT19), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n511), .B(new_n512), .C1(new_n516), .C2(new_n518), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n506), .B(new_n508), .C1(new_n519), .C2(new_n273), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n282), .A2(new_n283), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n472), .A2(new_n209), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n521), .A2(new_n472), .B1(new_n420), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(G238), .A2(G1698), .ZN(new_n524));
  INV_X1    g0324(.A(G244), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G1698), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n396), .A2(new_n526), .B1(G33), .B2(G116), .ZN(new_n527));
  OAI211_X1 g0327(.A(G190), .B(new_n523), .C1(new_n527), .C2(new_n420), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n389), .A3(new_n289), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n420), .B1(new_n531), .B2(new_n454), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n420), .A2(G274), .A3(new_n472), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n420), .A2(new_n522), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(KEYINPUT82), .A3(G190), .ZN(new_n537));
  OAI21_X1  g0337(.A(G200), .B1(new_n532), .B2(new_n535), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n520), .A2(new_n530), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n519), .A2(new_n273), .ZN(new_n540));
  INV_X1    g0340(.A(new_n506), .ZN(new_n541));
  INV_X1    g0341(.A(new_n448), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n505), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n523), .B1(new_n527), .B2(new_n420), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n362), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n536), .A2(new_n319), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n539), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n206), .B1(new_n408), .B2(new_n412), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n513), .B2(new_n514), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT6), .B1(new_n207), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(G20), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n265), .A2(G77), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n273), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n261), .A2(G97), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n542), .B2(G97), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n479), .A2(G257), .A3(new_n420), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT4), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n525), .A2(G1698), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n401), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(KEYINPUT4), .A2(G244), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n289), .A2(new_n291), .A3(new_n569), .A4(new_n292), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n289), .A2(new_n291), .A3(G250), .A4(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G283), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n564), .B1(new_n574), .B2(new_n282), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n477), .A2(new_n478), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n521), .A2(new_n576), .A3(new_n472), .A4(new_n475), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n562), .B1(G200), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT4), .B1(new_n396), .B2(new_n566), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n282), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n582), .A2(G190), .A3(new_n577), .A4(new_n563), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT80), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT80), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n575), .A2(new_n585), .A3(G190), .A4(new_n577), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n579), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT81), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n559), .A2(new_n589), .A3(new_n561), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n559), .B2(new_n561), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n362), .B1(new_n575), .B2(new_n577), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n420), .B1(new_n568), .B2(new_n573), .ZN(new_n594));
  NOR4_X1   g0394(.A1(new_n594), .A2(new_n319), .A3(new_n564), .A4(new_n481), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n591), .A2(new_n592), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n550), .A2(new_n588), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n217), .A2(G1698), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(G257), .B2(G1698), .ZN(new_n599));
  INV_X1    g0399(.A(G303), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n401), .A2(new_n599), .B1(new_n600), .B2(new_n309), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n282), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n479), .A2(G270), .A3(new_n420), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n577), .A2(KEYINPUT83), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT83), .B1(new_n577), .B2(new_n603), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n261), .A2(G116), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n542), .B2(G116), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G20), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n273), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT84), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n273), .A2(KEYINPUT84), .A3(new_n611), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n211), .B(new_n572), .C1(new_n510), .C2(G33), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(KEYINPUT20), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT20), .B1(new_n616), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n609), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n607), .A2(new_n621), .A3(G169), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n577), .A2(new_n603), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT83), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(new_n604), .B1(new_n282), .B2(new_n601), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(new_n621), .A3(G179), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n602), .B(G190), .C1(new_n605), .C2(new_n606), .ZN(new_n630));
  INV_X1    g0430(.A(new_n609), .ZN(new_n631));
  INV_X1    g0431(.A(new_n620), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n618), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n630), .B(new_n633), .C1(new_n628), .C2(new_n424), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n607), .A2(new_n621), .A3(KEYINPUT21), .A4(G169), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n624), .A2(new_n629), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n597), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n444), .A2(new_n504), .A3(new_n637), .ZN(G372));
  AND2_X1   g0438(.A1(new_n359), .A2(new_n369), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n379), .A2(new_n281), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n318), .A2(new_n330), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n307), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n642), .A2(new_n434), .ZN(new_n643));
  INV_X1    g0443(.A(new_n442), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n364), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT88), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n499), .A2(KEYINPUT87), .A3(new_n465), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT87), .B1(new_n499), .B2(new_n465), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n506), .B1(new_n519), .B2(new_n273), .ZN(new_n651));
  INV_X1    g0451(.A(new_n508), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n651), .A2(new_n538), .A3(new_n528), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n548), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n588), .A2(new_n596), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n647), .B1(new_n650), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n502), .A2(new_n503), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n588), .A2(new_n596), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT88), .A4(new_n655), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n464), .A2(new_n273), .ZN(new_n661));
  INV_X1    g0461(.A(new_n449), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n495), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n488), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n635), .A2(new_n629), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n624), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n657), .A2(new_n660), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n548), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n575), .A2(G179), .A3(new_n577), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n594), .A2(new_n481), .A3(new_n564), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n362), .B2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n562), .A3(new_n548), .A4(new_n653), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT89), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n596), .A2(new_n549), .A3(new_n674), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n673), .A2(KEYINPUT89), .A3(new_n674), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n669), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n668), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n444), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n646), .A2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n666), .A2(new_n624), .ZN(new_n683));
  INV_X1    g0483(.A(G13), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n684), .A2(G1), .A3(G20), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT90), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(G213), .B1(new_n687), .B2(KEYINPUT27), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT27), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(KEYINPUT91), .B(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n633), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n683), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n636), .B2(new_n696), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n504), .B1(new_n465), .B2(new_n695), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n665), .B2(new_n695), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n683), .A2(new_n695), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n706), .A2(new_n504), .B1(new_n496), .B2(new_n695), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(G399));
  NOR2_X1   g0508(.A1(new_n215), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n516), .A2(new_n610), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n222), .B2(new_n710), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n680), .A2(new_n716), .A3(new_n695), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n667), .A2(new_n658), .A3(new_n659), .A4(new_n655), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n562), .B1(new_n593), .B2(new_n595), .ZN(new_n719));
  OAI21_X1  g0519(.A(KEYINPUT26), .B1(new_n719), .B2(new_n654), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n548), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n596), .A2(new_n549), .A3(KEYINPUT26), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT93), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n593), .ZN(new_n724));
  INV_X1    g0524(.A(new_n592), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n724), .A2(new_n670), .B1(new_n725), .B2(new_n590), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n550), .A3(new_n674), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT93), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(new_n548), .A4(new_n720), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n718), .A2(new_n723), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n695), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n717), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT31), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n545), .A2(new_n594), .A3(new_n564), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n628), .A2(new_n494), .A3(new_n735), .A4(G179), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n736), .A2(KEYINPUT92), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n737), .B1(new_n736), .B2(KEYINPUT92), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n607), .A2(new_n578), .A3(new_n319), .A4(new_n545), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n494), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n734), .B1(new_n742), .B2(new_n695), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n637), .A2(new_n504), .A3(new_n695), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT30), .ZN(new_n746));
  INV_X1    g0546(.A(new_n741), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(KEYINPUT31), .B(new_n694), .C1(new_n748), .C2(new_n738), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n743), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n733), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n715), .B1(new_n753), .B2(G1), .ZN(G364));
  NOR2_X1   g0554(.A1(new_n684), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n210), .B1(new_n755), .B2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n709), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n699), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n219), .B1(G20), .B2(new_n362), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n215), .A2(new_n396), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n471), .B2(new_n223), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n471), .B2(new_n259), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n214), .A2(new_n309), .ZN(new_n771));
  INV_X1    g0571(.A(G355), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n771), .A2(new_n772), .B1(G116), .B2(new_n214), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT94), .Z(new_n774));
  AOI21_X1  g0574(.A(new_n766), .B1(new_n770), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n497), .A2(new_n424), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(G20), .A3(new_n319), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n600), .ZN(new_n778));
  NOR4_X1   g0578(.A1(new_n211), .A2(new_n424), .A3(G179), .A4(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n211), .A2(new_n319), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(new_n497), .A3(G200), .ZN(new_n783));
  XOR2_X1   g0583(.A(KEYINPUT33), .B(G317), .Z(new_n784));
  OAI22_X1  g0584(.A1(new_n780), .A2(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n782), .A2(new_n776), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n778), .B(new_n785), .C1(G326), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G190), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G294), .ZN(new_n792));
  NOR4_X1   g0592(.A1(new_n211), .A2(new_n319), .A3(G190), .A4(G200), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n309), .B1(new_n793), .B2(G311), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n211), .A2(new_n319), .A3(new_n497), .A4(G200), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n789), .A2(G20), .A3(new_n497), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n795), .A2(G322), .B1(new_n797), .B2(G329), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n788), .A2(new_n792), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n780), .A2(new_n206), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n309), .B1(new_n777), .B2(new_n507), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n800), .B1(KEYINPUT96), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(KEYINPUT96), .B2(new_n801), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT97), .Z(new_n804));
  INV_X1    g0604(.A(new_n783), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n805), .A2(G68), .B1(new_n795), .B2(G58), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n793), .A2(KEYINPUT95), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n806), .B1(new_n202), .B2(new_n786), .C1(new_n810), .C2(new_n270), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n796), .A2(KEYINPUT32), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT32), .B1(new_n796), .B2(new_n812), .ZN(new_n814));
  INV_X1    g0614(.A(new_n791), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n205), .ZN(new_n816));
  OR3_X1    g0616(.A1(new_n811), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n799), .B1(new_n804), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n775), .B1(new_n818), .B2(new_n764), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n759), .B1(new_n763), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n698), .B(G330), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n821), .B2(new_n759), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT98), .ZN(G396));
  AOI21_X1  g0623(.A(new_n694), .B1(new_n668), .B2(new_n679), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n694), .A2(new_n329), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n641), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n333), .B2(new_n825), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n824), .B(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n758), .B1(new_n829), .B2(new_n751), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n751), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n764), .A2(new_n760), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n759), .B1(new_n270), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n764), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G132), .A2(new_n797), .B1(new_n779), .B2(G68), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n202), .B2(new_n777), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n401), .B(new_n836), .C1(G58), .C2(new_n791), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n805), .A2(G150), .B1(new_n787), .B2(G137), .ZN(new_n838));
  INV_X1    g0638(.A(G143), .ZN(new_n839));
  INV_X1    g0639(.A(new_n795), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n838), .B1(new_n839), .B2(new_n840), .C1(new_n810), .C2(new_n812), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n837), .B1(new_n842), .B2(KEYINPUT34), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n810), .A2(new_n610), .B1(new_n781), .B2(new_n783), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT99), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n780), .A2(new_n507), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G303), .B2(new_n787), .ZN(new_n850));
  INV_X1    g0650(.A(G294), .ZN(new_n851));
  INV_X1    g0651(.A(G311), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n850), .B1(new_n851), .B2(new_n840), .C1(new_n852), .C2(new_n796), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n847), .A2(KEYINPUT99), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n308), .B1(new_n777), .B2(new_n206), .C1(new_n815), .C2(new_n205), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n846), .B1(new_n848), .B2(new_n856), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n833), .B1(new_n834), .B2(new_n857), .C1(new_n828), .C2(new_n761), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n831), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  NOR2_X1   g0660(.A1(new_n755), .A2(new_n210), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n640), .A2(new_n306), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n694), .A2(new_n281), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT100), .Z(new_n864));
  XNOR2_X1  g0664(.A(new_n862), .B(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n750), .A3(new_n828), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n430), .A2(new_n432), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n405), .A2(new_n273), .ZN(new_n869));
  OAI21_X1  g0669(.A(G68), .B1(new_n393), .B2(new_n397), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT76), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n398), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n872), .B2(new_n383), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n418), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT101), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(KEYINPUT101), .B(new_n418), .C1(new_n869), .C2(new_n873), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n691), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n437), .A3(new_n877), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n868), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT37), .B1(new_n435), .B2(new_n437), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n691), .B(KEYINPUT102), .Z(new_n883));
  NAND2_X1  g0683(.A1(new_n435), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n882), .A2(new_n430), .A3(new_n432), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n434), .A2(new_n442), .ZN(new_n887));
  INV_X1    g0687(.A(new_n878), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n885), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n880), .B2(KEYINPUT37), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n878), .B1(new_n434), .B2(new_n442), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n890), .A2(new_n895), .A3(KEYINPUT103), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT103), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n892), .B2(new_n893), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n867), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n434), .A2(KEYINPUT105), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT105), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n429), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n442), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n884), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n891), .A2(KEYINPUT104), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT104), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n438), .A2(new_n884), .A3(new_n427), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n885), .A2(new_n911), .B1(new_n912), .B2(KEYINPUT37), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n908), .A2(new_n909), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n898), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n866), .A2(new_n902), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n903), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n444), .A2(new_n750), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT107), .Z(new_n920));
  AOI21_X1  g0720(.A(new_n700), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT103), .B1(new_n890), .B2(new_n895), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n898), .A2(new_n897), .A3(new_n899), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n641), .A2(new_n694), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n824), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n827), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n925), .A2(new_n929), .A3(new_n865), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n907), .A2(new_n442), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n906), .A2(new_n905), .A3(new_n429), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n909), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n910), .A2(new_n913), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n931), .B1(new_n936), .B2(new_n895), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n640), .A2(new_n694), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n898), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n442), .A2(new_n883), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n930), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT106), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n716), .B1(new_n730), .B2(new_n695), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n716), .B2(new_n824), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n945), .B2(new_n443), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n733), .A2(new_n444), .A3(KEYINPUT106), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n646), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n942), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n861), .B1(new_n922), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n922), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n553), .A2(new_n555), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(KEYINPUT35), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(KEYINPUT35), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(G116), .A3(new_n220), .A4(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT36), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n381), .A2(new_n270), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n254), .B1(new_n222), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(G1), .A3(new_n684), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n952), .A2(new_n957), .A3(new_n960), .ZN(G367));
  INV_X1    g0761(.A(new_n562), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n659), .B1(new_n962), .B2(new_n695), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n672), .A2(new_n562), .A3(new_n694), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n707), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT44), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n707), .A2(new_n965), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT45), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n970), .B(new_n971), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n706), .A2(new_n504), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n703), .B2(new_n706), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(new_n701), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n753), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n977), .A2(new_n752), .A3(new_n733), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n709), .B(KEYINPUT41), .Z(new_n979));
  OAI21_X1  g0779(.A(new_n756), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n695), .A2(new_n520), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n669), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n654), .B2(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT108), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n973), .B1(new_n963), .B2(new_n964), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(KEYINPUT42), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n665), .B1(new_n963), .B2(new_n964), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n695), .B1(new_n989), .B2(new_n726), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT42), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n990), .B1(new_n986), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n985), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n704), .B1(new_n963), .B2(new_n964), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n980), .A2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n765), .B1(new_n214), .B2(new_n324), .C1(new_n768), .C2(new_n249), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n999), .A2(new_n758), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G317), .A2(new_n797), .B1(new_n779), .B2(new_n515), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n852), .B2(new_n786), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n840), .A2(new_n600), .B1(new_n851), .B2(new_n783), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1002), .A2(new_n396), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n777), .A2(new_n610), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n1005), .A2(KEYINPUT46), .B1(new_n815), .B2(new_n206), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT46), .B2(new_n1005), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1004), .B(new_n1007), .C1(new_n781), .C2(new_n810), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n309), .B1(new_n783), .B2(new_n812), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n780), .A2(new_n270), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(G137), .C2(new_n797), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n810), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(G50), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n791), .A2(G68), .ZN(new_n1014));
  INV_X1    g0814(.A(G150), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n840), .A2(new_n1015), .B1(new_n786), .B2(new_n839), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n777), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1016), .B1(G58), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1008), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  INV_X1    g0821(.A(new_n762), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1000), .B1(new_n1021), .B2(new_n834), .C1(new_n983), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n998), .A2(new_n1023), .ZN(G387));
  OR2_X1    g0824(.A1(new_n703), .A2(new_n1022), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n712), .A2(new_n771), .B1(G107), .B2(new_n214), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n246), .ZN(new_n1027));
  AOI21_X1  g0827(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1028));
  AOI21_X1  g0828(.A(KEYINPUT50), .B1(new_n322), .B2(new_n202), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n322), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n712), .B(new_n1028), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n767), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1027), .A2(G45), .B1(new_n1032), .B2(KEYINPUT110), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1032), .A2(KEYINPUT110), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1026), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n758), .B1(new_n1035), .B2(new_n766), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n815), .A2(new_n324), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G50), .B2(new_n795), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT111), .Z(new_n1039));
  OAI22_X1  g0839(.A1(new_n780), .A2(new_n205), .B1(new_n812), .B2(new_n786), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n783), .A2(new_n321), .B1(new_n1015), .B2(new_n796), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1017), .A2(G77), .B1(G68), .B2(new_n793), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1039), .A2(new_n396), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G326), .A2(new_n797), .B1(new_n779), .B2(G116), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n815), .A2(new_n781), .B1(new_n777), .B2(new_n851), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n805), .A2(G311), .B1(new_n787), .B2(G322), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT112), .ZN(new_n1048));
  INV_X1    g0848(.A(G317), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1048), .B1(new_n600), .B2(new_n810), .C1(new_n1049), .C2(new_n840), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n401), .B(new_n1045), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1044), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1036), .B1(new_n1057), .B2(new_n764), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n975), .A2(new_n757), .B1(new_n1025), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n976), .A2(new_n709), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n975), .A2(new_n753), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(G393));
  AND2_X1   g0862(.A1(new_n970), .A2(new_n704), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT113), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(KEYINPUT113), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n704), .C2(new_n970), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n976), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n709), .C1(new_n976), .C2(new_n972), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1066), .A2(new_n756), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n765), .B1(new_n214), .B2(new_n510), .C1(new_n768), .C2(new_n253), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n758), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n840), .A2(new_n852), .B1(new_n786), .B2(new_n1049), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n805), .A2(G303), .B1(G294), .B2(new_n793), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n309), .B(new_n800), .C1(G116), .C2(new_n791), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1017), .A2(G283), .B1(G322), .B2(new_n797), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n777), .A2(new_n255), .B1(new_n839), .B2(new_n796), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1078), .B(new_n849), .C1(G50), .C2(new_n805), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n401), .B1(G77), .B2(new_n791), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n1080), .C1(new_n321), .C2(new_n810), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n787), .A2(G150), .B1(new_n795), .B2(G159), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1077), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1071), .B1(new_n1084), .B2(new_n764), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n965), .B2(new_n1022), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1068), .A2(new_n1069), .A3(new_n1086), .ZN(G390));
  NAND2_X1  g0887(.A1(new_n752), .A2(new_n444), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT106), .B1(new_n733), .B2(new_n444), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n943), .B(new_n443), .C1(new_n717), .C2(new_n732), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n646), .B(new_n1088), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT114), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT116), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT115), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n827), .B1(new_n751), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n750), .A2(KEYINPUT115), .A3(G330), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n865), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n730), .A2(new_n695), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n926), .B1(new_n1099), .B2(new_n828), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n865), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n750), .A2(G330), .A3(new_n828), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1094), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n927), .B1(new_n731), .B2(new_n827), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1102), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n865), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n750), .A2(KEYINPUT115), .A3(G330), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT115), .B1(new_n750), .B2(G330), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n827), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1107), .B(KEYINPUT116), .C1(new_n1110), .C2(new_n865), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1106), .A2(new_n865), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n929), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1104), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n948), .A2(KEYINPUT114), .A3(new_n646), .A4(new_n1088), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1093), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1112), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n937), .A2(new_n939), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n929), .A2(new_n865), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n938), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n936), .A2(new_n895), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1121), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1118), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n937), .A2(new_n939), .B1(new_n1121), .B2(new_n1120), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1129), .A2(new_n1112), .A3(new_n1126), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1117), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1093), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1112), .B1(new_n1129), .B2(new_n1126), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1123), .A2(new_n1118), .A3(new_n1127), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1131), .A2(new_n709), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n759), .B1(new_n321), .B2(new_n832), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n787), .A2(G283), .B1(G68), .B2(new_n779), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n206), .B2(new_n783), .C1(new_n851), .C2(new_n796), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n309), .B(new_n1139), .C1(G87), .C2(new_n1017), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n795), .A2(G116), .B1(new_n791), .B2(G77), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT118), .Z(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n510), .C2(new_n810), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n805), .A2(G137), .B1(G125), .B2(new_n797), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n787), .A2(G128), .B1(new_n795), .B2(G132), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n1012), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n308), .B1(new_n779), .B2(G50), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT117), .Z(new_n1151));
  NAND2_X1  g0951(.A1(new_n1017), .A2(G150), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1152), .A2(KEYINPUT53), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1152), .A2(KEYINPUT53), .B1(G159), .B2(new_n791), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1149), .A2(new_n1151), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1143), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1137), .B1(new_n1156), .B2(new_n834), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1119), .B2(new_n760), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n757), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1136), .A2(new_n1160), .ZN(G378));
  INV_X1    g0961(.A(new_n942), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n639), .A2(new_n364), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n692), .A2(new_n361), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1163), .B(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n700), .B1(new_n915), .B2(new_n916), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1167), .B1(new_n903), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n866), .B1(new_n923), .B2(new_n924), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1167), .C1(new_n1170), .C2(KEYINPUT40), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1162), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1167), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1170), .A2(KEYINPUT40), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1168), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n942), .A3(new_n1171), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1173), .A2(KEYINPUT120), .A3(new_n1178), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1093), .A2(new_n1116), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1135), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT120), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1177), .A2(new_n1182), .A3(new_n942), .A4(new_n1171), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1179), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n710), .B1(new_n1187), .B2(new_n1181), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1179), .A2(new_n757), .A3(new_n1183), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n401), .A2(new_n474), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n779), .A2(G58), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n270), .B2(new_n777), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(G283), .C2(new_n797), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT119), .Z(new_n1195));
  AOI22_X1  g0995(.A1(new_n787), .A2(G116), .B1(new_n795), .B2(G107), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n805), .A2(G97), .B1(new_n793), .B2(new_n505), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1195), .A2(new_n1014), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT58), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1017), .A2(new_n1148), .B1(new_n795), .B2(G128), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n805), .A2(G132), .B1(G137), .B2(new_n793), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n787), .A2(G125), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n791), .A2(G150), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n797), .A2(G124), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(G33), .A2(G41), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n780), .C2(new_n812), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1206), .B2(KEYINPUT59), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1209), .A2(G50), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1207), .A2(new_n1211), .B1(new_n1191), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1200), .A2(new_n1201), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n764), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n759), .B1(new_n202), .B2(new_n832), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n1174), .C2(new_n761), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1190), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1189), .A2(new_n1218), .ZN(G375));
  AOI21_X1  g1019(.A(new_n759), .B1(new_n255), .B2(new_n832), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n805), .A2(new_n1148), .B1(new_n793), .B2(G150), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n787), .A2(G132), .B1(new_n795), .B2(G137), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1017), .A2(G159), .B1(G128), .B2(new_n797), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT122), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G50), .C2(new_n791), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1192), .A2(new_n396), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT121), .Z(new_n1228));
  OAI22_X1  g1028(.A1(new_n777), .A2(new_n205), .B1(new_n786), .B2(new_n851), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1010), .A2(new_n1037), .A3(new_n1229), .A4(new_n309), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n795), .A2(G283), .B1(new_n797), .B2(G303), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n610), .B2(new_n783), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1012), .B2(G107), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1226), .A2(new_n1228), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1220), .B1(new_n1234), .B2(new_n834), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1101), .B2(new_n760), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1115), .B2(new_n757), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1132), .A2(new_n979), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1115), .B1(new_n1093), .B2(new_n1116), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(G381));
  INV_X1    g1040(.A(G390), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n859), .ZN(new_n1242));
  OR4_X1    g1042(.A1(G396), .A2(new_n1242), .A3(G387), .A4(G393), .ZN(new_n1243));
  OR4_X1    g1043(.A1(G378), .A2(new_n1243), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1044(.A(G378), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n693), .A2(G213), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G407), .B(G213), .C1(G375), .C2(new_n1248), .ZN(G409));
  NOR2_X1   g1049(.A1(new_n1241), .A2(G387), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G390), .B1(new_n998), .B2(new_n1023), .ZN(new_n1251));
  XOR2_X1   g1051(.A(G393), .B(G396), .Z(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1253), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1239), .B1(KEYINPUT60), .B2(new_n1117), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1257), .A2(KEYINPUT125), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n710), .B1(new_n1239), .B2(KEYINPUT60), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1257), .B2(KEYINPUT125), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1237), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n859), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G384), .B(new_n1237), .C1(new_n1258), .C2(new_n1260), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(KEYINPUT62), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n979), .B1(new_n1135), .B2(new_n1180), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1179), .A2(new_n1265), .A3(new_n1183), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1217), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1173), .A2(new_n1178), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1268), .B2(new_n757), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G378), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT123), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1189), .A2(G378), .A3(new_n1218), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1247), .B(new_n1264), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT123), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1274), .B(G378), .C1(new_n1266), .C2(new_n1269), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT123), .B1(new_n1276), .B2(new_n1245), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1189), .A2(G378), .A3(new_n1218), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT124), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1262), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1263), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1272), .B(new_n1284), .C1(new_n1277), .C2(new_n1275), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1280), .A2(new_n1246), .A3(new_n1283), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1273), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1283), .B1(G2897), .B2(new_n1247), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1247), .A2(G2897), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1281), .A2(new_n1282), .A3(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1247), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1289), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1256), .B1(new_n1288), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1280), .A2(new_n1246), .A3(new_n1285), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1292), .B2(new_n1290), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1286), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1294), .A2(KEYINPUT63), .A3(new_n1283), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1256), .A2(KEYINPUT61), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1298), .A2(new_n1300), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1296), .A2(new_n1303), .ZN(G405));
  NAND2_X1  g1104(.A1(G375), .A2(new_n1245), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1272), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1283), .A2(new_n1307), .ZN(new_n1308));
  XOR2_X1   g1108(.A(new_n1306), .B(new_n1308), .Z(new_n1309));
  XNOR2_X1  g1109(.A(new_n1309), .B(new_n1256), .ZN(G402));
endmodule


