

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U556 ( .A(n763), .B(KEYINPUT98), .ZN(n777) );
  OR2_X1 U557 ( .A1(n732), .A2(n703), .ZN(n704) );
  AND2_X1 U558 ( .A1(G138), .A2(n899), .ZN(n571) );
  NOR2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n563) );
  NOR2_X4 U560 ( .A1(n701), .A2(G1384), .ZN(n789) );
  NAND2_X1 U561 ( .A1(n522), .A2(n820), .ZN(n837) );
  NAND2_X1 U562 ( .A1(n524), .A2(n523), .ZN(n522) );
  INV_X1 U563 ( .A(n786), .ZN(n523) );
  INV_X1 U564 ( .A(n787), .ZN(n524) );
  NAND2_X1 U565 ( .A1(n715), .A2(n876), .ZN(n714) );
  NOR2_X1 U566 ( .A1(n708), .A2(n709), .ZN(n715) );
  NAND2_X2 U567 ( .A1(G8), .A2(n747), .ZN(n785) );
  XNOR2_X1 U568 ( .A(n730), .B(n729), .ZN(n736) );
  NOR2_X2 U569 ( .A1(G651), .A2(n535), .ZN(n585) );
  NOR2_X2 U570 ( .A1(G2104), .A2(n556), .ZN(n565) );
  AND2_X1 U571 ( .A1(n987), .A2(n834), .ZN(n525) );
  OR2_X1 U572 ( .A1(n876), .A2(n715), .ZN(n716) );
  INV_X1 U573 ( .A(KEYINPUT29), .ZN(n729) );
  INV_X1 U574 ( .A(KEYINPUT31), .ZN(n743) );
  INV_X1 U575 ( .A(KEYINPUT66), .ZN(n537) );
  NOR2_X1 U576 ( .A1(n525), .A2(n819), .ZN(n820) );
  NOR2_X1 U577 ( .A1(G543), .A2(n536), .ZN(n530) );
  NOR2_X1 U578 ( .A1(G543), .A2(G651), .ZN(n660) );
  INV_X1 U579 ( .A(KEYINPUT0), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n526), .A2(G543), .ZN(n529) );
  INV_X1 U581 ( .A(G543), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n527), .A2(KEYINPUT0), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n529), .A2(n528), .ZN(n535) );
  NAND2_X1 U584 ( .A1(G51), .A2(n585), .ZN(n532) );
  INV_X1 U585 ( .A(G651), .ZN(n536) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n530), .Z(n664) );
  NAND2_X1 U587 ( .A1(G63), .A2(n664), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U589 ( .A(KEYINPUT6), .B(n533), .ZN(n544) );
  NAND2_X1 U590 ( .A1(n660), .A2(G89), .ZN(n534) );
  XNOR2_X1 U591 ( .A(n534), .B(KEYINPUT4), .ZN(n540) );
  OR2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n538) );
  XNOR2_X2 U593 ( .A(n538), .B(n537), .ZN(n665) );
  NAND2_X1 U594 ( .A1(G76), .A2(n665), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U596 ( .A(KEYINPUT5), .B(n541), .ZN(n542) );
  XNOR2_X1 U597 ( .A(KEYINPUT77), .B(n542), .ZN(n543) );
  NOR2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U599 ( .A(KEYINPUT7), .B(n545), .Z(G168) );
  XOR2_X1 U600 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  INV_X1 U605 ( .A(G120), .ZN(G236) );
  NAND2_X1 U606 ( .A1(G52), .A2(n585), .ZN(n546) );
  XNOR2_X1 U607 ( .A(n546), .B(KEYINPUT69), .ZN(n553) );
  NAND2_X1 U608 ( .A1(G90), .A2(n660), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G77), .A2(n665), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U611 ( .A(n549), .B(KEYINPUT9), .ZN(n551) );
  NAND2_X1 U612 ( .A1(G64), .A2(n664), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U614 ( .A1(n553), .A2(n552), .ZN(G171) );
  INV_X1 U615 ( .A(G171), .ZN(G301) );
  INV_X1 U616 ( .A(G2105), .ZN(n556) );
  AND2_X1 U617 ( .A1(G2105), .A2(G2104), .ZN(n903) );
  NAND2_X1 U618 ( .A1(G113), .A2(n903), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G125), .A2(n565), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n695) );
  AND2_X1 U621 ( .A1(G2104), .A2(n556), .ZN(n557) );
  XNOR2_X2 U622 ( .A(n557), .B(KEYINPUT64), .ZN(n900) );
  NAND2_X1 U623 ( .A1(n900), .A2(G101), .ZN(n559) );
  INV_X1 U624 ( .A(n559), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n558), .A2(KEYINPUT23), .ZN(n562) );
  INV_X1 U626 ( .A(KEYINPUT23), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n700) );
  XOR2_X2 U629 ( .A(KEYINPUT17), .B(n563), .Z(n899) );
  NAND2_X1 U630 ( .A1(n899), .A2(G137), .ZN(n697) );
  NAND2_X1 U631 ( .A1(n700), .A2(n697), .ZN(n564) );
  NOR2_X1 U632 ( .A1(n695), .A2(n564), .ZN(G160) );
  NAND2_X1 U633 ( .A1(G102), .A2(n900), .ZN(n569) );
  NAND2_X1 U634 ( .A1(G114), .A2(n903), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G126), .A2(n565), .ZN(n566) );
  AND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n701) );
  BUF_X1 U639 ( .A(n701), .Z(G164) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n572) );
  XOR2_X1 U641 ( .A(n572), .B(KEYINPUT10), .Z(n851) );
  NAND2_X1 U642 ( .A1(n851), .A2(G567), .ZN(n573) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  NAND2_X1 U644 ( .A1(n665), .A2(G68), .ZN(n574) );
  XNOR2_X1 U645 ( .A(KEYINPUT72), .B(n574), .ZN(n577) );
  NAND2_X1 U646 ( .A1(n660), .A2(G81), .ZN(n575) );
  XNOR2_X1 U647 ( .A(KEYINPUT12), .B(n575), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U649 ( .A(n578), .B(KEYINPUT13), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n664), .A2(G56), .ZN(n579) );
  XNOR2_X1 U651 ( .A(KEYINPUT14), .B(n579), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U653 ( .A(n582), .B(KEYINPUT73), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G43), .A2(n585), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n709) );
  INV_X1 U656 ( .A(n709), .ZN(n1002) );
  XNOR2_X1 U657 ( .A(G860), .B(KEYINPUT74), .ZN(n608) );
  NAND2_X1 U658 ( .A1(n1002), .A2(n608), .ZN(G153) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n585), .A2(G54), .ZN(n586) );
  XOR2_X1 U661 ( .A(KEYINPUT75), .B(n586), .Z(n588) );
  NAND2_X1 U662 ( .A1(G79), .A2(n665), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U664 ( .A(KEYINPUT76), .B(n589), .ZN(n593) );
  NAND2_X1 U665 ( .A1(G66), .A2(n664), .ZN(n591) );
  NAND2_X1 U666 ( .A1(G92), .A2(n660), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U669 ( .A(KEYINPUT15), .B(n594), .ZN(n999) );
  INV_X1 U670 ( .A(G868), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n999), .A2(n605), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(G284) );
  NAND2_X1 U673 ( .A1(n665), .A2(G78), .ZN(n597) );
  XOR2_X1 U674 ( .A(KEYINPUT70), .B(n597), .Z(n602) );
  NAND2_X1 U675 ( .A1(G53), .A2(n585), .ZN(n599) );
  NAND2_X1 U676 ( .A1(G65), .A2(n664), .ZN(n598) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U678 ( .A(KEYINPUT71), .B(n600), .Z(n601) );
  NOR2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n660), .A2(G91), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(G299) );
  NOR2_X1 U682 ( .A1(G286), .A2(n605), .ZN(n607) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(G297) );
  INV_X1 U685 ( .A(G559), .ZN(n609) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n999), .A2(n610), .ZN(n611) );
  XOR2_X1 U688 ( .A(KEYINPUT16), .B(n611), .Z(G148) );
  NOR2_X1 U689 ( .A1(G868), .A2(n709), .ZN(n614) );
  INV_X1 U690 ( .A(n999), .ZN(n876) );
  NAND2_X1 U691 ( .A1(n876), .A2(G868), .ZN(n612) );
  NOR2_X1 U692 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U694 ( .A(KEYINPUT78), .B(n615), .ZN(G282) );
  XOR2_X1 U695 ( .A(G2100), .B(KEYINPUT80), .Z(n625) );
  NAND2_X1 U696 ( .A1(G111), .A2(n903), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G135), .A2(n899), .ZN(n617) );
  NAND2_X1 U698 ( .A1(G99), .A2(n900), .ZN(n616) );
  NAND2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n565), .A2(G123), .ZN(n618) );
  XOR2_X1 U701 ( .A(KEYINPUT18), .B(n618), .Z(n619) );
  NOR2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n623), .B(KEYINPUT79), .ZN(n949) );
  XNOR2_X1 U705 ( .A(G2096), .B(n949), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(G156) );
  XOR2_X1 U707 ( .A(n1002), .B(KEYINPUT81), .Z(n627) );
  NAND2_X1 U708 ( .A1(G559), .A2(n876), .ZN(n626) );
  XOR2_X1 U709 ( .A(n627), .B(n626), .Z(n677) );
  NOR2_X1 U710 ( .A1(n677), .A2(G860), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G55), .A2(n585), .ZN(n629) );
  NAND2_X1 U712 ( .A1(G67), .A2(n664), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G93), .A2(n660), .ZN(n631) );
  NAND2_X1 U715 ( .A1(G80), .A2(n665), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n671) );
  XNOR2_X1 U718 ( .A(n634), .B(n671), .ZN(G145) );
  NAND2_X1 U719 ( .A1(n664), .A2(G60), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G72), .A2(n665), .ZN(n637) );
  NAND2_X1 U721 ( .A1(G47), .A2(n585), .ZN(n635) );
  XOR2_X1 U722 ( .A(KEYINPUT67), .B(n635), .Z(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G85), .A2(n660), .ZN(n638) );
  XNOR2_X1 U725 ( .A(KEYINPUT65), .B(n638), .ZN(n639) );
  NOR2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U728 ( .A(n643), .B(KEYINPUT68), .ZN(G290) );
  NAND2_X1 U729 ( .A1(G48), .A2(n585), .ZN(n645) );
  NAND2_X1 U730 ( .A1(G86), .A2(n660), .ZN(n644) );
  NAND2_X1 U731 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U732 ( .A1(n665), .A2(G73), .ZN(n646) );
  XOR2_X1 U733 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  NOR2_X1 U734 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n664), .A2(G61), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(G305) );
  NAND2_X1 U737 ( .A1(n585), .A2(G49), .ZN(n651) );
  XNOR2_X1 U738 ( .A(n651), .B(KEYINPUT82), .ZN(n653) );
  NAND2_X1 U739 ( .A1(G74), .A2(G651), .ZN(n652) );
  NAND2_X1 U740 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U741 ( .A(KEYINPUT83), .B(n654), .ZN(n658) );
  NAND2_X1 U742 ( .A1(G87), .A2(n535), .ZN(n655) );
  XOR2_X1 U743 ( .A(KEYINPUT84), .B(n655), .Z(n656) );
  NOR2_X1 U744 ( .A1(n664), .A2(n656), .ZN(n657) );
  NAND2_X1 U745 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U746 ( .A(KEYINPUT85), .B(n659), .Z(G288) );
  NAND2_X1 U747 ( .A1(G88), .A2(n660), .ZN(n661) );
  XNOR2_X1 U748 ( .A(n661), .B(KEYINPUT86), .ZN(n663) );
  NAND2_X1 U749 ( .A1(n585), .A2(G50), .ZN(n662) );
  NAND2_X1 U750 ( .A1(n663), .A2(n662), .ZN(n669) );
  NAND2_X1 U751 ( .A1(n664), .A2(G62), .ZN(n667) );
  NAND2_X1 U752 ( .A1(G75), .A2(n665), .ZN(n666) );
  NAND2_X1 U753 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U754 ( .A1(n669), .A2(n668), .ZN(G166) );
  INV_X1 U755 ( .A(G166), .ZN(G303) );
  NOR2_X1 U756 ( .A1(G868), .A2(n671), .ZN(n670) );
  XNOR2_X1 U757 ( .A(n670), .B(KEYINPUT87), .ZN(n680) );
  XNOR2_X1 U758 ( .A(n671), .B(G305), .ZN(n672) );
  XNOR2_X1 U759 ( .A(n672), .B(G288), .ZN(n673) );
  XOR2_X1 U760 ( .A(n673), .B(KEYINPUT19), .Z(n675) );
  INV_X1 U761 ( .A(G299), .ZN(n724) );
  XOR2_X1 U762 ( .A(G303), .B(n724), .Z(n674) );
  XNOR2_X1 U763 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U764 ( .A(G290), .B(n676), .ZN(n879) );
  XOR2_X1 U765 ( .A(n677), .B(n879), .Z(n678) );
  NAND2_X1 U766 ( .A1(G868), .A2(n678), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n680), .A2(n679), .ZN(G295) );
  XOR2_X1 U768 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n682) );
  NAND2_X1 U769 ( .A1(G2084), .A2(G2078), .ZN(n681) );
  XNOR2_X1 U770 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U771 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U772 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U774 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U775 ( .A1(G236), .A2(G237), .ZN(n686) );
  NAND2_X1 U776 ( .A1(G69), .A2(n686), .ZN(n687) );
  XNOR2_X1 U777 ( .A(KEYINPUT89), .B(n687), .ZN(n688) );
  NAND2_X1 U778 ( .A1(n688), .A2(G108), .ZN(n855) );
  NAND2_X1 U779 ( .A1(G567), .A2(n855), .ZN(n693) );
  NOR2_X1 U780 ( .A1(G220), .A2(G219), .ZN(n689) );
  XOR2_X1 U781 ( .A(KEYINPUT22), .B(n689), .Z(n690) );
  NOR2_X1 U782 ( .A1(G218), .A2(n690), .ZN(n691) );
  NAND2_X1 U783 ( .A1(G96), .A2(n691), .ZN(n856) );
  NAND2_X1 U784 ( .A1(G2106), .A2(n856), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n857) );
  NAND2_X1 U786 ( .A1(G483), .A2(G661), .ZN(n694) );
  NOR2_X1 U787 ( .A1(n857), .A2(n694), .ZN(n854) );
  NAND2_X1 U788 ( .A1(n854), .A2(G36), .ZN(G176) );
  INV_X1 U789 ( .A(G40), .ZN(n696) );
  NOR2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n698) );
  AND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n790) );
  INV_X1 U793 ( .A(n789), .ZN(n702) );
  NOR2_X4 U794 ( .A1(n790), .A2(n702), .ZN(n732) );
  INV_X1 U795 ( .A(G1341), .ZN(n703) );
  XNOR2_X1 U796 ( .A(n704), .B(KEYINPUT96), .ZN(n707) );
  NAND2_X1 U797 ( .A1(G1996), .A2(n732), .ZN(n705) );
  XNOR2_X1 U798 ( .A(KEYINPUT26), .B(n705), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n708) );
  INV_X1 U800 ( .A(n732), .ZN(n747) );
  AND2_X1 U801 ( .A1(n747), .A2(G1348), .ZN(n710) );
  XNOR2_X1 U802 ( .A(n710), .B(KEYINPUT97), .ZN(n712) );
  NAND2_X1 U803 ( .A1(n732), .A2(G2067), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n722) );
  NAND2_X1 U807 ( .A1(n732), .A2(G2072), .ZN(n718) );
  XNOR2_X1 U808 ( .A(n718), .B(KEYINPUT27), .ZN(n720) );
  XOR2_X1 U809 ( .A(G1956), .B(KEYINPUT94), .Z(n1010) );
  NOR2_X1 U810 ( .A1(n732), .A2(n1010), .ZN(n719) );
  NOR2_X1 U811 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n721) );
  NAND2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n728) );
  NOR2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n726) );
  XNOR2_X1 U815 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n725) );
  XNOR2_X1 U816 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n730) );
  OR2_X1 U818 ( .A1(n732), .A2(G1961), .ZN(n734) );
  XOR2_X1 U819 ( .A(G2078), .B(KEYINPUT25), .Z(n731) );
  XNOR2_X1 U820 ( .A(KEYINPUT93), .B(n731), .ZN(n964) );
  NAND2_X1 U821 ( .A1(n732), .A2(n964), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n740) );
  NAND2_X1 U823 ( .A1(n740), .A2(G171), .ZN(n735) );
  NAND2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n746) );
  NOR2_X1 U825 ( .A1(G1966), .A2(n785), .ZN(n758) );
  NOR2_X1 U826 ( .A1(G2084), .A2(n747), .ZN(n755) );
  NOR2_X1 U827 ( .A1(n758), .A2(n755), .ZN(n737) );
  NAND2_X1 U828 ( .A1(G8), .A2(n737), .ZN(n738) );
  XNOR2_X1 U829 ( .A(KEYINPUT30), .B(n738), .ZN(n739) );
  NOR2_X1 U830 ( .A1(G168), .A2(n739), .ZN(n742) );
  NOR2_X1 U831 ( .A1(G171), .A2(n740), .ZN(n741) );
  NOR2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n744) );
  XNOR2_X1 U833 ( .A(n744), .B(n743), .ZN(n745) );
  NAND2_X1 U834 ( .A1(n746), .A2(n745), .ZN(n756) );
  NAND2_X1 U835 ( .A1(n756), .A2(G286), .ZN(n752) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n785), .ZN(n749) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n750), .A2(G303), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n753), .A2(G8), .ZN(n754) );
  XNOR2_X1 U842 ( .A(n754), .B(KEYINPUT32), .ZN(n762) );
  NAND2_X1 U843 ( .A1(G8), .A2(n755), .ZN(n760) );
  INV_X1 U844 ( .A(n756), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U847 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U848 ( .A1(G1971), .A2(G303), .ZN(n764) );
  NOR2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n982) );
  NOR2_X1 U850 ( .A1(n764), .A2(n982), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n777), .A2(n765), .ZN(n767) );
  NAND2_X1 U852 ( .A1(G288), .A2(G1976), .ZN(n766) );
  XOR2_X1 U853 ( .A(KEYINPUT99), .B(n766), .Z(n983) );
  NAND2_X1 U854 ( .A1(n767), .A2(n983), .ZN(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(KEYINPUT100), .ZN(n769) );
  NOR2_X1 U856 ( .A1(n769), .A2(n785), .ZN(n770) );
  NOR2_X1 U857 ( .A1(KEYINPUT33), .A2(n770), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n982), .A2(KEYINPUT33), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n785), .A2(n771), .ZN(n772) );
  NOR2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n994) );
  NAND2_X1 U862 ( .A1(n774), .A2(n994), .ZN(n781) );
  NOR2_X1 U863 ( .A1(G2090), .A2(G303), .ZN(n775) );
  XOR2_X1 U864 ( .A(KEYINPUT101), .B(n775), .Z(n776) );
  NAND2_X1 U865 ( .A1(G8), .A2(n776), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n779), .A2(n785), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U869 ( .A(n782), .B(KEYINPUT102), .ZN(n787) );
  NOR2_X1 U870 ( .A1(G1981), .A2(G305), .ZN(n783) );
  XOR2_X1 U871 ( .A(n783), .B(KEYINPUT24), .Z(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U873 ( .A(G1986), .B(G290), .ZN(n987) );
  NOR2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n834) );
  XNOR2_X1 U875 ( .A(G2067), .B(KEYINPUT37), .ZN(n822) );
  NAND2_X1 U876 ( .A1(G140), .A2(n899), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G104), .A2(n900), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U879 ( .A(KEYINPUT34), .B(n793), .ZN(n799) );
  NAND2_X1 U880 ( .A1(G116), .A2(n903), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G128), .A2(n565), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U883 ( .A(KEYINPUT35), .B(n796), .Z(n797) );
  XNOR2_X1 U884 ( .A(KEYINPUT90), .B(n797), .ZN(n798) );
  NOR2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U886 ( .A(KEYINPUT36), .B(n800), .ZN(n922) );
  NOR2_X1 U887 ( .A1(n822), .A2(n922), .ZN(n933) );
  NAND2_X1 U888 ( .A1(n834), .A2(n933), .ZN(n831) );
  NAND2_X1 U889 ( .A1(G131), .A2(n899), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G95), .A2(n900), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U892 ( .A(KEYINPUT92), .B(n803), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G119), .A2(n565), .ZN(n804) );
  XNOR2_X1 U894 ( .A(KEYINPUT91), .B(n804), .ZN(n805) );
  NOR2_X1 U895 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U896 ( .A1(n903), .A2(G107), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n808), .A2(n807), .ZN(n915) );
  AND2_X1 U898 ( .A1(n915), .A2(G1991), .ZN(n817) );
  NAND2_X1 U899 ( .A1(G117), .A2(n903), .ZN(n810) );
  NAND2_X1 U900 ( .A1(G129), .A2(n565), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n900), .A2(G105), .ZN(n811) );
  XOR2_X1 U903 ( .A(KEYINPUT38), .B(n811), .Z(n812) );
  NOR2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n899), .A2(G141), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n909) );
  AND2_X1 U907 ( .A1(G1996), .A2(n909), .ZN(n816) );
  NOR2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n943) );
  INV_X1 U909 ( .A(n943), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n818), .A2(n834), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n831), .A2(n823), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n822), .A2(n922), .ZN(n935) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n909), .ZN(n945) );
  INV_X1 U914 ( .A(n823), .ZN(n827) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n915), .ZN(n824) );
  XOR2_X1 U916 ( .A(KEYINPUT103), .B(n824), .Z(n950) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n825) );
  NOR2_X1 U918 ( .A1(n950), .A2(n825), .ZN(n826) );
  NOR2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U920 ( .A1(n945), .A2(n828), .ZN(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT39), .B(n829), .ZN(n830) );
  XNOR2_X1 U922 ( .A(n830), .B(KEYINPUT104), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U924 ( .A1(n935), .A2(n833), .ZN(n835) );
  NAND2_X1 U925 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U926 ( .A1(n837), .A2(n836), .ZN(n839) );
  XOR2_X1 U927 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n838) );
  XNOR2_X1 U928 ( .A(n839), .B(n838), .ZN(G329) );
  XNOR2_X1 U929 ( .A(G2443), .B(G2446), .ZN(n849) );
  XOR2_X1 U930 ( .A(G2430), .B(KEYINPUT107), .Z(n841) );
  XNOR2_X1 U931 ( .A(G2454), .B(G2435), .ZN(n840) );
  XNOR2_X1 U932 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U933 ( .A(G2438), .B(G2427), .Z(n843) );
  XNOR2_X1 U934 ( .A(G1341), .B(G1348), .ZN(n842) );
  XNOR2_X1 U935 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U936 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U937 ( .A(G2451), .B(KEYINPUT106), .ZN(n846) );
  XNOR2_X1 U938 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U939 ( .A(n849), .B(n848), .ZN(n850) );
  NAND2_X1 U940 ( .A1(n850), .A2(G14), .ZN(n927) );
  XOR2_X1 U941 ( .A(KEYINPUT108), .B(n927), .Z(G401) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n851), .ZN(G217) );
  INV_X1 U943 ( .A(n851), .ZN(G223) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n852) );
  NAND2_X1 U945 ( .A1(G661), .A2(n852), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n853) );
  NAND2_X1 U947 ( .A1(n854), .A2(n853), .ZN(G188) );
  NOR2_X1 U948 ( .A1(n856), .A2(n855), .ZN(G325) );
  XNOR2_X1 U949 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U951 ( .A(G108), .ZN(G238) );
  INV_X1 U952 ( .A(G96), .ZN(G221) );
  XOR2_X1 U953 ( .A(KEYINPUT110), .B(n857), .Z(G319) );
  XOR2_X1 U954 ( .A(G2678), .B(G2084), .Z(n859) );
  XNOR2_X1 U955 ( .A(G2078), .B(G2072), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U957 ( .A(n860), .B(G2096), .Z(n862) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2090), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U960 ( .A(G2100), .B(KEYINPUT111), .Z(n864) );
  XNOR2_X1 U961 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U963 ( .A(n866), .B(n865), .Z(G227) );
  XOR2_X1 U964 ( .A(G1976), .B(G1961), .Z(n868) );
  XNOR2_X1 U965 ( .A(G1981), .B(G1966), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U967 ( .A(n869), .B(KEYINPUT41), .Z(n871) );
  XNOR2_X1 U968 ( .A(G1996), .B(G1991), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U970 ( .A(G2474), .B(G1971), .Z(n873) );
  XNOR2_X1 U971 ( .A(G1986), .B(G1956), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(G229) );
  XOR2_X1 U974 ( .A(n1002), .B(G286), .Z(n878) );
  XOR2_X1 U975 ( .A(G301), .B(n876), .Z(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n881) );
  NOR2_X1 U978 ( .A1(G37), .A2(n881), .ZN(G397) );
  NAND2_X1 U979 ( .A1(G100), .A2(n900), .ZN(n888) );
  NAND2_X1 U980 ( .A1(G136), .A2(n899), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G112), .A2(n903), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n886) );
  NAND2_X1 U983 ( .A1(n565), .A2(G124), .ZN(n884) );
  XOR2_X1 U984 ( .A(KEYINPUT44), .B(n884), .Z(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  NAND2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(KEYINPUT112), .B(n889), .Z(G162) );
  NAND2_X1 U988 ( .A1(G118), .A2(n903), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G130), .A2(n565), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n898) );
  XNOR2_X1 U991 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n896) );
  NAND2_X1 U992 ( .A1(G142), .A2(n899), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G106), .A2(n900), .ZN(n892) );
  NAND2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n894), .B(KEYINPUT45), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n914) );
  NAND2_X1 U998 ( .A1(G139), .A2(n899), .ZN(n902) );
  NAND2_X1 U999 ( .A1(G103), .A2(n900), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n908) );
  NAND2_X1 U1001 ( .A1(G115), .A2(n903), .ZN(n905) );
  NAND2_X1 U1002 ( .A1(G127), .A2(n565), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(KEYINPUT47), .B(n906), .Z(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n936) );
  XOR2_X1 U1006 ( .A(n936), .B(n949), .Z(n911) );
  XOR2_X1 U1007 ( .A(G160), .B(n909), .Z(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1009 ( .A(G162), .B(n912), .Z(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n924) );
  XOR2_X1 U1011 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n917) );
  XOR2_X1 U1012 ( .A(n915), .B(KEYINPUT116), .Z(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1014 ( .A(n918), .B(KEYINPUT46), .Z(n920) );
  XNOR2_X1 U1015 ( .A(G164), .B(KEYINPUT117), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n925), .ZN(n926) );
  XNOR2_X1 U1020 ( .A(KEYINPUT118), .B(n926), .ZN(G395) );
  NAND2_X1 U1021 ( .A1(G319), .A2(n927), .ZN(n930) );
  NOR2_X1 U1022 ( .A1(G227), .A2(G229), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(KEYINPUT49), .B(n928), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n932) );
  NOR2_X1 U1025 ( .A1(G397), .A2(G395), .ZN(n931) );
  NAND2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G69), .ZN(G235) );
  INV_X1 U1029 ( .A(n933), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n955) );
  XOR2_X1 U1031 ( .A(G2072), .B(n936), .Z(n938) );
  XOR2_X1 U1032 ( .A(G164), .B(G2078), .Z(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1034 ( .A(KEYINPUT50), .B(n939), .Z(n941) );
  XOR2_X1 U1035 ( .A(G160), .B(G2084), .Z(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n948) );
  XOR2_X1 U1038 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(n946), .B(KEYINPUT51), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n953) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1043 ( .A(KEYINPUT119), .B(n951), .Z(n952) );
  NAND2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1045 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n956), .ZN(n958) );
  INV_X1 U1047 ( .A(KEYINPUT55), .ZN(n957) );
  NAND2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1049 ( .A1(n959), .A2(G29), .ZN(n1039) );
  XNOR2_X1 U1050 ( .A(KEYINPUT54), .B(G34), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(n960), .B(KEYINPUT121), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G2084), .B(n961), .ZN(n977) );
  XNOR2_X1 U1053 ( .A(G2090), .B(G35), .ZN(n975) );
  XOR2_X1 U1054 ( .A(G2067), .B(G26), .Z(n963) );
  XOR2_X1 U1055 ( .A(G1991), .B(G25), .Z(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n972) );
  XNOR2_X1 U1057 ( .A(G27), .B(n964), .ZN(n970) );
  XOR2_X1 U1058 ( .A(G32), .B(G1996), .Z(n965) );
  NAND2_X1 U1059 ( .A1(n965), .A2(G28), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(KEYINPUT120), .B(G2072), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G33), .B(n966), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n973), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1068 ( .A(KEYINPUT55), .B(n978), .Z(n980) );
  INV_X1 U1069 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n981), .ZN(n1037) );
  INV_X1 U1072 ( .A(G16), .ZN(n1033) );
  XOR2_X1 U1073 ( .A(n1033), .B(KEYINPUT56), .Z(n1008) );
  INV_X1 U1074 ( .A(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1076 ( .A(KEYINPUT123), .B(n985), .Z(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G299), .B(G1956), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(G303), .B(G1971), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n992), .B(KEYINPUT124), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G168), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT122), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1086 ( .A(KEYINPUT57), .B(n996), .Z(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1006) );
  XOR2_X1 U1088 ( .A(n999), .B(G1348), .Z(n1001) );
  XOR2_X1 U1089 ( .A(G301), .B(G1961), .Z(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(G1341), .B(n1002), .Z(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1035) );
  XNOR2_X1 U1095 ( .A(KEYINPUT125), .B(G1966), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1009), .B(G21), .ZN(n1022) );
  XNOR2_X1 U1097 ( .A(n1010), .B(G20), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G1341), .B(G19), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(KEYINPUT59), .B(G1348), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(G4), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1018), .Z(n1020) );
  XNOR2_X1 U1106 ( .A(G1961), .B(G5), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1030) );
  XOR2_X1 U1109 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n1028) );
  XOR2_X1 U1110 ( .A(G1986), .B(G24), .Z(n1026) );
  XNOR2_X1 U1111 ( .A(G1971), .B(G22), .ZN(n1024) );
  XNOR2_X1 U1112 ( .A(G23), .B(G1976), .ZN(n1023) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1115 ( .A(n1028), .B(n1027), .Z(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(KEYINPUT61), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1120 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1121 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1122 ( .A(n1040), .B(KEYINPUT127), .ZN(n1041) );
  XOR2_X1 U1123 ( .A(KEYINPUT62), .B(n1041), .Z(G150) );
  INV_X1 U1124 ( .A(G150), .ZN(G311) );
endmodule

