

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743;

  OR2_X1 U377 ( .A1(n687), .A2(n551), .ZN(n504) );
  BUF_X1 U378 ( .A(n662), .Z(n357) );
  XNOR2_X1 U379 ( .A(n570), .B(n414), .ZN(n662) );
  AND2_X1 U380 ( .A1(n379), .A2(n585), .ZN(n569) );
  OR2_X1 U381 ( .A1(n699), .A2(G902), .ZN(n415) );
  XNOR2_X1 U382 ( .A(n524), .B(n458), .ZN(n494) );
  BUF_X1 U383 ( .A(G143), .Z(n358) );
  XNOR2_X1 U384 ( .A(n491), .B(n718), .ZN(n426) );
  XNOR2_X2 U385 ( .A(n722), .B(n484), .ZN(n491) );
  AND2_X2 U386 ( .A1(n641), .A2(n595), .ZN(n596) );
  XNOR2_X1 U387 ( .A(G113), .B(n358), .ZN(n511) );
  XNOR2_X1 U388 ( .A(n605), .B(n604), .ZN(n619) );
  NOR2_X1 U389 ( .A1(n538), .A2(n539), .ZN(n544) );
  INV_X2 U390 ( .A(G953), .ZN(n560) );
  AND2_X1 U391 ( .A1(n740), .A2(KEYINPUT84), .ZN(n359) );
  XNOR2_X2 U392 ( .A(n432), .B(n611), .ZN(n448) );
  XNOR2_X2 U393 ( .A(n388), .B(n387), .ZN(n740) );
  XNOR2_X2 U394 ( .A(n728), .B(G146), .ZN(n485) );
  NOR2_X2 U395 ( .A1(n416), .A2(n737), .ZN(n543) );
  XNOR2_X2 U396 ( .A(n421), .B(KEYINPUT35), .ZN(n737) );
  XNOR2_X1 U397 ( .A(n594), .B(KEYINPUT105), .ZN(n738) );
  AND2_X1 U398 ( .A1(n431), .A2(n680), .ZN(n605) );
  NOR2_X2 U399 ( .A1(n705), .A2(G902), .ZN(n480) );
  XOR2_X1 U400 ( .A(G146), .B(G125), .Z(n492) );
  NOR2_X1 U401 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U402 ( .A1(KEYINPUT77), .A2(n596), .ZN(n597) );
  NOR2_X1 U403 ( .A1(n540), .A2(n537), .ZN(n637) );
  AND2_X1 U404 ( .A1(n591), .A2(n590), .ZN(n431) );
  NAND2_X1 U405 ( .A1(n571), .A2(n430), .ZN(n429) );
  BUF_X1 U406 ( .A(n592), .Z(n617) );
  XOR2_X1 U407 ( .A(n481), .B(n480), .Z(n540) );
  XNOR2_X1 U408 ( .A(n407), .B(G110), .ZN(n490) );
  XOR2_X1 U409 ( .A(G113), .B(G116), .Z(n367) );
  INV_X1 U410 ( .A(KEYINPUT80), .ZN(n385) );
  XNOR2_X1 U411 ( .A(n569), .B(n568), .ZN(n389) );
  OR2_X2 U412 ( .A1(n625), .A2(G902), .ZN(n489) );
  XNOR2_X1 U413 ( .A(n518), .B(n517), .ZN(n519) );
  NOR2_X1 U414 ( .A1(n359), .A2(n360), .ZN(n420) );
  INV_X1 U415 ( .A(KEYINPUT4), .ZN(n458) );
  NOR2_X1 U416 ( .A1(G953), .A2(G237), .ZN(n507) );
  XNOR2_X1 U417 ( .A(n411), .B(G140), .ZN(n478) );
  INV_X1 U418 ( .A(G137), .ZN(n411) );
  XNOR2_X1 U419 ( .A(n376), .B(n375), .ZN(n521) );
  INV_X1 U420 ( .A(KEYINPUT8), .ZN(n375) );
  NAND2_X1 U421 ( .A1(n560), .A2(G234), .ZN(n376) );
  NAND2_X1 U422 ( .A1(G234), .A2(G237), .ZN(n503) );
  XNOR2_X1 U423 ( .A(n392), .B(n391), .ZN(n687) );
  INV_X1 U424 ( .A(KEYINPUT33), .ZN(n391) );
  XNOR2_X1 U425 ( .A(n535), .B(KEYINPUT22), .ZN(n538) );
  NOR2_X1 U426 ( .A1(n601), .A2(n602), .ZN(n435) );
  NAND2_X1 U427 ( .A1(n383), .A2(n433), .ZN(n432) );
  XNOR2_X1 U428 ( .A(n434), .B(KEYINPUT46), .ZN(n433) );
  XNOR2_X1 U429 ( .A(n435), .B(n603), .ZN(n383) );
  NOR2_X1 U430 ( .A1(n743), .A2(n741), .ZN(n434) );
  NOR2_X1 U431 ( .A1(n629), .A2(n556), .ZN(n557) );
  NOR2_X1 U432 ( .A1(n555), .A2(n684), .ZN(n556) );
  NOR2_X1 U433 ( .A1(n634), .A2(n645), .ZN(n555) );
  XNOR2_X1 U434 ( .A(n467), .B(KEYINPUT91), .ZN(n665) );
  XNOR2_X1 U435 ( .A(KEYINPUT88), .B(KEYINPUT23), .ZN(n473) );
  XNOR2_X1 U436 ( .A(G119), .B(G128), .ZN(n471) );
  INV_X1 U437 ( .A(G122), .ZN(n525) );
  XOR2_X1 U438 ( .A(G134), .B(KEYINPUT9), .Z(n523) );
  XOR2_X1 U439 ( .A(G902), .B(KEYINPUT15), .Z(n624) );
  OR2_X2 U440 ( .A1(n729), .A2(n715), .ZN(n452) );
  XNOR2_X1 U441 ( .A(n516), .B(n515), .ZN(n701) );
  XNOR2_X1 U442 ( .A(n408), .B(n490), .ZN(n461) );
  XNOR2_X1 U443 ( .A(n393), .B(n364), .ZN(n497) );
  NAND2_X1 U444 ( .A1(n380), .A2(n381), .ZN(n655) );
  NOR2_X1 U445 ( .A1(n623), .A2(n451), .ZN(n381) );
  BUF_X1 U446 ( .A(n622), .Z(n623) );
  INV_X1 U447 ( .A(n377), .ZN(n606) );
  XNOR2_X1 U448 ( .A(n581), .B(KEYINPUT103), .ZN(n612) );
  INV_X1 U449 ( .A(KEYINPUT0), .ZN(n428) );
  AND2_X1 U450 ( .A1(n502), .A2(n363), .ZN(n430) );
  XNOR2_X1 U451 ( .A(n554), .B(KEYINPUT95), .ZN(n675) );
  XNOR2_X1 U452 ( .A(n531), .B(G478), .ZN(n549) );
  NAND2_X1 U453 ( .A1(n548), .A2(n549), .ZN(n377) );
  INV_X1 U454 ( .A(KEYINPUT1), .ZN(n414) );
  XNOR2_X1 U455 ( .A(n491), .B(n439), .ZN(n443) );
  XNOR2_X1 U456 ( .A(n442), .B(n440), .ZN(n439) );
  XNOR2_X1 U457 ( .A(n486), .B(n441), .ZN(n440) );
  AND2_X1 U458 ( .A1(n660), .A2(n560), .ZN(n438) );
  XNOR2_X1 U459 ( .A(n738), .B(KEYINPUT78), .ZN(n599) );
  OR2_X1 U460 ( .A1(G237), .A2(G902), .ZN(n500) );
  XNOR2_X1 U461 ( .A(n494), .B(n361), .ZN(n728) );
  XOR2_X1 U462 ( .A(G140), .B(G131), .Z(n512) );
  XOR2_X1 U463 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n509) );
  XNOR2_X1 U464 ( .A(n478), .B(n409), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n410), .B(G104), .ZN(n409) );
  INV_X1 U466 ( .A(KEYINPUT72), .ZN(n410) );
  XNOR2_X1 U467 ( .A(KEYINPUT64), .B(G101), .ZN(n484) );
  XNOR2_X1 U468 ( .A(G107), .B(KEYINPUT86), .ZN(n407) );
  XOR2_X1 U469 ( .A(KEYINPUT18), .B(KEYINPUT73), .Z(n496) );
  XNOR2_X1 U470 ( .A(KEYINPUT17), .B(KEYINPUT85), .ZN(n495) );
  XNOR2_X1 U471 ( .A(n494), .B(n493), .ZN(n393) );
  INV_X1 U472 ( .A(n742), .ZN(n447) );
  INV_X1 U473 ( .A(n665), .ZN(n532) );
  INV_X1 U474 ( .A(KEYINPUT5), .ZN(n441) );
  XNOR2_X1 U475 ( .A(n487), .B(n488), .ZN(n442) );
  XOR2_X1 U476 ( .A(KEYINPUT93), .B(KEYINPUT70), .Z(n487) );
  XNOR2_X1 U477 ( .A(n608), .B(n395), .ZN(n678) );
  XNOR2_X1 U478 ( .A(n607), .B(n396), .ZN(n395) );
  INV_X1 U479 ( .A(KEYINPUT108), .ZN(n396) );
  XNOR2_X1 U480 ( .A(n587), .B(n586), .ZN(n591) );
  INV_X1 U481 ( .A(KEYINPUT30), .ZN(n586) );
  NAND2_X1 U482 ( .A1(n450), .A2(n449), .ZN(n453) );
  AND2_X1 U483 ( .A1(n655), .A2(n374), .ZN(n449) );
  XNOR2_X1 U484 ( .A(KEYINPUT3), .B(G119), .ZN(n483) );
  XNOR2_X1 U485 ( .A(n390), .B(n362), .ZN(n479) );
  XNOR2_X1 U486 ( .A(n476), .B(n475), .ZN(n390) );
  XNOR2_X1 U487 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U488 ( .A(n445), .B(n444), .ZN(n741) );
  XNOR2_X1 U489 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n444) );
  AND2_X1 U490 ( .A1(n612), .A2(n378), .ZN(n583) );
  XNOR2_X1 U491 ( .A(n504), .B(n370), .ZN(n422) );
  INV_X1 U492 ( .A(KEYINPUT32), .ZN(n387) );
  XNOR2_X1 U493 ( .A(n413), .B(n412), .ZN(n645) );
  XNOR2_X1 U494 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n412) );
  NOR2_X1 U495 ( .A1(n538), .A2(n614), .ZN(n536) );
  XNOR2_X1 U496 ( .A(n377), .B(KEYINPUT101), .ZN(n643) );
  XNOR2_X1 U497 ( .A(n382), .B(KEYINPUT94), .ZN(n634) );
  NOR2_X1 U498 ( .A1(n552), .A2(n588), .ZN(n382) );
  INV_X1 U499 ( .A(KEYINPUT60), .ZN(n402) );
  INV_X1 U500 ( .A(KEYINPUT122), .ZN(n398) );
  INV_X1 U501 ( .A(KEYINPUT56), .ZN(n423) );
  INV_X1 U502 ( .A(KEYINPUT53), .ZN(n436) );
  AND2_X1 U503 ( .A1(n637), .A2(KEYINPUT84), .ZN(n360) );
  XOR2_X1 U504 ( .A(G134), .B(G131), .Z(n361) );
  AND2_X1 U505 ( .A1(G221), .A2(n521), .ZN(n362) );
  XNOR2_X1 U506 ( .A(KEYINPUT14), .B(n503), .ZN(n363) );
  XOR2_X1 U507 ( .A(n496), .B(n495), .Z(n364) );
  OR2_X1 U508 ( .A1(n693), .A2(n692), .ZN(n365) );
  XNOR2_X1 U509 ( .A(n593), .B(KEYINPUT74), .ZN(n366) );
  XOR2_X1 U510 ( .A(KEYINPUT38), .B(n617), .Z(n680) );
  AND2_X1 U511 ( .A1(n617), .A2(n593), .ZN(n368) );
  AND2_X1 U512 ( .A1(n365), .A2(n438), .ZN(n369) );
  XNOR2_X1 U513 ( .A(KEYINPUT67), .B(KEYINPUT34), .ZN(n370) );
  XOR2_X1 U514 ( .A(n699), .B(n455), .Z(n371) );
  XNOR2_X1 U515 ( .A(n696), .B(n695), .ZN(n372) );
  XOR2_X1 U516 ( .A(n701), .B(n700), .Z(n373) );
  AND2_X1 U517 ( .A1(n624), .A2(G472), .ZN(n374) );
  INV_X1 U518 ( .A(KEYINPUT2), .ZN(n451) );
  INV_X1 U519 ( .A(n710), .ZN(n404) );
  NAND2_X1 U520 ( .A1(n675), .A2(n534), .ZN(n413) );
  NOR2_X1 U521 ( .A1(n739), .A2(n447), .ZN(n446) );
  XNOR2_X1 U522 ( .A(n453), .B(n626), .ZN(n627) );
  NAND2_X1 U523 ( .A1(n706), .A2(G210), .ZN(n425) );
  AND2_X4 U524 ( .A1(n450), .A2(n454), .ZN(n706) );
  INV_X1 U525 ( .A(n582), .ZN(n378) );
  XNOR2_X1 U526 ( .A(n437), .B(n436), .ZN(G75) );
  XNOR2_X1 U527 ( .A(n520), .B(n519), .ZN(n547) );
  XNOR2_X1 U528 ( .A(n514), .B(n513), .ZN(n515) );
  NAND2_X1 U529 ( .A1(n448), .A2(n446), .ZN(n622) );
  NAND2_X2 U530 ( .A1(n452), .A2(n451), .ZN(n450) );
  NOR2_X4 U531 ( .A1(n609), .A2(n572), .ZN(n641) );
  NAND2_X2 U532 ( .A1(n389), .A2(n570), .ZN(n609) );
  INV_X1 U533 ( .A(n585), .ZN(n567) );
  XNOR2_X2 U534 ( .A(n670), .B(KEYINPUT100), .ZN(n585) );
  INV_X1 U535 ( .A(n578), .ZN(n379) );
  XNOR2_X1 U536 ( .A(n425), .B(n372), .ZN(n386) );
  INV_X1 U537 ( .A(n715), .ZN(n380) );
  NAND2_X1 U538 ( .A1(n544), .A2(n541), .ZN(n388) );
  XNOR2_X1 U539 ( .A(n506), .B(KEYINPUT16), .ZN(n427) );
  NAND2_X1 U540 ( .A1(n729), .A2(n653), .ZN(n652) );
  XNOR2_X2 U541 ( .A(n622), .B(n621), .ZN(n729) );
  NOR2_X1 U542 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U543 ( .A1(n384), .A2(n369), .ZN(n437) );
  XNOR2_X1 U544 ( .A(n658), .B(n385), .ZN(n384) );
  NAND2_X1 U545 ( .A1(n386), .A2(n404), .ZN(n424) );
  NAND2_X1 U546 ( .A1(n422), .A2(n366), .ZN(n421) );
  NAND2_X1 U547 ( .A1(n553), .A2(n539), .ZN(n392) );
  XNOR2_X1 U548 ( .A(n485), .B(n443), .ZN(n625) );
  NAND2_X1 U549 ( .A1(n619), .A2(n606), .ZN(n445) );
  NOR2_X2 U550 ( .A1(n394), .A2(n558), .ZN(n397) );
  XNOR2_X1 U551 ( .A(n543), .B(n542), .ZN(n394) );
  XNOR2_X1 U552 ( .A(n528), .B(n527), .ZN(n530) );
  NAND2_X1 U553 ( .A1(n468), .A2(G221), .ZN(n465) );
  XNOR2_X1 U554 ( .A(n464), .B(KEYINPUT20), .ZN(n468) );
  XNOR2_X2 U555 ( .A(n397), .B(n559), .ZN(n715) );
  XNOR2_X1 U556 ( .A(n424), .B(n423), .ZN(G51) );
  XNOR2_X1 U557 ( .A(n399), .B(n398), .ZN(G54) );
  NAND2_X1 U558 ( .A1(n400), .A2(n404), .ZN(n399) );
  XNOR2_X1 U559 ( .A(n401), .B(n371), .ZN(n400) );
  NAND2_X1 U560 ( .A1(n706), .A2(G469), .ZN(n401) );
  XNOR2_X1 U561 ( .A(n403), .B(n402), .ZN(G60) );
  NAND2_X1 U562 ( .A1(n405), .A2(n404), .ZN(n403) );
  XNOR2_X1 U563 ( .A(n406), .B(n373), .ZN(n405) );
  NAND2_X1 U564 ( .A1(n706), .A2(G475), .ZN(n406) );
  XNOR2_X2 U565 ( .A(n415), .B(G469), .ZN(n570) );
  NAND2_X1 U566 ( .A1(n420), .A2(n417), .ZN(n416) );
  NAND2_X1 U567 ( .A1(n419), .A2(n418), .ZN(n417) );
  INV_X1 U568 ( .A(n637), .ZN(n418) );
  NOR2_X1 U569 ( .A1(n740), .A2(KEYINPUT84), .ZN(n419) );
  XNOR2_X1 U570 ( .A(n426), .B(n497), .ZN(n694) );
  XNOR2_X1 U571 ( .A(n427), .B(n490), .ZN(n718) );
  XNOR2_X2 U572 ( .A(n367), .B(n483), .ZN(n722) );
  XNOR2_X2 U573 ( .A(n429), .B(n428), .ZN(n534) );
  XNOR2_X2 U574 ( .A(n582), .B(KEYINPUT19), .ZN(n571) );
  AND2_X2 U575 ( .A1(n655), .A2(n624), .ZN(n454) );
  NAND2_X1 U576 ( .A1(n431), .A2(n368), .ZN(n594) );
  INV_X2 U577 ( .A(G143), .ZN(n457) );
  XOR2_X1 U578 ( .A(n698), .B(n697), .Z(n455) );
  AND2_X1 U579 ( .A1(G224), .A2(n560), .ZN(n456) );
  INV_X1 U580 ( .A(KEYINPUT65), .ZN(n603) );
  XNOR2_X1 U581 ( .A(n492), .B(n456), .ZN(n493) );
  INV_X1 U582 ( .A(KEYINPUT44), .ZN(n542) );
  XNOR2_X1 U583 ( .A(n459), .B(n484), .ZN(n460) );
  INV_X1 U584 ( .A(G475), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U586 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n559) );
  INV_X1 U587 ( .A(KEYINPUT39), .ZN(n604) );
  NOR2_X1 U588 ( .A1(G952), .A2(n560), .ZN(n710) );
  XNOR2_X2 U589 ( .A(n457), .B(G128), .ZN(n524) );
  NAND2_X1 U590 ( .A1(G227), .A2(n560), .ZN(n459) );
  XNOR2_X1 U591 ( .A(n485), .B(n462), .ZN(n699) );
  XOR2_X1 U592 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n466) );
  INV_X1 U593 ( .A(n624), .ZN(n463) );
  NAND2_X1 U594 ( .A1(G234), .A2(n463), .ZN(n464) );
  XNOR2_X1 U595 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U596 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n470) );
  NAND2_X1 U597 ( .A1(G217), .A2(n468), .ZN(n469) );
  XNOR2_X1 U598 ( .A(n470), .B(n469), .ZN(n481) );
  XOR2_X1 U599 ( .A(KEYINPUT24), .B(G110), .Z(n472) );
  XNOR2_X1 U600 ( .A(n472), .B(n471), .ZN(n476) );
  XOR2_X1 U601 ( .A(KEYINPUT89), .B(KEYINPUT71), .Z(n474) );
  XNOR2_X1 U602 ( .A(n474), .B(n473), .ZN(n475) );
  INV_X1 U603 ( .A(n492), .ZN(n477) );
  XNOR2_X1 U604 ( .A(KEYINPUT10), .B(n477), .ZN(n505) );
  XNOR2_X1 U605 ( .A(n478), .B(n505), .ZN(n727) );
  XNOR2_X1 U606 ( .A(n479), .B(n727), .ZN(n705) );
  NAND2_X1 U607 ( .A1(n532), .A2(n540), .ZN(n661) );
  NOR2_X1 U608 ( .A1(n662), .A2(n661), .ZN(n482) );
  XNOR2_X1 U609 ( .A(n482), .B(KEYINPUT68), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n507), .A2(G210), .ZN(n486) );
  XNOR2_X1 U611 ( .A(G137), .B(KEYINPUT69), .ZN(n488) );
  XNOR2_X2 U612 ( .A(n489), .B(G472), .ZN(n670) );
  XNOR2_X1 U613 ( .A(KEYINPUT6), .B(n670), .ZN(n577) );
  INV_X1 U614 ( .A(n577), .ZN(n539) );
  XOR2_X2 U615 ( .A(G122), .B(G104), .Z(n506) );
  NOR2_X1 U616 ( .A1(n624), .A2(n694), .ZN(n499) );
  NAND2_X1 U617 ( .A1(G210), .A2(n500), .ZN(n498) );
  XNOR2_X1 U618 ( .A(n499), .B(n498), .ZN(n592) );
  NAND2_X1 U619 ( .A1(G214), .A2(n500), .ZN(n679) );
  NAND2_X1 U620 ( .A1(n592), .A2(n679), .ZN(n582) );
  XOR2_X1 U621 ( .A(KEYINPUT87), .B(G898), .Z(n712) );
  NOR2_X1 U622 ( .A1(n712), .A2(n560), .ZN(n724) );
  NAND2_X1 U623 ( .A1(n724), .A2(G902), .ZN(n501) );
  NAND2_X1 U624 ( .A1(G952), .A2(n560), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n501), .A2(n562), .ZN(n502) );
  INV_X1 U626 ( .A(n534), .ZN(n551) );
  XNOR2_X1 U627 ( .A(n506), .B(n505), .ZN(n516) );
  NAND2_X1 U628 ( .A1(G214), .A2(n507), .ZN(n508) );
  XNOR2_X1 U629 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U630 ( .A(n510), .B(KEYINPUT12), .Z(n514) );
  XNOR2_X1 U631 ( .A(n512), .B(n511), .ZN(n513) );
  NOR2_X1 U632 ( .A1(G902), .A2(n701), .ZN(n520) );
  XNOR2_X1 U633 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n518) );
  NAND2_X1 U634 ( .A1(G217), .A2(n521), .ZN(n522) );
  XNOR2_X1 U635 ( .A(n523), .B(n522), .ZN(n528) );
  XNOR2_X1 U636 ( .A(n524), .B(G107), .ZN(n526) );
  XOR2_X1 U637 ( .A(G116), .B(KEYINPUT7), .Z(n529) );
  XNOR2_X1 U638 ( .A(n530), .B(n529), .ZN(n703) );
  NOR2_X1 U639 ( .A1(n703), .A2(G902), .ZN(n531) );
  NOR2_X1 U640 ( .A1(n547), .A2(n549), .ZN(n593) );
  NAND2_X1 U641 ( .A1(n547), .A2(n549), .ZN(n682) );
  NOR2_X1 U642 ( .A1(n682), .A2(n665), .ZN(n533) );
  NAND2_X1 U643 ( .A1(n534), .A2(n533), .ZN(n535) );
  INV_X1 U644 ( .A(n357), .ZN(n614) );
  NAND2_X1 U645 ( .A1(n567), .A2(n536), .ZN(n537) );
  INV_X1 U646 ( .A(n540), .ZN(n666) );
  AND2_X1 U647 ( .A1(n666), .A2(n614), .ZN(n541) );
  AND2_X1 U648 ( .A1(n357), .A2(n544), .ZN(n545) );
  XNOR2_X1 U649 ( .A(n545), .B(KEYINPUT83), .ZN(n546) );
  NOR2_X1 U650 ( .A1(n666), .A2(n546), .ZN(n629) );
  INV_X1 U651 ( .A(n547), .ZN(n548) );
  NOR2_X1 U652 ( .A1(n549), .A2(n548), .ZN(n646) );
  NOR2_X1 U653 ( .A1(n646), .A2(n606), .ZN(n684) );
  INV_X1 U654 ( .A(n661), .ZN(n550) );
  NAND2_X1 U655 ( .A1(n570), .A2(n550), .ZN(n588) );
  OR2_X1 U656 ( .A1(n670), .A2(n551), .ZN(n552) );
  NAND2_X1 U657 ( .A1(n553), .A2(n670), .ZN(n554) );
  XNOR2_X1 U658 ( .A(KEYINPUT99), .B(n557), .ZN(n558) );
  INV_X1 U659 ( .A(n684), .ZN(n595) );
  OR2_X1 U660 ( .A1(KEYINPUT77), .A2(n595), .ZN(n573) );
  NOR2_X1 U661 ( .A1(G900), .A2(n560), .ZN(n561) );
  NAND2_X1 U662 ( .A1(n561), .A2(G902), .ZN(n563) );
  NAND2_X1 U663 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U664 ( .A1(n564), .A2(n363), .ZN(n589) );
  NOR2_X1 U665 ( .A1(n589), .A2(n665), .ZN(n565) );
  XNOR2_X1 U666 ( .A(n565), .B(KEYINPUT66), .ZN(n566) );
  NAND2_X1 U667 ( .A1(n566), .A2(n666), .ZN(n578) );
  XNOR2_X1 U668 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n568) );
  INV_X1 U669 ( .A(n571), .ZN(n572) );
  NAND2_X1 U670 ( .A1(n573), .A2(n641), .ZN(n574) );
  NAND2_X1 U671 ( .A1(n574), .A2(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U672 ( .A1(n595), .A2(KEYINPUT77), .ZN(n575) );
  NAND2_X1 U673 ( .A1(n576), .A2(n575), .ZN(n602) );
  XNOR2_X1 U674 ( .A(KEYINPUT102), .B(n579), .ZN(n580) );
  NAND2_X1 U675 ( .A1(n580), .A2(n643), .ZN(n581) );
  XNOR2_X1 U676 ( .A(n583), .B(KEYINPUT36), .ZN(n584) );
  NAND2_X1 U677 ( .A1(n584), .A2(n614), .ZN(n651) );
  NAND2_X1 U678 ( .A1(n585), .A2(n679), .ZN(n587) );
  NOR2_X1 U679 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U680 ( .A1(KEYINPUT47), .A2(n597), .ZN(n598) );
  NOR2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U682 ( .A1(n651), .A2(n600), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n680), .A2(n679), .ZN(n683) );
  NOR2_X1 U684 ( .A1(n683), .A2(n682), .ZN(n608) );
  XNOR2_X1 U685 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n607) );
  NOR2_X1 U686 ( .A1(n609), .A2(n678), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n610), .B(KEYINPUT42), .ZN(n743) );
  INV_X1 U688 ( .A(KEYINPUT48), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n679), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT43), .ZN(n616) );
  NOR2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U693 ( .A(KEYINPUT104), .B(n618), .ZN(n739) );
  NAND2_X1 U694 ( .A1(n619), .A2(n646), .ZN(n620) );
  XNOR2_X1 U695 ( .A(KEYINPUT110), .B(n620), .ZN(n742) );
  INV_X1 U696 ( .A(KEYINPUT81), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n625), .B(KEYINPUT62), .ZN(n626) );
  NOR2_X1 U698 ( .A1(n710), .A2(n627), .ZN(n628) );
  XOR2_X1 U699 ( .A(KEYINPUT63), .B(n628), .Z(G57) );
  XOR2_X1 U700 ( .A(G101), .B(n629), .Z(G3) );
  NAND2_X1 U701 ( .A1(n634), .A2(n643), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n630), .B(G104), .ZN(G6) );
  XOR2_X1 U703 ( .A(KEYINPUT112), .B(KEYINPUT27), .Z(n632) );
  XNOR2_X1 U704 ( .A(G107), .B(KEYINPUT26), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(n633) );
  XOR2_X1 U706 ( .A(KEYINPUT111), .B(n633), .Z(n636) );
  NAND2_X1 U707 ( .A1(n646), .A2(n634), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(G9) );
  XOR2_X1 U709 ( .A(G110), .B(n637), .Z(G12) );
  XOR2_X1 U710 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n639) );
  NAND2_X1 U711 ( .A1(n641), .A2(n646), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(n640) );
  XOR2_X1 U713 ( .A(G128), .B(n640), .Z(G30) );
  NAND2_X1 U714 ( .A1(n641), .A2(n643), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n642), .B(G146), .ZN(G48) );
  NAND2_X1 U716 ( .A1(n645), .A2(n643), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n644), .B(G113), .ZN(G15) );
  XOR2_X1 U718 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n648) );
  NAND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U720 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U721 ( .A(G116), .B(n649), .ZN(G18) );
  XOR2_X1 U722 ( .A(G125), .B(KEYINPUT37), .Z(n650) );
  XNOR2_X1 U723 ( .A(n651), .B(n650), .ZN(G27) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(KEYINPUT76), .Z(n653) );
  XNOR2_X1 U725 ( .A(KEYINPUT79), .B(n652), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n715), .A2(n653), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U728 ( .A1(n678), .A2(n687), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n659), .B(KEYINPUT119), .ZN(n660) );
  XOR2_X1 U730 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n664) );
  NAND2_X1 U731 ( .A1(n357), .A2(n661), .ZN(n663) );
  XNOR2_X1 U732 ( .A(n664), .B(n663), .ZN(n673) );
  NAND2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(KEYINPUT116), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n668), .B(KEYINPUT49), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT117), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U740 ( .A(KEYINPUT51), .B(n676), .Z(n677) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n690) );
  NOR2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n688) );
  NOR2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U747 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U748 ( .A(KEYINPUT52), .B(n691), .ZN(n693) );
  NAND2_X1 U749 ( .A1(n363), .A2(G952), .ZN(n692) );
  XOR2_X1 U750 ( .A(KEYINPUT75), .B(KEYINPUT55), .Z(n696) );
  XNOR2_X1 U751 ( .A(n694), .B(KEYINPUT54), .ZN(n695) );
  XOR2_X1 U752 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n698) );
  XNOR2_X1 U753 ( .A(KEYINPUT121), .B(KEYINPUT120), .ZN(n697) );
  INV_X1 U754 ( .A(KEYINPUT59), .ZN(n700) );
  NAND2_X1 U755 ( .A1(G478), .A2(n706), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U757 ( .A1(n710), .A2(n704), .ZN(G63) );
  XOR2_X1 U758 ( .A(n705), .B(KEYINPUT123), .Z(n708) );
  NAND2_X1 U759 ( .A1(n706), .A2(G217), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U761 ( .A1(n710), .A2(n709), .ZN(G66) );
  NAND2_X1 U762 ( .A1(G953), .A2(G224), .ZN(n711) );
  XNOR2_X1 U763 ( .A(KEYINPUT61), .B(n711), .ZN(n713) );
  NAND2_X1 U764 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U765 ( .A(KEYINPUT124), .B(n714), .Z(n717) );
  NOR2_X1 U766 ( .A1(G953), .A2(n715), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(n726) );
  XOR2_X1 U768 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n720) );
  XNOR2_X1 U769 ( .A(G101), .B(n718), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U772 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U773 ( .A(n726), .B(n725), .Z(G69) );
  XOR2_X1 U774 ( .A(n728), .B(n727), .Z(n732) );
  XOR2_X1 U775 ( .A(n732), .B(n729), .Z(n730) );
  NOR2_X1 U776 ( .A1(G953), .A2(n730), .ZN(n731) );
  XNOR2_X1 U777 ( .A(n731), .B(KEYINPUT127), .ZN(n736) );
  XNOR2_X1 U778 ( .A(G227), .B(n732), .ZN(n733) );
  NAND2_X1 U779 ( .A1(n733), .A2(G900), .ZN(n734) );
  NAND2_X1 U780 ( .A1(n734), .A2(G953), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n736), .A2(n735), .ZN(G72) );
  XOR2_X1 U782 ( .A(n737), .B(G122), .Z(G24) );
  XOR2_X1 U783 ( .A(n358), .B(n738), .Z(G45) );
  XOR2_X1 U784 ( .A(G140), .B(n739), .Z(G42) );
  XOR2_X1 U785 ( .A(n740), .B(G119), .Z(G21) );
  XOR2_X1 U786 ( .A(n741), .B(G131), .Z(G33) );
  XNOR2_X1 U787 ( .A(G134), .B(n742), .ZN(G36) );
  XOR2_X1 U788 ( .A(n743), .B(G137), .Z(G39) );
endmodule

