//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT16), .A3(new_n203), .ZN(new_n204));
  OAI221_X1 g003(.A(new_n204), .B1(KEYINPUT92), .B2(G8gat), .C1(new_n203), .C2(new_n202), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OR3_X1    g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT88), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n214), .B1(new_n211), .B2(KEYINPUT88), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n210), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217));
  INV_X1    g016(.A(G43gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G50gat), .ZN(new_n219));
  INV_X1    g018(.A(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G43gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n217), .B1(new_n222), .B2(KEYINPUT87), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(KEYINPUT87), .B2(new_n222), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n216), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT89), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT90), .B(G43gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n220), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT15), .B1(new_n228), .B2(new_n219), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT91), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n210), .B1(new_n211), .B2(new_n213), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n207), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n226), .A2(KEYINPUT17), .A3(new_n232), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n207), .A2(KEYINPUT93), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n207), .A2(KEYINPUT93), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n233), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(KEYINPUT18), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n240), .B(new_n233), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n244), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT18), .ZN(new_n249));
  INV_X1    g048(.A(new_n244), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n242), .B2(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n245), .A2(new_n248), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT11), .ZN(new_n254));
  INV_X1    g053(.A(G169gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G197gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT86), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n252), .A2(new_n259), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n264));
  INV_X1    g063(.A(G228gat), .ZN(new_n265));
  INV_X1    g064(.A(G233gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269));
  INV_X1    g068(.A(G211gat), .ZN(new_n270));
  INV_X1    g069(.A(G218gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n268), .A3(new_n272), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT76), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT29), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n278), .B(new_n279), .C1(KEYINPUT76), .C2(new_n276), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  INV_X1    g086(.A(G162gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290));
  AOI211_X1 g089(.A(new_n283), .B(new_n285), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT79), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n285), .B2(new_n283), .ZN(new_n293));
  INV_X1    g092(.A(G141gat), .ZN(new_n294));
  INV_X1    g093(.A(G148gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(KEYINPUT79), .A3(new_n284), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n297), .A3(new_n286), .ZN(new_n298));
  XOR2_X1   g097(.A(G155gat), .B(G162gat), .Z(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT80), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT80), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n291), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n267), .B1(new_n282), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT83), .ZN(new_n306));
  INV_X1    g105(.A(new_n291), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n298), .A2(new_n302), .A3(new_n299), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n302), .B1(new_n298), .B2(new_n299), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n281), .B(new_n307), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n310), .B2(new_n279), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n278), .B1(KEYINPUT76), .B2(new_n276), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n306), .A3(new_n279), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n305), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n279), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n312), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT29), .B1(new_n276), .B2(new_n277), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(KEYINPUT3), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n267), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(G22gat), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n321), .ZN(new_n324));
  INV_X1    g123(.A(new_n267), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G22gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n315), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n328), .A2(new_n313), .A3(new_n311), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n326), .B(new_n327), .C1(new_n329), .C2(new_n305), .ZN(new_n330));
  XNOR2_X1  g129(.A(G78gat), .B(G106gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT31), .B(G50gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n323), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n323), .B2(new_n330), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT32), .ZN(new_n338));
  OR2_X1    g137(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(G127gat), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G127gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G134gat), .ZN(new_n343));
  INV_X1    g142(.A(G120gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G113gat), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT1), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n341), .A2(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n345), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT69), .B(G113gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(G120gat), .ZN(new_n354));
  INV_X1    g153(.A(G134gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G127gat), .ZN(new_n356));
  AND2_X1   g155(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n357));
  NOR2_X1   g156(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n343), .B(new_n356), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n354), .A2(KEYINPUT71), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT71), .ZN(new_n361));
  INV_X1    g160(.A(new_n359), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n346), .A2(KEYINPUT69), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G113gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n365), .A3(G120gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n345), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n361), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n351), .B1(new_n360), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT72), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT71), .B1(new_n354), .B2(new_n359), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n362), .A2(new_n367), .A3(new_n361), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n350), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT72), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT24), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT24), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(G183gat), .A3(G190gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT66), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(G183gat), .B2(G190gat), .ZN(new_n383));
  INV_X1    g182(.A(G183gat), .ZN(new_n384));
  INV_X1    g183(.A(G190gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT66), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n381), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(KEYINPUT65), .ZN(new_n389));
  NOR2_X1   g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT23), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n387), .A2(KEYINPUT25), .A3(new_n389), .A4(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(G169gat), .B2(G176gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n388), .A2(KEYINPUT65), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n393), .B(new_n391), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n378), .A2(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT67), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n390), .B(KEYINPUT26), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n389), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT27), .B(G183gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n385), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT28), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT28), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n410), .A3(new_n385), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n406), .A2(new_n409), .A3(new_n411), .A4(new_n377), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT67), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n402), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n404), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT73), .B1(new_n376), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n371), .A2(new_n372), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n374), .B1(new_n417), .B2(new_n351), .ZN(new_n418));
  AOI211_X1 g217(.A(KEYINPUT72), .B(new_n350), .C1(new_n371), .C2(new_n372), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n395), .A2(new_n402), .A3(new_n413), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n413), .B1(new_n395), .B2(new_n402), .ZN(new_n422));
  INV_X1    g221(.A(new_n412), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT73), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n420), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n376), .A2(new_n415), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n416), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n429), .B(KEYINPUT64), .Z(new_n430));
  AOI21_X1  g229(.A(new_n338), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n430), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G15gat), .B(G43gat), .Z(new_n436));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n432), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n416), .A2(new_n426), .A3(new_n429), .A4(new_n427), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT34), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n430), .A2(KEYINPUT34), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n416), .A2(new_n426), .A3(new_n427), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT74), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(KEYINPUT74), .A3(new_n443), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT33), .B1(new_n428), .B2(new_n430), .ZN(new_n448));
  INV_X1    g247(.A(new_n438), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n431), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n439), .A2(new_n446), .A3(new_n447), .A4(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT74), .B1(new_n441), .B2(new_n443), .ZN(new_n453));
  AOI221_X4 g252(.A(new_n338), .B1(KEYINPUT33), .B2(new_n438), .C1(new_n428), .C2(new_n430), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n447), .B1(new_n455), .B2(new_n439), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n264), .B(new_n337), .C1(new_n452), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n458));
  XNOR2_X1  g257(.A(G1gat), .B(G29gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT0), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G57gat), .ZN(new_n461));
  XOR2_X1   g260(.A(new_n461), .B(G85gat), .Z(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n304), .A2(new_n281), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n310), .A2(new_n369), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n304), .A2(new_n373), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT4), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT4), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n370), .A2(new_n375), .A3(new_n472), .A4(new_n304), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n463), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n467), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n319), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n465), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n470), .A2(KEYINPUT4), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n370), .A2(new_n304), .A3(new_n375), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT4), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n480), .B1(new_n482), .B2(KEYINPUT81), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n484), .A3(KEYINPUT4), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n479), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n319), .A2(new_n369), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n470), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT5), .B1(new_n488), .B2(new_n465), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n458), .B(new_n475), .C1(new_n486), .C2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n418), .A2(new_n419), .A3(new_n319), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT81), .B1(new_n493), .B2(new_n472), .ZN(new_n494));
  INV_X1    g293(.A(new_n480), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n485), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n479), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n489), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n469), .A2(new_n474), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n463), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(G226gat), .A2(G233gat), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n404), .A2(new_n412), .A3(new_n503), .A4(new_n414), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n403), .A2(new_n412), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n503), .A2(KEYINPUT29), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n313), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n403), .A2(new_n412), .A3(new_n503), .ZN(new_n510));
  INV_X1    g309(.A(new_n506), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n510), .B(new_n312), .C1(new_n424), .C2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G36gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT77), .B(G8gat), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n514), .B(new_n515), .Z(new_n516));
  NAND3_X1  g315(.A1(new_n509), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(KEYINPUT78), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n512), .ZN(new_n520));
  INV_X1    g319(.A(new_n516), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(KEYINPUT78), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT30), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n499), .A2(new_n462), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT82), .B1(new_n498), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n501), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n502), .B(new_n527), .C1(new_n530), .C2(KEYINPUT6), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT35), .B1(new_n457), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT6), .B1(new_n501), .B2(new_n529), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n499), .B1(new_n486), .B2(new_n489), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n490), .A2(new_n491), .B1(new_n534), .B2(new_n463), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n533), .A2(new_n535), .A3(new_n526), .ZN(new_n536));
  INV_X1    g335(.A(new_n444), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n431), .A2(new_n448), .A3(new_n449), .ZN(new_n538));
  OAI211_X1 g337(.A(KEYINPUT74), .B(new_n537), .C1(new_n538), .C2(new_n454), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n336), .B1(new_n539), .B2(new_n451), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n536), .A2(new_n540), .A3(new_n264), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n532), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT36), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n544), .A3(new_n451), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT75), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n539), .A2(new_n451), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT75), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n539), .A2(new_n451), .A3(new_n549), .A4(new_n544), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT38), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT84), .B(KEYINPUT37), .Z(new_n553));
  NAND3_X1  g352(.A1(new_n509), .A2(new_n512), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n554), .A2(new_n521), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n520), .A2(KEYINPUT37), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n508), .A2(new_n312), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n510), .B(new_n313), .C1(new_n424), .C2(new_n511), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(KEYINPUT37), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(new_n554), .A3(new_n552), .A4(new_n521), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n517), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n533), .B2(new_n535), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n523), .A2(new_n525), .B1(new_n534), .B2(new_n463), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n465), .B1(new_n474), .B2(new_n478), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT39), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n463), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n567), .B1(new_n488), .B2(new_n465), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n471), .A2(new_n473), .B1(new_n476), .B2(new_n477), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n570), .B2(new_n465), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT40), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT40), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n568), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n336), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n531), .A2(new_n336), .B1(new_n564), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n551), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n263), .B1(new_n543), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G64gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G57gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT95), .B(G57gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n584), .B2(new_n581), .ZN(new_n585));
  NOR2_X1   g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n581), .A2(G57gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT9), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n591), .A2(new_n582), .B1(new_n592), .B2(new_n588), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n586), .B1(KEYINPUT94), .B2(new_n588), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(KEYINPUT94), .B2(new_n588), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n590), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n240), .B1(KEYINPUT21), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G183gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n596), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G127gat), .B(G155gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G211gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n603), .A2(new_n610), .A3(new_n604), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n233), .A2(new_n234), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT98), .B(G85gat), .Z(new_n616));
  INV_X1    g415(.A(G92gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n616), .A2(new_n617), .B1(KEYINPUT8), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n620));
  NAND2_X1  g419(.A1(G85gat), .A2(G92gat), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G99gat), .B(G106gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT99), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n627), .A2(KEYINPUT100), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n624), .A2(new_n626), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(KEYINPUT100), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n236), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  AND2_X1   g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n633), .A2(new_n233), .B1(KEYINPUT41), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n634), .A2(KEYINPUT41), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT96), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G134gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n636), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G190gat), .B(G218gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G162gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n614), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(G230gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n266), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n624), .B2(KEYINPUT102), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n652), .A2(new_n626), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n626), .B2(KEYINPUT103), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n655), .A2(new_n624), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n597), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n631), .A2(KEYINPUT101), .A3(new_n596), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n631), .B2(new_n596), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n650), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n633), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n649), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n663), .A2(new_n649), .ZN(new_n664));
  XNOR2_X1  g463(.A(G120gat), .B(G148gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G176gat), .ZN(new_n666));
  INV_X1    g465(.A(G204gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OR3_X1    g468(.A1(new_n662), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n662), .B2(new_n664), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n647), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n580), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n533), .A2(new_n535), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n526), .ZN(new_n679));
  NOR2_X1   g478(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT16), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n683), .A2(G8gat), .B1(new_n684), .B2(new_n679), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(G8gat), .B2(new_n683), .ZN(G1325gat));
  AOI21_X1  g485(.A(G15gat), .B1(new_n674), .B2(new_n547), .ZN(new_n687));
  INV_X1    g486(.A(new_n551), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT105), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n687), .B1(new_n674), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n336), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT106), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT43), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(new_n327), .ZN(G1327gat));
  NOR3_X1   g494(.A1(new_n614), .A2(new_n646), .A3(new_n672), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n580), .A2(new_n208), .A3(new_n676), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT45), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n543), .A2(new_n579), .ZN(new_n700));
  INV_X1    g499(.A(new_n646), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n564), .A2(new_n577), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n536), .A2(KEYINPUT108), .A3(new_n337), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n531), .B2(new_n336), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n551), .B(new_n704), .C1(new_n705), .C2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n703), .B1(new_n708), .B2(new_n543), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n702), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n672), .B(KEYINPUT107), .Z(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR4_X1   g511(.A1(new_n710), .A2(new_n263), .A3(new_n614), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n676), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n698), .B1(new_n715), .B2(new_n208), .ZN(G1328gat));
  NAND4_X1  g515(.A1(new_n580), .A2(new_n209), .A3(new_n526), .A4(new_n696), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT46), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n713), .A2(new_n526), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n719), .B2(G36gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT109), .ZN(G1329gat));
  NAND2_X1  g520(.A1(new_n713), .A2(new_n688), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n227), .ZN(new_n723));
  INV_X1    g522(.A(new_n227), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n580), .A2(new_n724), .A3(new_n547), .A4(new_n696), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n723), .A2(new_n725), .B1(KEYINPUT110), .B2(KEYINPUT47), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1330gat));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n336), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G50gat), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n580), .A2(new_n220), .A3(new_n336), .A4(new_n696), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n729), .A3(new_n732), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n734), .A2(KEYINPUT48), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT48), .B1(new_n734), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n708), .A2(new_n543), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n711), .A2(new_n647), .A3(new_n262), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n676), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT112), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n583), .ZN(G1332gat));
  XOR2_X1   g543(.A(new_n526), .B(KEYINPUT113), .Z(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  NAND2_X1  g549(.A1(new_n741), .A2(new_n688), .ZN(new_n751));
  AOI21_X1  g550(.A(G71gat), .B1(new_n539), .B2(new_n451), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n751), .A2(G71gat), .B1(new_n741), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT114), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n741), .A2(new_n336), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  INV_X1    g556(.A(new_n614), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n263), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n646), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n739), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n739), .A2(new_n760), .A3(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n672), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n767), .A2(new_n676), .A3(new_n616), .ZN(new_n768));
  INV_X1    g567(.A(new_n672), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n759), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n702), .B2(new_n709), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT115), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n773), .B(new_n770), .C1(new_n702), .C2(new_n709), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n675), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n768), .B1(new_n616), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT116), .ZN(G1336gat));
  NAND4_X1  g577(.A1(new_n765), .A2(new_n617), .A3(new_n712), .A4(new_n746), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n771), .B2(new_n745), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n779), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n772), .A2(new_n526), .A3(new_n774), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(G92gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n785), .B2(new_n780), .ZN(G1337gat));
  INV_X1    g585(.A(G99gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n767), .A2(new_n787), .A3(new_n547), .ZN(new_n788));
  OAI21_X1  g587(.A(G99gat), .B1(new_n775), .B2(new_n551), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  INV_X1    g589(.A(G106gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n336), .A2(new_n791), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n711), .B(new_n792), .C1(new_n763), .C2(new_n764), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  OAI21_X1  g594(.A(G106gat), .B1(new_n771), .B2(new_n337), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n772), .A2(new_n336), .A3(new_n774), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G106gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n794), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT117), .B1(new_n800), .B2(KEYINPUT53), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n793), .B1(new_n798), .B2(G106gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n802), .A2(new_n803), .A3(new_n795), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n797), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(KEYINPUT118), .B(new_n797), .C1(new_n801), .C2(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1339gat));
  INV_X1    g608(.A(new_n662), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n660), .A2(new_n649), .A3(new_n661), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n668), .B1(new_n662), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT55), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n814), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n670), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n262), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT119), .B1(new_n243), .B2(new_n244), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n242), .A2(new_n822), .A3(new_n250), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n246), .A2(new_n247), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n252), .A2(new_n259), .B1(new_n825), .B2(new_n257), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n672), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n701), .B1(new_n820), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n257), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n261), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n818), .A2(new_n646), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n758), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n673), .A2(new_n263), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n675), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n540), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n746), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n353), .A3(new_n262), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n336), .B1(new_n832), .B2(new_n833), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n746), .A2(new_n675), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(new_n547), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n263), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n841), .ZN(G1340gat));
  NOR3_X1   g641(.A1(new_n840), .A2(new_n344), .A3(new_n711), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n836), .A2(new_n672), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n344), .ZN(G1341gat));
  NAND3_X1  g644(.A1(new_n836), .A2(new_n342), .A3(new_n614), .ZN(new_n846));
  OAI21_X1  g645(.A(G127gat), .B1(new_n840), .B2(new_n758), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1342gat));
  INV_X1    g647(.A(new_n835), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n646), .A2(new_n526), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n339), .A3(new_n340), .A4(new_n850), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n852));
  OAI21_X1  g651(.A(G134gat), .B1(new_n840), .B2(new_n646), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n832), .A2(new_n833), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n857), .A3(new_n336), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n839), .A2(new_n551), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n831), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n818), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n816), .A2(KEYINPUT121), .A3(new_n670), .A4(new_n817), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n262), .A3(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n830), .A2(new_n769), .A3(KEYINPUT120), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n826), .B2(new_n672), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT122), .B(new_n861), .C1(new_n870), .C2(new_n701), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n701), .B1(new_n865), .B2(new_n869), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n614), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n871), .A2(new_n874), .A3(KEYINPUT123), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n833), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT123), .B1(new_n871), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n336), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n860), .B1(new_n878), .B2(KEYINPUT57), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n294), .B1(new_n879), .B2(new_n262), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n688), .A2(new_n337), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n834), .A2(new_n881), .ZN(new_n882));
  NOR4_X1   g681(.A1(new_n882), .A2(G141gat), .A3(new_n263), .A4(new_n746), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT58), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  INV_X1    g684(.A(new_n883), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n263), .B(new_n860), .C1(new_n878), .C2(KEYINPUT57), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n294), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n884), .A2(new_n888), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n882), .A2(new_n746), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n295), .A3(new_n672), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT124), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n295), .C1(new_n879), .C2(new_n672), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n857), .B1(new_n856), .B2(new_n336), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n758), .B1(new_n872), .B2(new_n831), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n833), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n857), .A3(new_n336), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n896), .A2(new_n672), .A3(new_n859), .A4(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n894), .B1(new_n900), .B2(G148gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n892), .B1(new_n893), .B2(new_n901), .ZN(G1345gat));
  NAND3_X1  g701(.A1(new_n890), .A2(new_n287), .A3(new_n614), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n879), .A2(new_n614), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n287), .ZN(G1346gat));
  AND2_X1   g704(.A1(new_n879), .A2(new_n701), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n850), .A2(new_n288), .ZN(new_n907));
  OAI22_X1  g706(.A1(new_n906), .A2(new_n288), .B1(new_n882), .B2(new_n907), .ZN(G1347gat));
  AOI21_X1  g707(.A(new_n676), .B1(new_n832), .B2(new_n833), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n746), .A2(new_n540), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT125), .Z(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(G169gat), .B1(new_n913), .B2(new_n262), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n676), .A2(new_n527), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n838), .A2(new_n547), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n263), .A2(new_n255), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  INV_X1    g717(.A(G176gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n913), .A2(new_n919), .A3(new_n672), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n916), .A2(new_n712), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n919), .ZN(G1349gat));
  AOI21_X1  g721(.A(new_n384), .B1(new_n916), .B2(new_n614), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n614), .A2(new_n407), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n913), .B2(new_n924), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g725(.A1(new_n913), .A2(new_n385), .A3(new_n701), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n385), .B1(new_n916), .B2(new_n701), .ZN(new_n928));
  XOR2_X1   g727(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n928), .A2(new_n930), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  AND3_X1   g732(.A1(new_n909), .A2(new_n746), .A3(new_n881), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n262), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n896), .A2(new_n899), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n551), .A2(new_n915), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n262), .A2(G197gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n667), .A3(new_n672), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT62), .Z(new_n942));
  NOR3_X1   g741(.A1(new_n936), .A2(new_n711), .A3(new_n937), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n667), .B2(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n934), .A2(new_n270), .A3(new_n614), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n938), .A2(new_n614), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n946), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT63), .B1(new_n946), .B2(G211gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(G1354gat));
  AOI21_X1  g748(.A(G218gat), .B1(new_n934), .B2(new_n701), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n646), .A2(new_n271), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n938), .B2(new_n951), .ZN(G1355gat));
endmodule


