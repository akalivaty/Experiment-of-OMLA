//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1316, new_n1317, new_n1318, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406, new_n1407,
    new_n1408;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT65), .B(G50), .ZN(new_n208));
  AND3_X1   g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT66), .Z(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n212), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n206), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT67), .Z(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n214), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT68), .Z(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n223), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT69), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT70), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  AOI21_X1  g0052(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n255), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(G226), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G222), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G223), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n266), .B(new_n253), .C1(G77), .C2(new_n262), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G169), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n219), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n212), .B1(new_n206), .B2(new_n208), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n212), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI22_X1  g0078(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n272), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n272), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n221), .B1(new_n211), .B2(G20), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n283), .A2(new_n284), .B1(new_n221), .B2(new_n282), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G179), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n261), .A2(new_n287), .A3(new_n267), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n270), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n268), .A2(G200), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n280), .A2(KEYINPUT9), .A3(new_n285), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n268), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT9), .B1(new_n280), .B2(new_n285), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT10), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT72), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT72), .B(KEYINPUT10), .C1(new_n294), .C2(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n268), .A2(new_n293), .ZN(new_n301));
  AOI211_X1 g0101(.A(KEYINPUT10), .B(new_n301), .C1(KEYINPUT71), .C2(new_n291), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n291), .A2(KEYINPUT71), .ZN(new_n303));
  INV_X1    g0103(.A(new_n295), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n292), .A4(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n290), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n211), .A2(G20), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n283), .A2(G77), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G77), .B2(new_n281), .ZN(new_n309));
  INV_X1    g0109(.A(new_n274), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n310), .A2(new_n277), .B1(G20), .B2(G77), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n275), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n309), .B1(new_n272), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n256), .B1(G244), .B2(new_n260), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G232), .A2(G1698), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n264), .A2(G238), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n262), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n253), .C1(G107), .C2(new_n262), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n314), .B1(new_n269), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n315), .A2(new_n287), .A3(new_n319), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(G200), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n314), .B(new_n324), .C1(new_n293), .C2(new_n320), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT73), .B1(new_n306), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n283), .A2(G68), .A3(new_n307), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT75), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n282), .B2(new_n203), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n330), .A2(KEYINPUT12), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(KEYINPUT12), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(KEYINPUT76), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n278), .A2(new_n221), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n275), .A2(new_n207), .B1(new_n212), .B2(G68), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n272), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT11), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n237), .A2(G1698), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n262), .B(new_n341), .C1(G226), .C2(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n258), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n219), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n254), .B1(new_n345), .B2(new_n257), .ZN(new_n346));
  INV_X1    g0146(.A(new_n255), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G238), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n259), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  OR3_X1    g0154(.A1(new_n344), .A2(new_n350), .A3(new_n353), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT14), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n357), .A3(G169), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n351), .A2(KEYINPUT13), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(G179), .A3(new_n355), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n357), .B1(new_n356), .B2(G169), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n340), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n340), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n356), .A2(G200), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(G190), .A3(new_n355), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n327), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n348), .B1(new_n237), .B2(new_n259), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G33), .ZN(new_n372));
  INV_X1    g0172(.A(G87), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT77), .B1(new_n372), .B2(KEYINPUT3), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT77), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT3), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(G33), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n372), .A2(KEYINPUT3), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n264), .A2(G223), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n375), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n379), .A2(new_n380), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  AND2_X1   g0185(.A1(G226), .A2(G1698), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n376), .A4(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n376), .A2(new_n379), .A3(new_n380), .A4(new_n386), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT79), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n383), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(G179), .B(new_n371), .C1(new_n390), .C2(new_n258), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n392));
  INV_X1    g0192(.A(new_n382), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n374), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n388), .A2(KEYINPUT79), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n388), .A2(KEYINPUT79), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n370), .B1(new_n397), .B2(new_n253), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n391), .B1(new_n398), .B2(new_n269), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n262), .B2(G20), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n378), .A2(G33), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n380), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n203), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n202), .A2(new_n203), .ZN(new_n408));
  OAI21_X1  g0208(.A(G20), .B1(new_n206), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n277), .A2(G159), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n401), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n272), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n381), .A2(new_n402), .A3(new_n212), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G68), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n402), .B1(new_n381), .B2(new_n212), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT78), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT7), .B1(new_n392), .B2(G20), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT78), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n419), .A3(G68), .A4(new_n414), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n411), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n413), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  INV_X1    g0222(.A(new_n283), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n310), .A2(new_n307), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n423), .A2(new_n424), .B1(new_n281), .B2(new_n310), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n399), .B(new_n400), .C1(new_n422), .C2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n425), .ZN(new_n428));
  AOI211_X1 g0228(.A(new_n401), .B(new_n411), .C1(new_n417), .C2(new_n420), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(new_n413), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n400), .B1(new_n430), .B2(new_n399), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT80), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n293), .B(new_n371), .C1(new_n390), .C2(new_n258), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n398), .B2(G200), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n428), .C1(new_n429), .C2(new_n413), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT81), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n417), .A2(new_n420), .ZN(new_n438));
  INV_X1    g0238(.A(new_n411), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(KEYINPUT16), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n413), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n425), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n437), .B1(new_n442), .B2(new_n434), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT17), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT17), .B1(new_n442), .B2(new_n434), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n399), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT18), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT80), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n426), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n432), .A2(new_n444), .A3(new_n446), .A4(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n326), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n369), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(G257), .A2(G1698), .ZN(new_n456));
  INV_X1    g0256(.A(G264), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(G1698), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(new_n376), .A3(new_n380), .A4(new_n379), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n405), .A2(G303), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n258), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT5), .B(G41), .ZN(new_n462));
  INV_X1    g0262(.A(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(G270), .A3(new_n258), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n211), .A2(G45), .ZN(new_n467));
  OR2_X1    g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n346), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT83), .B1(new_n461), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  INV_X1    g0274(.A(G97), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n474), .B(new_n212), .C1(G33), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G20), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n272), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT20), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n476), .A2(KEYINPUT20), .A3(new_n272), .A4(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n281), .A2(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n211), .A2(G33), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n281), .A2(new_n485), .A3(new_n219), .A4(new_n271), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(new_n487), .B2(G116), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n269), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n457), .A2(G1698), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(G257), .B2(G1698), .ZN(new_n491));
  INV_X1    g0291(.A(G303), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n381), .A2(new_n491), .B1(new_n492), .B2(new_n262), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n253), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n462), .A2(new_n464), .B1(new_n345), .B2(new_n257), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(G270), .B1(new_n346), .B2(new_n470), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT83), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n473), .A2(new_n489), .A3(new_n498), .A4(KEYINPUT21), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n483), .A2(new_n488), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(G179), .A3(new_n494), .A4(new_n496), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT84), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n473), .A2(new_n498), .A3(new_n489), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT84), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n499), .A2(new_n507), .A3(new_n501), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n503), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n473), .A2(new_n498), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n500), .B1(new_n510), .B2(G190), .ZN(new_n511));
  INV_X1    g0311(.A(G200), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n495), .A2(G257), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n471), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n405), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n517), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n262), .A2(new_n519), .A3(KEYINPUT82), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n264), .A2(G244), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n381), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(G250), .A2(G1698), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n404), .A2(new_n380), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n474), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n521), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n515), .B1(new_n529), .B2(new_n253), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n287), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n527), .B1(new_n518), .B2(new_n520), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n258), .B1(new_n532), .B2(new_n524), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n269), .B1(new_n533), .B2(new_n515), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT6), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n535), .A2(new_n475), .A3(G107), .ZN(new_n536));
  XNOR2_X1  g0336(.A(G97), .B(G107), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI22_X1  g0338(.A1(new_n538), .A2(new_n212), .B1(new_n207), .B2(new_n278), .ZN(new_n539));
  INV_X1    g0339(.A(G107), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n403), .B2(new_n406), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n272), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n282), .A2(new_n475), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n487), .A2(G97), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n531), .A2(new_n534), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n212), .A2(G87), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT22), .B1(new_n262), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT23), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n212), .B2(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n540), .A2(KEYINPUT23), .A3(G20), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT22), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n373), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n392), .A2(new_n212), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n547), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n558), .B1(new_n405), .B2(new_n548), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G116), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(G20), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n552), .B2(new_n553), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n376), .A2(new_n379), .A3(new_n212), .A4(new_n380), .ZN(new_n567));
  INV_X1    g0367(.A(new_n559), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n566), .A2(new_n569), .A3(KEYINPUT24), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n272), .B1(new_n561), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n282), .A2(KEYINPUT25), .A3(new_n540), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT25), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n281), .B2(G107), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n487), .A2(G107), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G294), .ZN(new_n576));
  OR2_X1    g0376(.A1(G250), .A2(G1698), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G257), .B2(new_n264), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n381), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(new_n253), .B1(G264), .B2(new_n495), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(G190), .A3(new_n471), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n253), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n495), .A2(G264), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n471), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n571), .A2(new_n575), .A3(new_n581), .A4(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(G200), .B1(new_n533), .B2(new_n515), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n529), .A2(new_n253), .ZN(new_n588));
  INV_X1    g0388(.A(new_n515), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(G190), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n544), .A2(new_n543), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n278), .A2(new_n207), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n475), .A2(new_n540), .ZN(new_n593));
  NOR2_X1   g0393(.A1(G97), .A2(G107), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n535), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n536), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n592), .B1(new_n597), .B2(G20), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n262), .A2(new_n402), .A3(G20), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT7), .B1(new_n405), .B2(new_n212), .ZN(new_n600));
  OAI21_X1  g0400(.A(G107), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n591), .B1(new_n602), .B2(new_n272), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n587), .A2(new_n590), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n546), .A2(new_n586), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n571), .A2(new_n575), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n287), .A2(new_n582), .A3(new_n471), .A4(new_n583), .ZN(new_n607));
  AOI21_X1  g0407(.A(G169), .B1(new_n580), .B2(new_n471), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n312), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(new_n281), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT19), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n373), .A2(new_n475), .A3(new_n540), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n343), .A2(new_n212), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n613), .A2(new_n212), .A3(G33), .A4(G97), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n203), .A2(new_n567), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n618), .B2(new_n272), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n487), .A2(new_n611), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n258), .A2(G274), .A3(new_n464), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n258), .A2(G250), .A3(new_n467), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n349), .A2(new_n264), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G244), .B2(new_n264), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n563), .B1(new_n381), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n626), .B2(new_n253), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n619), .A2(new_n620), .B1(new_n287), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(G169), .B2(new_n627), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n567), .A2(new_n203), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n614), .A2(new_n615), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n617), .B1(new_n631), .B2(KEYINPUT19), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n272), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n612), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n487), .A2(G87), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n626), .A2(new_n253), .ZN(new_n637));
  INV_X1    g0437(.A(new_n623), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G190), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n636), .B(new_n639), .C1(new_n512), .C2(new_n627), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n629), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n605), .A2(new_n610), .A3(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n455), .A2(new_n509), .A3(new_n513), .A4(new_n642), .ZN(G372));
  NAND2_X1  g0443(.A1(new_n300), .A2(new_n305), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n442), .A2(new_n437), .A3(new_n434), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n445), .B1(new_n647), .B2(KEYINPUT17), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n323), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n367), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n649), .B1(new_n363), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n448), .A2(KEYINPUT87), .A3(new_n426), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT87), .B1(new_n448), .B2(new_n426), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n644), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n289), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n633), .A2(new_n634), .A3(new_n620), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n627), .A2(new_n287), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n626), .A2(KEYINPUT85), .A3(new_n253), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT85), .B1(new_n626), .B2(new_n253), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n638), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n662), .B1(new_n269), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n639), .A2(new_n619), .A3(new_n635), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(G200), .B2(new_n666), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT86), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT85), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n637), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n623), .B1(new_n672), .B2(new_n663), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n639), .B(new_n636), .C1(new_n673), .C2(new_n512), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n628), .B1(new_n673), .B2(G169), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT86), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n546), .B1(new_n670), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n605), .B1(new_n670), .B2(new_n677), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n506), .A2(new_n499), .A3(new_n501), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n610), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n588), .A2(new_n589), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n603), .B1(new_n269), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n531), .A3(new_n629), .A4(new_n640), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n667), .B1(new_n687), .B2(KEYINPUT26), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n680), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n659), .B1(new_n454), .B2(new_n690), .ZN(G369));
  NAND3_X1  g0491(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n500), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n682), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n509), .A2(new_n513), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g0501(.A(KEYINPUT88), .B(G330), .Z(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n606), .A2(new_n697), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n610), .B1(new_n586), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n697), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n610), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n509), .A2(new_n697), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n708), .A3(new_n713), .ZN(G399));
  INV_X1    g0514(.A(G41), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n215), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n614), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n222), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(new_n716), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n675), .B1(new_n687), .B2(KEYINPUT26), .ZN(new_n723));
  INV_X1    g0523(.A(new_n546), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n676), .B1(new_n674), .B2(new_n675), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n723), .B1(new_n727), .B2(KEYINPUT26), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n606), .A2(new_n609), .B1(new_n505), .B2(new_n504), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n503), .A3(new_n508), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT93), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT93), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n729), .A2(new_n503), .A3(new_n732), .A4(new_n508), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n681), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n722), .B1(new_n735), .B2(new_n707), .ZN(new_n736));
  AOI211_X1 g0536(.A(KEYINPUT94), .B(new_n697), .C1(new_n728), .C2(new_n734), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT95), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT95), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n741), .B(KEYINPUT29), .C1(new_n736), .C2(new_n737), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n689), .A2(new_n707), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n740), .A2(new_n742), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n642), .A2(new_n509), .A3(new_n513), .A4(new_n707), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n287), .B(new_n584), .C1(new_n533), .C2(new_n515), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(new_n510), .A3(new_n673), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n494), .A2(new_n496), .A3(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT89), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n580), .A2(new_n627), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT89), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n494), .A2(new_n496), .A3(new_n752), .A4(G179), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n530), .A2(KEYINPUT30), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT91), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n580), .A2(new_n627), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(KEYINPUT89), .B2(new_n749), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT91), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT30), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n533), .A2(new_n760), .A3(new_n515), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n758), .A2(new_n759), .A3(new_n753), .A4(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n748), .B1(new_n756), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT90), .B1(new_n754), .B2(new_n685), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT90), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n758), .A2(new_n765), .A3(new_n530), .A4(new_n753), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n764), .A2(new_n766), .A3(new_n760), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n746), .B1(new_n768), .B2(new_n697), .ZN(new_n769));
  AOI211_X1 g0569(.A(KEYINPUT31), .B(new_n707), .C1(new_n763), .C2(new_n767), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n745), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n702), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT92), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT92), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n771), .A2(new_n774), .A3(new_n702), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n744), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n721), .B1(new_n777), .B2(G1), .ZN(G364));
  INV_X1    g0578(.A(new_n716), .ZN(new_n779));
  INV_X1    g0579(.A(G13), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n211), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n704), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n702), .B2(new_n701), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n215), .A2(new_n262), .ZN(new_n787));
  INV_X1    g0587(.A(G355), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n788), .B1(G116), .B2(new_n215), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n251), .A2(G45), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n215), .A2(new_n381), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n463), .B2(new_n222), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n219), .B1(G20), .B2(new_n269), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n784), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n212), .A2(new_n287), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n802), .A2(new_n512), .A3(G190), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n802), .A2(new_n293), .A3(new_n512), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n804), .A2(new_n203), .B1(new_n806), .B2(new_n221), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G190), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n807), .B1(G77), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n212), .A2(G179), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(new_n293), .A3(G200), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT96), .Z(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G107), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n812), .A2(G190), .A3(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n373), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n812), .A2(new_n808), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT32), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n819), .A2(new_n820), .A3(G159), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n293), .A2(G179), .A3(G200), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n212), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n817), .B(new_n821), .C1(G97), .C2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n820), .B1(new_n819), .B2(G159), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n802), .A2(new_n293), .A3(G200), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n405), .B(new_n826), .C1(G58), .C2(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n811), .A2(new_n815), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  INV_X1    g0630(.A(G294), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n405), .B1(new_n809), .B2(new_n830), .C1(new_n823), .C2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n816), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G303), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT33), .B(G317), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G326), .A2(new_n805), .B1(new_n803), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n827), .A2(G322), .B1(G329), .B2(new_n819), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n814), .ZN(new_n839));
  INV_X1    g0639(.A(G283), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n829), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n800), .B1(new_n842), .B2(new_n797), .ZN(new_n843));
  INV_X1    g0643(.A(new_n796), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n701), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n786), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G396));
  NAND2_X1  g0647(.A1(new_n650), .A2(new_n707), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n325), .B1(new_n314), .B2(new_n707), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n323), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n743), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n851), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n689), .A2(new_n707), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n776), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n784), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n776), .A2(new_n852), .A3(new_n854), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n814), .A2(G87), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n830), .B2(new_n818), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT98), .Z(new_n861));
  AOI22_X1  g0661(.A1(new_n803), .A2(G283), .B1(G116), .B2(new_n810), .ZN(new_n862));
  INV_X1    g0662(.A(new_n827), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n831), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n262), .B1(new_n805), .B2(G303), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n865), .B1(new_n475), .B2(new_n823), .C1(new_n540), .C2(new_n816), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n861), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n839), .A2(new_n203), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n381), .B1(new_n819), .B2(G132), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n824), .A2(G58), .B1(new_n833), .B2(G50), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n803), .A2(G150), .B1(G159), .B2(new_n810), .ZN(new_n871));
  INV_X1    g0671(.A(G137), .ZN(new_n872));
  INV_X1    g0672(.A(G143), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n871), .B1(new_n872), .B2(new_n806), .C1(new_n873), .C2(new_n863), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT34), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n869), .B(new_n870), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n868), .B(new_n876), .C1(new_n875), .C2(new_n874), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n797), .B1(new_n867), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n784), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n797), .A2(new_n794), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT97), .Z(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n879), .B1(new_n882), .B2(new_n207), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n878), .B(new_n883), .C1(new_n853), .C2(new_n795), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n858), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(G384));
  NOR2_X1   g0686(.A1(new_n781), .A2(new_n211), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n743), .A2(new_n739), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n888), .A2(new_n452), .A3(new_n369), .A4(new_n453), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n740), .B2(new_n742), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n658), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT101), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n421), .A2(KEYINPUT16), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n440), .A3(new_n272), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n896), .A2(new_n428), .B1(new_n447), .B2(new_n695), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT37), .B1(new_n647), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT37), .B1(new_n430), .B2(new_n399), .ZN(new_n899));
  INV_X1    g0699(.A(new_n695), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n430), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n899), .A2(new_n645), .A3(new_n646), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n695), .B1(new_n896), .B2(new_n428), .ZN(new_n903));
  AOI221_X4 g0703(.A(new_n894), .B1(new_n898), .B2(new_n902), .C1(new_n451), .C2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT87), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n427), .B2(new_n431), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n448), .A2(KEYINPUT87), .A3(new_n426), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n906), .A2(new_n444), .A3(new_n446), .A4(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n901), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n901), .B(new_n435), .C1(new_n442), .C2(new_n447), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n902), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n893), .B1(new_n904), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n363), .A2(new_n697), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT100), .ZN(new_n917));
  INV_X1    g0717(.A(new_n903), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n448), .A2(new_n449), .A3(new_n426), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n449), .B1(new_n448), .B2(new_n426), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n918), .B1(new_n921), .B2(new_n648), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n898), .A2(new_n902), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n894), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n451), .A2(new_n903), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n898), .A2(new_n902), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(KEYINPUT38), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n915), .A2(new_n917), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n924), .A2(new_n927), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n340), .A2(new_n697), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n363), .A2(new_n367), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n363), .B2(new_n367), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n854), .B2(new_n848), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n930), .A2(new_n936), .B1(new_n656), .B2(new_n695), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n929), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n892), .B(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n934), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n851), .B1(new_n941), .B2(new_n932), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n942), .A2(new_n771), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT38), .B1(new_n925), .B2(new_n926), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n904), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n942), .A2(KEYINPUT40), .A3(new_n771), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n904), .B2(new_n914), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n455), .A2(new_n771), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n702), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n887), .B1(new_n940), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n940), .B2(new_n954), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n719), .A2(new_n207), .A3(new_n408), .ZN(new_n957));
  INV_X1    g0757(.A(new_n208), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n203), .ZN(new_n959));
  OAI211_X1 g0759(.A(G1), .B(new_n780), .C1(new_n957), .C2(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n597), .A2(KEYINPUT35), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n597), .A2(KEYINPUT35), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n961), .A2(G116), .A3(new_n220), .A4(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n956), .A2(new_n960), .A3(new_n965), .ZN(G367));
  NOR2_X1   g0766(.A1(new_n823), .A2(new_n203), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n405), .B(new_n967), .C1(G159), .C2(new_n803), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n827), .A2(G150), .B1(new_n805), .B2(G143), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n958), .A2(new_n810), .B1(new_n819), .B2(G137), .ZN(new_n970));
  INV_X1    g0770(.A(new_n813), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n833), .A2(G58), .B1(new_n971), .B2(G77), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n863), .A2(new_n492), .B1(new_n806), .B2(new_n830), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT107), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n381), .B1(new_n813), .B2(new_n475), .C1(new_n823), .C2(new_n540), .ZN(new_n977));
  XNOR2_X1  g0777(.A(KEYINPUT108), .B(G317), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G283), .A2(new_n810), .B1(new_n819), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n831), .B2(new_n804), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n976), .A2(new_n977), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n833), .A2(KEYINPUT46), .A3(G116), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT46), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n816), .B2(new_n477), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(new_n974), .C2(new_n975), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n973), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n797), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n798), .B1(new_n215), .B2(new_n312), .C1(new_n243), .C2(new_n791), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n784), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n725), .A2(new_n726), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n636), .A2(new_n707), .ZN(new_n993));
  MUX2_X1   g0793(.A(new_n992), .B(new_n675), .S(new_n993), .Z(new_n994));
  AND2_X1   g0794(.A1(new_n994), .A2(new_n796), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n546), .A2(new_n604), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n545), .A2(new_n697), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n998), .A2(new_n999), .B1(new_n724), .B2(new_n697), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT102), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(KEYINPUT102), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n610), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n697), .B1(new_n1005), .B2(new_n546), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1003), .A2(new_n713), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1006), .B1(KEYINPUT42), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(KEYINPUT42), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT43), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n994), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n994), .A2(new_n1011), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n994), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n711), .A2(new_n1003), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT103), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1020), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n713), .A2(new_n708), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n1003), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT44), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT105), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT104), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(KEYINPUT105), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1026), .A2(new_n1003), .A3(KEYINPUT104), .A4(KEYINPUT44), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1026), .A2(new_n1003), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT45), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n711), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(KEYINPUT106), .A3(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n710), .B(new_n712), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(new_n703), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1039), .A2(KEYINPUT106), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1035), .A2(new_n1037), .A3(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1040), .A2(new_n777), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n777), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n716), .B(KEYINPUT41), .Z(new_n1048));
  AOI21_X1  g0848(.A(new_n783), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n997), .B1(new_n1025), .B2(new_n1049), .ZN(G387));
  NAND2_X1  g0850(.A1(new_n777), .A2(new_n1043), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1042), .B1(new_n744), .B2(new_n776), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n779), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1042), .A2(new_n782), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT109), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n796), .B1(new_n706), .B2(new_n709), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n787), .A2(new_n717), .B1(G107), .B2(new_n215), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT110), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n240), .A2(new_n463), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n717), .ZN(new_n1060));
  AOI211_X1 g0860(.A(G45), .B(new_n1060), .C1(G68), .C2(G77), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n274), .A2(G50), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n791), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1058), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n784), .B1(new_n1065), .B2(new_n799), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n979), .A2(new_n827), .B1(new_n803), .B2(G311), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(KEYINPUT111), .B(G322), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1067), .B1(new_n492), .B2(new_n809), .C1(new_n806), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n824), .A2(G283), .B1(new_n833), .B2(G294), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n392), .B1(G326), .B2(new_n819), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n477), .B2(new_n813), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT112), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1076), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n839), .A2(new_n475), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n310), .A2(new_n803), .B1(new_n805), .B2(G159), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n221), .B2(new_n863), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G68), .A2(new_n810), .B1(new_n819), .B2(G150), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n823), .A2(new_n312), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G77), .B2(new_n833), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n392), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1081), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1066), .B1(new_n1090), .B2(new_n797), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT113), .Z(new_n1092));
  AOI21_X1  g0892(.A(new_n1055), .B1(new_n1056), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1053), .A2(new_n1093), .ZN(G393));
  XNOR2_X1  g0894(.A(new_n1038), .B(new_n711), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n783), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n248), .A2(new_n791), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n798), .B1(new_n475), .B2(new_n215), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n784), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n827), .A2(G159), .B1(new_n805), .B2(G150), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT51), .Z(new_n1101));
  OAI22_X1  g0901(.A1(new_n804), .A2(new_n208), .B1(new_n818), .B2(new_n873), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n310), .B2(new_n810), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n823), .A2(new_n207), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n381), .B(new_n1104), .C1(G68), .C2(new_n833), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n859), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n804), .A2(new_n492), .B1(new_n818), .B2(new_n1068), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n262), .B(new_n1107), .C1(G294), .C2(new_n810), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n824), .A2(G116), .B1(new_n833), .B2(G283), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n815), .A3(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n827), .A2(G311), .B1(new_n805), .B2(G317), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT52), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1106), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1099), .B1(new_n1113), .B2(new_n797), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1004), .B2(new_n844), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1095), .B1(new_n777), .B2(new_n1043), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1046), .A2(new_n779), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1096), .B(new_n1115), .C1(new_n1116), .C2(new_n1117), .ZN(G390));
  AND3_X1   g0918(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n901), .B1(new_n655), .B2(new_n648), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n913), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n894), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT39), .B1(new_n1122), .B2(new_n927), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n794), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n784), .B1(new_n881), .B2(new_n310), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT117), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n868), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G107), .A2(new_n803), .B1(new_n827), .B2(G116), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n805), .A2(G283), .B1(G294), .B2(new_n819), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n405), .B1(new_n809), .B2(new_n475), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1104), .A2(new_n1130), .A3(new_n817), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n816), .A2(new_n276), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT53), .Z(new_n1134));
  OAI21_X1  g0934(.A(new_n262), .B1(new_n804), .B2(new_n872), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G159), .B2(new_n824), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n827), .A2(G132), .B1(new_n805), .B2(G128), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n810), .A2(new_n1139), .B1(new_n819), .B2(G125), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n971), .A2(new_n958), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1136), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1132), .B1(new_n1134), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1126), .B1(new_n1144), .B2(new_n797), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1124), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n942), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n771), .A2(G330), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n917), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n904), .B2(new_n914), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n850), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n738), .B2(new_n848), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n941), .A2(KEYINPUT114), .A3(new_n932), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT114), .B1(new_n941), .B2(new_n932), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1151), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n936), .A2(new_n917), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n915), .B2(new_n928), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1149), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n771), .A2(new_n774), .A3(new_n702), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n774), .B1(new_n771), .B2(new_n702), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n942), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT115), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT115), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1165), .B(new_n942), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n936), .A2(new_n917), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n731), .A2(new_n681), .A3(new_n733), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n641), .A2(new_n546), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n667), .B1(new_n1171), .B2(new_n679), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n678), .B2(new_n679), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n707), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT94), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n735), .A2(new_n722), .A3(new_n707), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n848), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n850), .A3(new_n1156), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1122), .A2(new_n927), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n1150), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1167), .A2(new_n1169), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1160), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1146), .B1(new_n1182), .B2(new_n782), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1156), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n771), .A2(G330), .A3(new_n853), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1185), .A2(new_n1186), .B1(new_n1177), .B2(new_n850), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1165), .B1(new_n776), .B2(new_n942), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1166), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n854), .A2(new_n848), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n941), .A2(new_n932), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n776), .B2(new_n853), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1191), .B1(new_n1193), .B2(new_n1149), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n454), .A2(new_n1148), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n890), .A2(new_n658), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(new_n1182), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n716), .B1(new_n1198), .B2(new_n1182), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1199), .A2(KEYINPUT116), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT116), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1184), .B1(new_n1201), .B2(new_n1202), .ZN(G378));
  INV_X1    g1003(.A(KEYINPUT121), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n851), .B1(new_n773), .B2(new_n775), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1205), .A2(new_n1192), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1167), .A2(new_n1187), .B1(new_n1206), .B2(new_n1191), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1197), .B1(new_n1182), .B2(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n929), .A2(new_n937), .ZN(new_n1209));
  INV_X1    g1009(.A(G330), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1179), .B2(new_n948), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n286), .A2(new_n900), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n306), .B(new_n1212), .Z(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1213), .B(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n947), .A2(new_n1211), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n947), .B2(new_n1211), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1209), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT119), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1216), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n949), .A2(G330), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT40), .B1(new_n930), .B2(new_n943), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n947), .A2(new_n1211), .A3(new_n1216), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(new_n938), .A3(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1219), .A2(new_n1220), .A3(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(KEYINPUT119), .B(new_n1209), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1208), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT120), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1230), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1231), .B1(new_n1219), .B2(new_n1226), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n716), .B1(new_n1234), .B2(new_n1208), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1232), .A2(new_n1233), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1227), .A2(new_n783), .A3(new_n1228), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n863), .A2(new_n540), .B1(new_n806), .B2(new_n477), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n611), .A2(new_n810), .B1(new_n819), .B2(G283), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n475), .B2(new_n804), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n813), .A2(new_n202), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1239), .A2(new_n1241), .A3(new_n967), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n381), .A2(new_n715), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G77), .B2(new_n833), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT118), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1243), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT58), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1244), .B(new_n221), .C1(G33), .C2(G41), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n803), .A2(G132), .B1(new_n805), .B2(G125), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n827), .A2(G128), .B1(G137), .B2(new_n810), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n824), .A2(G150), .B1(new_n833), .B2(new_n1139), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(KEYINPUT59), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(KEYINPUT59), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n971), .A2(G159), .ZN(new_n1259));
  AOI211_X1 g1059(.A(G33), .B(G41), .C1(new_n819), .C2(G124), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1251), .B(new_n1252), .C1(new_n1257), .C2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n797), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n879), .B1(new_n208), .B2(new_n880), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n1221), .C2(new_n795), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1238), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1204), .B1(new_n1237), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT120), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n1271), .A3(new_n1235), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1267), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(KEYINPUT121), .A3(new_n1273), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1268), .A2(new_n1274), .ZN(G375));
  AOI211_X1 g1075(.A(new_n262), .B(new_n1087), .C1(G303), .C2(new_n819), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n475), .B2(new_n816), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n839), .A2(new_n207), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n804), .A2(new_n477), .B1(new_n809), .B2(new_n540), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n863), .A2(new_n840), .B1(new_n806), .B2(new_n831), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1139), .A2(new_n803), .B1(new_n805), .B2(G132), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n276), .B2(new_n809), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1242), .B1(G159), .B2(new_n833), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n221), .B2(new_n823), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n819), .A2(G128), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n863), .B2(new_n872), .ZN(new_n1287));
  NOR4_X1   g1087(.A1(new_n1283), .A2(new_n1285), .A3(new_n381), .A4(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n797), .B1(new_n1281), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n879), .B1(new_n882), .B2(new_n203), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1289), .B(new_n1290), .C1(new_n1156), .C2(new_n795), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1207), .B2(new_n782), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n889), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n741), .B1(new_n1295), .B2(KEYINPUT29), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n742), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1196), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n659), .A3(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1194), .A3(new_n1190), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1198), .A2(new_n1048), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1293), .A2(new_n1302), .ZN(new_n1303));
  XOR2_X1   g1103(.A(new_n1303), .B(KEYINPUT122), .Z(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(G381));
  INV_X1    g1105(.A(new_n1049), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n996), .B1(new_n1306), .B2(new_n1024), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(G390), .A2(G384), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(G393), .A2(G396), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1304), .A2(new_n1307), .A3(new_n1308), .A4(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT123), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1183), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1314));
  OR3_X1    g1114(.A1(G375), .A2(new_n1312), .A3(new_n1314), .ZN(G407));
  NAND2_X1  g1115(.A1(new_n696), .A2(G213), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1313), .A2(new_n1317), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G407), .B(G213), .C1(G375), .C2(new_n1318), .ZN(G409));
  NAND3_X1  g1119(.A1(new_n1272), .A2(G378), .A3(new_n1273), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1208), .A2(new_n1227), .A3(new_n1048), .A4(new_n1228), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1266), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1322), .B1(new_n1323), .B2(new_n783), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(KEYINPUT124), .A3(new_n1313), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT124), .B1(new_n1325), .B2(new_n1313), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1320), .A2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n779), .B1(new_n1207), .B2(new_n1300), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT60), .ZN(new_n1333));
  AOI211_X1 g1133(.A(KEYINPUT125), .B(new_n1333), .C1(new_n1207), .C2(new_n1300), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT125), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT60), .B1(new_n1301), .B2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1332), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(KEYINPUT126), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1335), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1333), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1301), .A2(new_n1335), .A3(KEYINPUT60), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT126), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(new_n1343), .A3(new_n1332), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1338), .A2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(G384), .B1(new_n1345), .B2(new_n1293), .ZN(new_n1346));
  AOI211_X1 g1146(.A(new_n885), .B(new_n1292), .C1(new_n1338), .C2(new_n1344), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1330), .A2(new_n1348), .A3(new_n1316), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(KEYINPUT62), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1343), .B1(new_n1342), .B2(new_n1332), .ZN(new_n1351));
  AOI211_X1 g1151(.A(KEYINPUT126), .B(new_n1331), .C1(new_n1340), .C2(new_n1341), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1293), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n885), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1345), .A2(G384), .A3(new_n1293), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1317), .A2(G2897), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1354), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  OAI211_X1 g1157(.A(G2897), .B(new_n1317), .C1(new_n1346), .C2(new_n1347), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1325), .A2(new_n1313), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT124), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1326), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1267), .B1(new_n1363), .B2(new_n1271), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1362), .B1(G378), .B2(new_n1364), .ZN(new_n1365));
  OAI211_X1 g1165(.A(new_n1357), .B(new_n1358), .C1(new_n1365), .C2(new_n1317), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT61), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1317), .B1(new_n1320), .B2(new_n1329), .ZN(new_n1368));
  INV_X1    g1168(.A(KEYINPUT62), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1368), .A2(new_n1369), .A3(new_n1348), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1350), .A2(new_n1366), .A3(new_n1367), .A4(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1307), .A2(G390), .ZN(new_n1372));
  INV_X1    g1172(.A(G390), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(G387), .A2(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n846), .B1(new_n1053), .B2(new_n1093), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1309), .A2(new_n1375), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1372), .A2(new_n1374), .A3(new_n1376), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1376), .B1(new_n1372), .B2(new_n1374), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1379), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1371), .A2(new_n1380), .ZN(new_n1381));
  AND3_X1   g1181(.A1(new_n1354), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1356), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1383));
  NOR2_X1   g1183(.A1(new_n1382), .A2(new_n1383), .ZN(new_n1384));
  INV_X1    g1184(.A(new_n1368), .ZN(new_n1385));
  AOI21_X1  g1185(.A(KEYINPUT61), .B1(new_n1384), .B2(new_n1385), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT63), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1349), .A2(new_n1387), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1368), .A2(KEYINPUT63), .A3(new_n1348), .ZN(new_n1389));
  NAND4_X1  g1189(.A1(new_n1386), .A2(new_n1379), .A3(new_n1388), .A4(new_n1389), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1381), .A2(new_n1390), .ZN(G405));
  INV_X1    g1191(.A(KEYINPUT127), .ZN(new_n1392));
  OAI21_X1  g1192(.A(new_n1392), .B1(new_n1377), .B2(new_n1378), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1372), .A2(new_n1374), .ZN(new_n1394));
  INV_X1    g1194(.A(new_n1376), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1394), .A2(new_n1395), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1372), .A2(new_n1374), .A3(new_n1376), .ZN(new_n1397));
  NAND3_X1  g1197(.A1(new_n1396), .A2(KEYINPUT127), .A3(new_n1397), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1393), .A2(new_n1398), .ZN(new_n1399));
  NAND3_X1  g1199(.A1(new_n1268), .A2(new_n1274), .A3(new_n1313), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1400), .A2(new_n1320), .ZN(new_n1401));
  NAND2_X1  g1201(.A1(new_n1401), .A2(new_n1348), .ZN(new_n1402));
  INV_X1    g1202(.A(new_n1348), .ZN(new_n1403));
  NAND3_X1  g1203(.A1(new_n1400), .A2(new_n1403), .A3(new_n1320), .ZN(new_n1404));
  NAND3_X1  g1204(.A1(new_n1399), .A2(new_n1402), .A3(new_n1404), .ZN(new_n1405));
  AND3_X1   g1205(.A1(new_n1400), .A2(new_n1403), .A3(new_n1320), .ZN(new_n1406));
  AOI21_X1  g1206(.A(new_n1403), .B1(new_n1400), .B2(new_n1320), .ZN(new_n1407));
  OAI21_X1  g1207(.A(new_n1393), .B1(new_n1406), .B2(new_n1407), .ZN(new_n1408));
  AND2_X1   g1208(.A1(new_n1405), .A2(new_n1408), .ZN(G402));
endmodule


