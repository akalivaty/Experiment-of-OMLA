//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g029(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  OR4_X1    g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G567), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(new_n456), .B2(G2106), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(new_n461), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n474), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n484), .B2(G112), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT70), .B1(new_n469), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n480), .A2(new_n488), .A3(new_n484), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(new_n490), .B2(G136), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n491), .B(new_n492), .ZN(G162));
  NAND2_X1  g068(.A1(new_n472), .A2(G102), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G126), .B1(new_n467), .B2(new_n468), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n484), .C1(new_n467), .C2(new_n468), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n480), .A2(new_n502), .A3(G138), .A4(new_n484), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n509), .A2(new_n511), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(new_n518), .A3(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR3_X1    g098(.A1(new_n515), .A2(KEYINPUT72), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT72), .B1(new_n515), .B2(new_n523), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(G166));
  AND2_X1   g101(.A1(new_n516), .A2(new_n518), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n512), .A2(new_n527), .A3(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n527), .A2(G51), .A3(G543), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n509), .A2(new_n511), .A3(G63), .A4(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n509), .A2(new_n511), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  INV_X1    g114(.A(new_n519), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G90), .ZN(new_n541));
  INV_X1    g116(.A(new_n521), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G52), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  INV_X1    g121(.A(G68), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n536), .A2(new_n546), .B1(new_n547), .B2(new_n508), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI221_X1 g125(.A(KEYINPUT73), .B1(new_n547), .B2(new_n508), .C1(new_n536), .C2(new_n546), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(G651), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT74), .B(G81), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n540), .A2(new_n553), .B1(new_n542), .B2(G43), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n516), .A2(new_n518), .A3(G53), .A4(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n536), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n540), .A2(G91), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(G166), .ZN(G303));
  NAND2_X1  g146(.A1(new_n542), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n512), .A2(new_n527), .A3(G87), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G288));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n519), .A2(new_n579), .B1(new_n521), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n509), .A2(new_n511), .A3(G61), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n507), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(KEYINPUT76), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(KEYINPUT76), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n507), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n519), .A2(new_n591), .B1(new_n521), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  INV_X1    g172(.A(G79), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n536), .A2(new_n597), .B1(new_n598), .B2(new_n508), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI221_X1 g176(.A(KEYINPUT77), .B1(new_n598), .B2(new_n508), .C1(new_n536), .C2(new_n597), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n601), .A2(G651), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n542), .A2(G54), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n519), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n512), .A2(new_n527), .A3(KEYINPUT10), .A4(G92), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n603), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n596), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n596), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  AND3_X1   g189(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G860), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n610), .B1(G559), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT78), .Z(G148));
  OR2_X1    g195(.A1(new_n610), .A2(G559), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(KEYINPUT79), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(KEYINPUT79), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n623), .B(new_n624), .C1(G868), .C2(new_n556), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT80), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n480), .A2(new_n472), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT13), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n490), .A2(G135), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n484), .A2(G111), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n471), .B1(new_n633), .B2(KEYINPUT81), .ZN(new_n634));
  OAI221_X1 g209(.A(new_n634), .B1(KEYINPUT81), .B2(new_n633), .C1(G99), .C2(G2105), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n480), .A2(G123), .A3(G2105), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n631), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT84), .B(G2438), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2443), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2446), .Z(new_n651));
  OR2_X1    g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n641), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n640), .A3(new_n656), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n661), .A3(G14), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT85), .ZN(new_n665));
  XOR2_X1   g240(.A(G2067), .B(G2678), .Z(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT18), .ZN(new_n668));
  NOR2_X1   g243(.A1(G2072), .A2(G2078), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n444), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n671), .A3(KEYINPUT17), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT86), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT87), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(new_n687), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n684), .A2(new_n691), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n690), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1981), .B(G1986), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g276(.A1(new_n690), .A2(new_n697), .A3(new_n694), .A4(new_n695), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(new_n699), .B2(new_n702), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n680), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n705), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n707), .A2(new_n679), .A3(new_n703), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n706), .A2(new_n708), .ZN(G229));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G6), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G305), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT32), .B(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G22), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G166), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1971), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n710), .A2(G23), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT89), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n575), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(KEYINPUT89), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n719), .B1(new_n723), .B2(new_n710), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT33), .B(G1976), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n714), .A2(new_n718), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT34), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n714), .A2(new_n718), .A3(new_n729), .A4(new_n726), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n490), .A2(G131), .ZN(new_n733));
  INV_X1    g308(.A(G119), .ZN(new_n734));
  NOR2_X1   g309(.A1(G95), .A2(G2105), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(new_n484), .B2(G107), .ZN(new_n736));
  OAI22_X1  g311(.A1(new_n481), .A2(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n732), .B1(new_n738), .B2(new_n731), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n710), .A2(G24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n594), .B2(new_n710), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT88), .B(G1986), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n728), .A2(new_n730), .A3(new_n741), .A4(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT91), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n731), .A2(G27), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n731), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT97), .B(G2078), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT98), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n753), .B(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n750), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n746), .A2(new_n757), .A3(new_n747), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n472), .A2(G105), .ZN(new_n759));
  INV_X1    g334(.A(G129), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n481), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n490), .B2(G141), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT26), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  MUX2_X1   g341(.A(G32), .B(new_n766), .S(G29), .Z(new_n767));
  XOR2_X1   g342(.A(KEYINPUT27), .B(G1996), .Z(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n710), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n710), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G1966), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n769), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n772), .A2(G1966), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n556), .A2(G16), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G16), .B2(G19), .ZN(new_n777));
  INV_X1    g352(.A(G1341), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(KEYINPUT24), .A2(G34), .ZN(new_n780));
  NOR2_X1   g355(.A1(KEYINPUT24), .A2(G34), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n780), .A2(new_n781), .A3(G29), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n478), .B2(G29), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  INV_X1    g361(.A(G1961), .ZN(new_n787));
  OAI21_X1  g362(.A(KEYINPUT96), .B1(G5), .B2(G16), .ZN(new_n788));
  OR3_X1    g363(.A1(KEYINPUT96), .A2(G5), .A3(G16), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n788), .B(new_n789), .C1(G301), .C2(new_n710), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n790), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n774), .A2(new_n775), .A3(new_n779), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT31), .B(G11), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(G28), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(G28), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n795), .A2(new_n796), .A3(new_n731), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n793), .B(new_n797), .C1(new_n637), .C2(new_n731), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n777), .A2(new_n778), .ZN(new_n800));
  OR2_X1    g375(.A1(G29), .A2(G33), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n490), .A2(G139), .ZN(new_n802));
  NAND2_X1  g377(.A1(G115), .A2(G2104), .ZN(new_n803));
  INV_X1    g378(.A(G127), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n469), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G2105), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT94), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n484), .A2(G2104), .ZN(new_n808));
  INV_X1    g383(.A(G103), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT93), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n472), .A2(new_n811), .A3(G103), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT25), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n810), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n805), .A2(new_n818), .A3(G2105), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n802), .A2(new_n807), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n801), .B1(new_n820), .B2(new_n731), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n799), .B(new_n800), .C1(new_n442), .C2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n442), .B2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n790), .A2(new_n787), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n710), .A2(G20), .ZN(new_n825));
  OAI211_X1 g400(.A(KEYINPUT23), .B(new_n825), .C1(new_n615), .C2(new_n710), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(KEYINPUT23), .B2(new_n825), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1956), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n792), .A2(new_n823), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(G162), .A2(G29), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G29), .B2(G35), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT29), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT29), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n830), .B(new_n833), .C1(G29), .C2(G35), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G2090), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n731), .A2(G26), .ZN(new_n838));
  INV_X1    g413(.A(G128), .ZN(new_n839));
  NOR2_X1   g414(.A1(G104), .A2(G2105), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(new_n484), .B2(G116), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n481), .A2(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n490), .B2(G140), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n838), .B1(new_n843), .B2(new_n731), .ZN(new_n844));
  MUX2_X1   g419(.A(new_n838), .B(new_n844), .S(KEYINPUT28), .Z(new_n845));
  INV_X1    g420(.A(G2067), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT92), .B1(G4), .B2(G16), .ZN(new_n848));
  OR3_X1    g423(.A1(KEYINPUT92), .A2(G4), .A3(G16), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n848), .B(new_n849), .C1(new_n610), .C2(new_n710), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G1348), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n832), .A2(G2090), .A3(new_n834), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n837), .A2(new_n847), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n829), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n751), .A2(new_n756), .A3(new_n758), .A4(new_n854), .ZN(G150));
  NAND2_X1  g430(.A1(G150), .A2(KEYINPUT99), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n758), .A2(new_n854), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n857), .A2(new_n858), .A3(new_n756), .A4(new_n751), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(G311));
  NAND3_X1  g435(.A1(new_n509), .A2(new_n511), .A3(G67), .ZN(new_n861));
  NAND2_X1  g436(.A1(G80), .A2(G543), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n507), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n540), .A2(G93), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT100), .B(G55), .Z(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(new_n521), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT101), .A4(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n869));
  INV_X1    g444(.A(G93), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n519), .A2(new_n870), .B1(new_n866), .B2(new_n521), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n871), .B2(new_n863), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(new_n618), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n611), .A2(G559), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT38), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n868), .A2(new_n872), .B1(new_n552), .B2(new_n554), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n879), .A2(new_n552), .A3(new_n554), .ZN(new_n880));
  OAI21_X1  g455(.A(KEYINPUT102), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(new_n555), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n877), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT39), .ZN(new_n887));
  AOI21_X1  g462(.A(G860), .B1(new_n887), .B2(KEYINPUT103), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(KEYINPUT103), .B2(new_n887), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n886), .A2(KEYINPUT39), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n875), .B1(new_n889), .B2(new_n890), .ZN(G145));
  XNOR2_X1  g466(.A(new_n637), .B(G160), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G162), .ZN(new_n893));
  XNOR2_X1  g468(.A(G164), .B(new_n843), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n807), .A2(new_n819), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n802), .A4(new_n817), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n820), .A2(KEYINPUT105), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n897), .A2(new_n629), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n629), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n894), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n898), .ZN(new_n902));
  INV_X1    g477(.A(new_n629), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n897), .A2(new_n629), .A3(new_n898), .ZN(new_n905));
  INV_X1    g480(.A(new_n894), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(KEYINPUT104), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(KEYINPUT104), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n909), .B(new_n910), .C1(G118), .C2(new_n484), .ZN(new_n911));
  INV_X1    g486(.A(G130), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n912), .B2(new_n481), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(G142), .B2(new_n490), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n733), .B2(new_n737), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n490), .A2(G142), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n738), .B1(new_n916), .B2(new_n913), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n915), .A2(new_n917), .A3(new_n766), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n766), .B1(new_n915), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n901), .A2(new_n907), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n907), .B2(new_n901), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n893), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n901), .A2(new_n907), .ZN(new_n924));
  INV_X1    g499(.A(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n901), .A2(new_n907), .A3(new_n920), .ZN(new_n927));
  INV_X1    g502(.A(new_n893), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n923), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g507(.A1(G305), .A2(KEYINPUT108), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(new_n586), .B2(new_n587), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n524), .A2(new_n525), .A3(new_n721), .A4(new_n722), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n524), .A2(new_n525), .B1(new_n721), .B2(new_n722), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n938), .A2(new_n594), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(G166), .A2(new_n723), .ZN(new_n941));
  AOI21_X1  g516(.A(G290), .B1(new_n941), .B2(new_n937), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n936), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n594), .B1(new_n938), .B2(new_n939), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n933), .A2(new_n935), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(G290), .A3(new_n937), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT42), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n948), .B(KEYINPUT109), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n885), .B(new_n621), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n610), .A2(new_n615), .ZN(new_n956));
  NAND4_X1  g531(.A1(G299), .A2(new_n604), .A3(new_n603), .A4(new_n609), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT41), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT106), .ZN(new_n961));
  INV_X1    g536(.A(new_n958), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n958), .A2(new_n965), .A3(new_n959), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n955), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n955), .B2(new_n962), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n951), .A2(new_n954), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n951), .B2(new_n954), .ZN(new_n971));
  OAI21_X1  g546(.A(G868), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n873), .A2(G868), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(G295));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n973), .ZN(G331));
  AND2_X1   g550(.A1(G286), .A2(KEYINPUT110), .ZN(new_n976));
  NOR2_X1   g551(.A1(G286), .A2(KEYINPUT110), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(G301), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n528), .A2(new_n530), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n529), .A4(new_n532), .ZN(new_n981));
  NAND2_X1  g556(.A1(G286), .A2(KEYINPUT110), .ZN(new_n982));
  AOI21_X1  g557(.A(G171), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n978), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n879), .A2(new_n552), .A3(new_n554), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n883), .B1(new_n882), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n878), .A2(KEYINPUT102), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(G301), .B1(new_n976), .B2(new_n977), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n981), .A2(G171), .A3(new_n982), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n881), .A2(new_n991), .A3(new_n884), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(KEYINPUT111), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n885), .A2(new_n994), .A3(new_n984), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n993), .A2(new_n967), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n988), .A2(new_n958), .A3(new_n992), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n948), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n930), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n948), .B1(new_n996), .B2(new_n997), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT43), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n962), .B1(new_n993), .B2(new_n995), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n958), .A2(KEYINPUT41), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n958), .A2(new_n963), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n1003), .B(new_n1004), .C1(new_n988), .C2(new_n992), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n947), .B(new_n943), .C1(new_n1002), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1006), .A2(new_n1007), .A3(new_n930), .A4(new_n998), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1001), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(new_n930), .A3(new_n998), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(new_n1012), .B2(KEYINPUT43), .ZN(new_n1013));
  OR3_X1    g588(.A1(new_n999), .A2(KEYINPUT43), .A3(new_n1000), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1011), .B1(new_n1016), .B2(new_n1017), .ZN(G397));
  NAND3_X1  g593(.A1(new_n473), .A2(G40), .A3(new_n477), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n501), .A2(new_n503), .ZN(new_n1022));
  INV_X1    g597(.A(new_n497), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n480), .B2(G126), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n494), .B1(new_n1024), .B2(new_n484), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1020), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT113), .Z(new_n1029));
  XNOR2_X1  g604(.A(new_n843), .B(new_n846), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1028), .A2(G1996), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n766), .ZN(new_n1034));
  INV_X1    g609(.A(G1996), .ZN(new_n1035));
  OAI221_X1 g610(.A(new_n1031), .B1(new_n766), .B2(new_n1033), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n738), .B(new_n740), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1037), .B2(new_n1029), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1028), .A2(G1986), .A3(G290), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n1039), .B(KEYINPUT48), .Z(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1032), .B1(KEYINPUT126), .B2(KEYINPUT46), .ZN(new_n1042));
  NOR2_X1   g617(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1043));
  AND2_X1   g618(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1034), .A2(new_n1031), .A3(new_n1042), .A4(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT47), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n843), .A2(new_n846), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n738), .A2(new_n740), .ZN(new_n1049));
  XOR2_X1   g624(.A(new_n1049), .B(KEYINPUT125), .Z(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1036), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1029), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1041), .A2(new_n1047), .A3(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT115), .B1(new_n505), .B2(new_n1021), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n1057), .B(G1384), .C1(new_n499), .C2(new_n504), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1055), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1019), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1059), .A2(new_n784), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1026), .A2(new_n1057), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1384), .B1(new_n499), .B2(new_n504), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT115), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1027), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n1021), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1020), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1966), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G8), .ZN(new_n1071));
  NOR2_X1   g646(.A1(G168), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT51), .B1(new_n1072), .B2(KEYINPUT121), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1059), .A2(new_n784), .A3(new_n1060), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1067), .B1(new_n1078), .B2(new_n1027), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1079), .B2(G1966), .ZN(new_n1080));
  OAI211_X1 g655(.A(G8), .B(new_n1074), .C1(new_n1080), .C2(G286), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(G8), .A3(G286), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1076), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT62), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n581), .A2(G1981), .A3(new_n584), .ZN(new_n1085));
  OAI21_X1  g660(.A(G1981), .B1(new_n581), .B2(new_n584), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1088), .A2(KEYINPUT118), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(KEYINPUT118), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(KEYINPUT118), .A3(new_n1088), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1020), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G8), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1976), .B1(new_n576), .B2(new_n577), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1098), .A3(G8), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n723), .A2(G1976), .ZN(new_n1103));
  AND4_X1   g678(.A1(new_n1102), .A2(new_n1095), .A3(G8), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1095), .A2(new_n1103), .A3(new_n1102), .A4(G8), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n1100), .A3(new_n1099), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1097), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(G166), .A2(new_n1071), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT55), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1019), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1066), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1063), .A2(KEYINPUT114), .A3(KEYINPUT45), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n717), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(G2090), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1110), .A2(new_n1118), .A3(G8), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1062), .A2(new_n1064), .A3(new_n1054), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1120), .A2(new_n836), .A3(new_n1020), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(G8), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT55), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1109), .B(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1108), .A2(new_n1119), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1117), .A2(new_n787), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1111), .A2(new_n1113), .A3(new_n443), .A4(new_n1114), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1079), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1134));
  AOI21_X1  g709(.A(G301), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1076), .A2(new_n1081), .A3(new_n1136), .A4(new_n1082), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1084), .A2(new_n1128), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1139));
  INV_X1    g714(.A(G1966), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g716(.A(new_n1071), .B(G286), .C1(new_n1141), .C2(new_n1077), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1108), .A2(new_n1127), .A3(new_n1119), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1118), .A2(G8), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1144), .B1(new_n1146), .B2(new_n1126), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1147), .A2(new_n1119), .A3(new_n1108), .A4(new_n1142), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(G1976), .ZN(new_n1150));
  INV_X1    g725(.A(G288), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1150), .B(new_n1151), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1096), .B1(new_n1152), .B2(new_n1085), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1119), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n1108), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1138), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1128), .A2(new_n1083), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1158), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1111), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(new_n1132), .A3(new_n1129), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(G171), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT124), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1133), .A2(G301), .A3(new_n1134), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1160), .A2(new_n1164), .A3(G171), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1162), .A2(KEYINPUT54), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1167));
  NOR2_X1   g742(.A1(new_n1160), .A2(G171), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(new_n1135), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT57), .ZN(new_n1171));
  NAND2_X1  g746(.A1(G299), .A2(KEYINPUT119), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(G299), .A2(KEYINPUT119), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1174), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1176), .A2(KEYINPUT57), .A3(new_n1172), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1120), .A2(new_n1020), .A3(new_n1121), .ZN(new_n1179));
  INV_X1    g754(.A(G1956), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT56), .B(G2072), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1158), .A2(new_n1111), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1178), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1181), .A2(new_n1183), .A3(new_n1178), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(KEYINPUT61), .B1(new_n1186), .B2(new_n1184), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1178), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1190), .A2(new_n1191), .A3(new_n1185), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT59), .ZN(new_n1194));
  XOR2_X1   g769(.A(KEYINPUT58), .B(G1341), .Z(new_n1195));
  NAND2_X1  g770(.A1(new_n1095), .A2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(KEYINPUT120), .B(G1996), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1194), .B1(new_n1199), .B2(new_n556), .ZN(new_n1200));
  AOI211_X1 g775(.A(KEYINPUT59), .B(new_n555), .C1(new_n1196), .C2(new_n1198), .ZN(new_n1201));
  AOI21_X1  g776(.A(G1348), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n846), .B(new_n1020), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1203), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT60), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n611), .A2(new_n1206), .ZN(new_n1207));
  OAI22_X1  g782(.A1(new_n1200), .A2(new_n1201), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  OR3_X1    g783(.A1(new_n1202), .A2(new_n611), .A3(new_n1204), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n611), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1206), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1184), .B1(new_n1193), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1185), .A2(new_n611), .A3(new_n1205), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1170), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1156), .B1(new_n1157), .B2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n594), .B(G1986), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1038), .B1(new_n1028), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1053), .B1(new_n1216), .B2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g794(.A1(new_n931), .A2(new_n662), .A3(new_n677), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n465), .B1(new_n706), .B2(new_n708), .ZN(new_n1222));
  NAND3_X1  g796(.A1(new_n1009), .A2(new_n1221), .A3(new_n1222), .ZN(G225));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n1224));
  NAND2_X1  g798(.A1(G225), .A2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g799(.A1(new_n1009), .A2(new_n1221), .A3(new_n1222), .A4(KEYINPUT127), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n1225), .A2(new_n1226), .ZN(G308));
endmodule


