//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n638, new_n640,
    new_n641, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1232;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT65), .A3(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n467), .A2(G137), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT66), .B1(new_n468), .B2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G101), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n470), .A2(KEYINPUT67), .A3(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n481), .A2(new_n469), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n482), .A2(G125), .ZN(new_n483));
  AND2_X1   g058(.A1(G113), .A2(G2104), .ZN(new_n484));
  OAI21_X1  g059(.A(G2105), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n480), .A2(new_n485), .ZN(G160));
  NAND3_X1  g061(.A1(new_n467), .A2(G2105), .A3(new_n469), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  OR2_X1    g067(.A1(G100), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G162));
  NAND4_X1  g071(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n498), .B1(new_n497), .B2(new_n500), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT4), .A2(G138), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n481), .A2(new_n469), .A3(G138), .A4(new_n468), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n501), .A2(new_n502), .A3(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n511), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(G543), .B1(new_n514), .B2(new_n515), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT69), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n511), .A2(new_n513), .ZN(new_n527));
  INV_X1    g102(.A(G62), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n523), .A2(new_n525), .B1(G651), .B2(new_n529), .ZN(G166));
  OAI21_X1  g105(.A(G89), .B1(new_n514), .B2(new_n515), .ZN(new_n531));
  INV_X1    g106(.A(G63), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n527), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n534), .A2(new_n535), .B1(new_n520), .B2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  OAI211_X1 g115(.A(G52), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n516), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n511), .A2(new_n513), .A3(G64), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n533), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT70), .B1(new_n543), .B2(new_n548), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(G171));
  OAI211_X1 g127(.A(G43), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n516), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n511), .A2(new_n513), .A3(G56), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n533), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  NAND3_X1  g140(.A1(new_n511), .A2(new_n513), .A3(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n568), .A2(KEYINPUT72), .A3(G651), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n571), .A2(new_n572), .B1(G91), .B2(new_n517), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n519), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n575), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n520), .A2(G53), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n573), .A2(new_n577), .A3(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n517), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n520), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT73), .Z(G288));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT74), .B1(new_n527), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n511), .A2(new_n513), .A3(new_n592), .A4(G61), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n520), .A2(G48), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n516), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n594), .A2(KEYINPUT75), .A3(G651), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT76), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G651), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n520), .A2(G47), .ZN(new_n607));
  INV_X1    g182(.A(G85), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n516), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n607), .B(KEYINPUT77), .C1(new_n608), .C2(new_n516), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n617));
  OR3_X1    g192(.A1(new_n516), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n527), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G651), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n520), .A2(G54), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n516), .B2(new_n616), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n618), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT79), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n615), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n615), .B1(new_n626), .B2(G868), .ZN(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  INV_X1    g204(.A(G91), .ZN(new_n630));
  AOI21_X1  g205(.A(KEYINPUT72), .B1(new_n568), .B2(G651), .ZN(new_n631));
  AOI211_X1 g206(.A(new_n570), .B(new_n533), .C1(new_n566), .C2(new_n567), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n577), .B1(new_n630), .B2(new_n516), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n580), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n629), .B1(new_n635), .B2(G868), .ZN(G297));
  OAI21_X1  g211(.A(new_n629), .B1(new_n635), .B2(G868), .ZN(G280));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n626), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n626), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(G868), .B2(new_n559), .ZN(G323));
  XOR2_X1   g217(.A(G323), .B(KEYINPUT80), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g219(.A(new_n471), .B(new_n472), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(new_n482), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  INV_X1    g222(.A(G2100), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n488), .A2(G123), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n491), .A2(G135), .ZN(new_n653));
  NOR2_X1   g228(.A1(G99), .A2(G2105), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2096), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n651), .A2(new_n657), .ZN(G156));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2435), .ZN(new_n660));
  XOR2_X1   g235(.A(G2427), .B(G2438), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT14), .ZN(new_n663));
  XOR2_X1   g238(.A(G2451), .B(G2454), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n663), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2443), .B(G2446), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OR3_X1    g246(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n668), .B2(new_n669), .ZN(new_n673));
  AND3_X1   g248(.A1(new_n672), .A2(G14), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT82), .ZN(G401));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2072), .B(G2078), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT83), .ZN(new_n679));
  XOR2_X1   g254(.A(G2067), .B(G2678), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(KEYINPUT84), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT17), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n677), .B(new_n681), .C1(new_n683), .C2(new_n680), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n680), .A3(new_n676), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n680), .A3(new_n677), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT18), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2096), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n689), .A2(new_n648), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n648), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G227));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT85), .ZN(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT86), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1971), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT19), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n695), .A2(new_n697), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(new_n700), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n698), .A2(new_n700), .A3(new_n703), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n705), .B(new_n706), .C1(new_n702), .C2(new_n704), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1981), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT87), .B(G1986), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(G229));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G35), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G162), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT29), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(G2090), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n720), .A2(KEYINPUT23), .A3(G20), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n722));
  INV_X1    g297(.A(G20), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G16), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n721), .B(new_n724), .C1(new_n635), .C2(new_n720), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1956), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n719), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n718), .A2(G2090), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n645), .A2(G105), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT96), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n488), .A2(G129), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n491), .A2(G141), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT97), .B(KEYINPUT26), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n737), .B(new_n738), .Z(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n736), .A2(KEYINPUT98), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n735), .B2(new_n739), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G29), .ZN(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G32), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT27), .B(G1996), .Z(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n748), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n715), .B1(new_n741), .B2(new_n743), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n746), .ZN(new_n752));
  NAND2_X1  g327(.A1(G171), .A2(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G5), .B2(G16), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G1961), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G1961), .ZN(new_n756));
  NOR2_X1   g331(.A1(G164), .A2(new_n715), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G27), .B2(new_n715), .ZN(new_n758));
  INV_X1    g333(.A(G2078), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n755), .A2(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G16), .A2(G21), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G168), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT30), .B(G28), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n762), .A2(G1966), .B1(new_n715), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n749), .A2(new_n752), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n656), .A2(new_n715), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n762), .A2(G1966), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT24), .A2(G34), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n770), .A2(new_n715), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G160), .B2(new_n715), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2084), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n715), .A2(G33), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT25), .Z(new_n777));
  INV_X1    g352(.A(G139), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n777), .B1(new_n490), .B2(new_n778), .C1(new_n779), .C2(new_n468), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n775), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2072), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G11), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n782), .B(new_n783), .C1(new_n758), .C2(new_n759), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n774), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n766), .A2(new_n767), .A3(new_n769), .A4(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n785), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n765), .A2(new_n789), .A3(new_n768), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n790), .A2(KEYINPUT99), .A3(new_n767), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n729), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n720), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(new_n587), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n720), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n795), .A2(KEYINPUT33), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(KEYINPUT33), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G6), .B(G305), .S(G16), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n720), .A2(G22), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G166), .B2(new_n720), .ZN(new_n805));
  INV_X1    g380(.A(G1971), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n800), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT34), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n800), .A2(new_n803), .A3(new_n810), .A4(new_n807), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n488), .A2(G119), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n491), .A2(G131), .ZN(new_n813));
  NOR2_X1   g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(new_n468), .B2(G107), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT88), .ZN(new_n817));
  MUX2_X1   g392(.A(G25), .B(new_n817), .S(G29), .Z(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT35), .B(G1991), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT89), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G24), .B(G290), .S(G16), .Z(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT90), .B(G1986), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n809), .A2(new_n811), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(KEYINPUT91), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n720), .A2(G19), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n559), .B2(new_n720), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT94), .B(G1341), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n720), .A2(G4), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n626), .B2(new_n720), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT92), .B(G1348), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT93), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n834), .B(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n792), .A2(new_n828), .A3(new_n832), .A4(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT28), .ZN(new_n839));
  INV_X1    g414(.A(G26), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(G29), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(G29), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n488), .A2(G128), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n491), .A2(G140), .ZN(new_n844));
  NOR2_X1   g419(.A1(G104), .A2(G2105), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n842), .B1(new_n847), .B2(G29), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n841), .B1(new_n848), .B2(new_n839), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT95), .B(G2067), .Z(new_n850));
  XOR2_X1   g425(.A(new_n849), .B(new_n850), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n838), .A2(new_n851), .ZN(G311));
  AND2_X1   g427(.A1(new_n792), .A2(new_n828), .ZN(new_n853));
  INV_X1    g428(.A(new_n851), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n832), .A4(new_n837), .ZN(G150));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  INV_X1    g431(.A(G67), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n527), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G651), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g436(.A(G55), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n862));
  INV_X1    g437(.A(G93), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n516), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n858), .A2(KEYINPUT100), .A3(G651), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n861), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n626), .A2(G559), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT39), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n858), .A2(KEYINPUT100), .A3(G651), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT100), .B1(new_n858), .B2(G651), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n873), .A2(new_n874), .A3(new_n864), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT101), .B1(new_n555), .B2(new_n558), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n559), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n559), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n867), .A2(KEYINPUT101), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n872), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n869), .B1(new_n884), .B2(G860), .ZN(G145));
  NAND4_X1  g460(.A1(new_n504), .A2(new_n497), .A3(new_n507), .A4(new_n500), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n816), .B(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(G160), .A2(new_n656), .ZN(new_n888));
  NAND2_X1  g463(.A1(G160), .A2(new_n656), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(G162), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(G162), .B1(new_n888), .B2(new_n889), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  INV_X1    g469(.A(new_n887), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n890), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n736), .A2(new_n780), .A3(new_n740), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n744), .B2(new_n780), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n893), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n893), .B2(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n488), .A2(G130), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n491), .A2(G142), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n468), .A2(G118), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT102), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n904), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n647), .B(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n847), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  OR3_X1    g484(.A1(new_n899), .A2(new_n900), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n899), .B2(new_n900), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g489(.A1(G305), .A2(new_n794), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n597), .A2(new_n587), .A3(new_n601), .A4(new_n602), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(G303), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(G290), .A2(KEYINPUT104), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n606), .A2(new_n613), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G303), .B1(new_n915), .B2(new_n916), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n606), .A2(new_n613), .A3(new_n920), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n606), .B2(new_n613), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n923), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n917), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT42), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n883), .B(new_n640), .ZN(new_n932));
  INV_X1    g507(.A(new_n625), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n633), .B2(new_n634), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n573), .A2(new_n577), .A3(new_n580), .A4(new_n625), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT41), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n635), .A2(KEYINPUT103), .A3(new_n625), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n932), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(new_n932), .B2(new_n936), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n931), .B(new_n945), .Z(new_n946));
  MUX2_X1   g521(.A(new_n867), .B(new_n946), .S(G868), .Z(G295));
  MUX2_X1   g522(.A(new_n867), .B(new_n946), .S(G868), .Z(G331));
  NAND2_X1  g523(.A1(G171), .A2(G168), .ZN(new_n949));
  NAND3_X1  g524(.A1(G286), .A2(new_n550), .A3(new_n551), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n882), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n879), .A2(new_n949), .A3(new_n881), .A4(new_n950), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n954), .A2(new_n937), .A3(new_n942), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(new_n936), .A3(new_n953), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n929), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n928), .A2(new_n927), .A3(new_n917), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(KEYINPUT41), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n936), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n954), .A2(KEYINPUT41), .A3(new_n941), .A4(new_n939), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n962), .B(new_n963), .C1(new_n924), .C2(new_n929), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n964), .A3(new_n911), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n911), .B1(new_n930), .B2(new_n957), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT105), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n969), .B(new_n911), .C1(new_n930), .C2(new_n957), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n960), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n966), .B1(new_n971), .B2(KEYINPUT43), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n972), .A2(KEYINPUT44), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n968), .A2(new_n974), .A3(new_n960), .A4(new_n970), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(KEYINPUT44), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT106), .B1(new_n965), .B2(KEYINPUT43), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n965), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT107), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n982));
  AOI21_X1  g557(.A(G37), .B1(new_n930), .B2(new_n957), .ZN(new_n983));
  AOI211_X1 g558(.A(new_n982), .B(new_n974), .C1(new_n983), .C2(new_n964), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n975), .B(KEYINPUT44), .C1(new_n984), .C2(new_n977), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n973), .B1(new_n981), .B2(new_n987), .ZN(G397));
  NAND2_X1  g563(.A1(new_n736), .A2(new_n740), .ZN(new_n989));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n886), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n470), .A2(KEYINPUT67), .A3(new_n475), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT67), .B1(new_n470), .B2(new_n475), .ZN(new_n995));
  OAI211_X1 g570(.A(G40), .B(new_n485), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n989), .A2(G1996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1996), .B1(new_n741), .B2(new_n743), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n847), .B(G2067), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n997), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n816), .B(new_n819), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n997), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1000), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(G290), .B(G1986), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1006), .B1(new_n997), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n991), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(new_n480), .A3(G40), .A4(new_n485), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G8), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n597), .A2(new_n1012), .A3(new_n601), .A4(new_n602), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT113), .ZN(new_n1015));
  INV_X1    g590(.A(new_n595), .ZN(new_n1016));
  OAI21_X1  g591(.A(G1981), .B1(new_n1016), .B2(new_n600), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1014), .A2(KEYINPUT113), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1019), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1013), .A2(new_n1017), .A3(new_n1021), .A4(new_n1015), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G288), .A2(G1976), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1011), .B1(new_n1025), .B2(new_n1013), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n794), .A2(G1976), .ZN(new_n1028));
  OAI211_X1 g603(.A(G8), .B(new_n1028), .C1(new_n996), .C2(new_n991), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(KEYINPUT112), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(G288), .A2(new_n1030), .A3(new_n799), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1030), .A2(KEYINPUT112), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1010), .A2(G8), .A3(new_n1028), .A4(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1011), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1027), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT114), .B(new_n1038), .C1(new_n1023), .C2(new_n1011), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n497), .A2(new_n500), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT68), .ZN(new_n1043));
  INV_X1    g618(.A(new_n508), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n990), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n996), .B1(new_n1047), .B2(KEYINPUT50), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT110), .B(G2090), .Z(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n886), .A2(new_n1051), .A3(new_n990), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1048), .A2(new_n1050), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT45), .B1(new_n1046), .B2(new_n990), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n886), .A2(KEYINPUT45), .A3(new_n990), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n480), .A2(new_n1057), .A3(G40), .A4(new_n485), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n806), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1041), .B1(new_n1055), .B2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(G303), .B2(G8), .ZN(new_n1063));
  NOR4_X1   g638(.A1(G166), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(new_n1041), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1026), .B1(new_n1040), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G168), .A2(new_n1041), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT51), .B1(new_n1069), .B2(KEYINPUT122), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1073));
  INV_X1    g648(.A(new_n996), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1052), .A2(KEYINPUT109), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1052), .A2(KEYINPUT109), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G2084), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1046), .A2(KEYINPUT45), .A3(new_n990), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n996), .B1(new_n992), .B2(new_n991), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1046), .A2(KEYINPUT115), .A3(KEYINPUT45), .A4(new_n990), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1966), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1078), .A2(new_n1079), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1070), .B(new_n1072), .C1(new_n1087), .C2(new_n1041), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1048), .A2(new_n1079), .A3(new_n1054), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(G8), .B(new_n1071), .C1(new_n1091), .C2(G286), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(G8), .A3(G286), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT62), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1046), .A2(new_n1051), .A3(new_n990), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(new_n1074), .A3(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n1049), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n992), .B1(G164), .B2(G1384), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n886), .A2(KEYINPUT45), .A3(new_n990), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n996), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1971), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(G8), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1065), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1100), .A2(new_n1111), .A3(new_n1066), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1961), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1077), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1105), .A2(new_n1107), .A3(new_n759), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(G2078), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1115), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1113), .B(new_n1123), .C1(new_n1094), .C2(KEYINPUT62), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1068), .B1(new_n1099), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1091), .A2(G8), .A3(G168), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT63), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1037), .A2(new_n1039), .A3(new_n1066), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1112), .B2(new_n1127), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1040), .A2(new_n1134), .A3(KEYINPUT116), .A4(new_n1066), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n835), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1010), .A2(G2067), .ZN(new_n1139));
  NOR4_X1   g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n626), .ZN(new_n1140));
  NAND2_X1  g715(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n1141));
  OAI221_X1 g716(.A(KEYINPUT117), .B1(new_n630), .B2(new_n516), .C1(new_n631), .C2(new_n632), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n635), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(G299), .A2(new_n1143), .A3(new_n1142), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1141), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(G1956), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1103), .A2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT56), .B(G2072), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1105), .A2(new_n1107), .A3(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1151), .A2(new_n1147), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1147), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1149), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1147), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1151), .A2(new_n1147), .A3(new_n1153), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n1141), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1140), .B1(new_n1156), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1056), .A2(new_n1058), .A3(G1996), .ZN(new_n1164));
  XNOR2_X1  g739(.A(KEYINPUT118), .B(G1341), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT58), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1010), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n559), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1163), .B1(new_n1168), .B2(KEYINPUT59), .ZN(new_n1169));
  INV_X1    g744(.A(G1996), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1105), .A2(new_n1107), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1010), .A2(new_n1166), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n880), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1173), .A2(KEYINPUT120), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(KEYINPUT119), .B1(new_n1168), .B2(KEYINPUT59), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1173), .A2(new_n1177), .A3(new_n1174), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1169), .B(new_n1175), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1138), .ZN(new_n1181));
  OR3_X1    g756(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n626), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1162), .A2(new_n1179), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1180), .A2(new_n626), .A3(new_n1160), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1184), .A2(new_n1185), .A3(new_n1159), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1114), .A2(new_n1077), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1083), .A2(new_n1057), .A3(new_n1119), .ZN(new_n1188));
  AOI21_X1  g763(.A(G301), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AND4_X1   g764(.A1(G301), .A2(new_n1115), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1112), .B1(new_n1191), .B2(KEYINPUT54), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1187), .A2(G301), .A3(new_n1188), .ZN(new_n1193));
  AOI21_X1  g768(.A(KEYINPUT54), .B1(new_n1122), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1194), .A2(KEYINPUT123), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT123), .ZN(new_n1196));
  AOI211_X1 g771(.A(new_n1196), .B(KEYINPUT54), .C1(new_n1122), .C2(new_n1193), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1192), .B(new_n1094), .C1(new_n1195), .C2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1136), .B1(new_n1186), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1008), .B1(new_n1125), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1006), .A2(KEYINPUT126), .ZN(new_n1201));
  INV_X1    g776(.A(new_n997), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1202), .A2(G1986), .A3(G290), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1203), .B(KEYINPUT48), .Z(new_n1204));
  INV_X1    g779(.A(KEYINPUT126), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1000), .A2(new_n1205), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1201), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n997), .A2(new_n1170), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT46), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n997), .B1(new_n989), .B2(new_n1002), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT47), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1207), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n817), .A2(new_n819), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1000), .A2(new_n1003), .A3(new_n1214), .ZN(new_n1215));
  OR2_X1    g790(.A1(new_n847), .A2(G2067), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(KEYINPUT125), .B1(new_n1217), .B2(new_n997), .ZN(new_n1218));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n1219));
  AOI211_X1 g794(.A(new_n1219), .B(new_n1202), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1220));
  OAI211_X1 g795(.A(new_n1213), .B(KEYINPUT127), .C1(new_n1218), .C2(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1207), .A2(new_n1212), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1221), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1200), .A2(new_n1226), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g802(.A(new_n674), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n913), .A2(new_n1229), .A3(new_n692), .ZN(new_n1230));
  NOR4_X1   g804(.A1(new_n1230), .A2(new_n972), .A3(new_n460), .A4(G229), .ZN(G308));
  NOR3_X1   g805(.A1(new_n972), .A2(G229), .A3(new_n460), .ZN(new_n1232));
  NAND4_X1  g806(.A1(new_n1232), .A2(new_n1229), .A3(new_n692), .A4(new_n913), .ZN(G225));
endmodule


