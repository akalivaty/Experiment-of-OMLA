

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590;

  XNOR2_X2 U323 ( .A(n458), .B(KEYINPUT119), .ZN(n459) );
  NOR2_X4 U324 ( .A1(n540), .A2(n459), .ZN(n570) );
  XNOR2_X1 U325 ( .A(n335), .B(n334), .ZN(n337) );
  XNOR2_X1 U326 ( .A(n327), .B(n372), .ZN(n328) );
  NOR2_X1 U327 ( .A1(n576), .A2(n385), .ZN(n387) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U329 ( .A(n418), .B(n291), .ZN(n327) );
  INV_X1 U330 ( .A(KEYINPUT9), .ZN(n332) );
  XNOR2_X1 U331 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U332 ( .A(KEYINPUT47), .B(KEYINPUT108), .ZN(n392) );
  AND2_X1 U333 ( .A1(n477), .A2(n454), .ZN(n455) );
  XNOR2_X1 U334 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U335 ( .A(G36GAT), .B(G218GAT), .Z(n398) );
  XNOR2_X1 U336 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n396) );
  XNOR2_X1 U337 ( .A(KEYINPUT99), .B(KEYINPUT36), .ZN(n345) );
  XOR2_X1 U338 ( .A(n383), .B(n382), .Z(n579) );
  XNOR2_X1 U339 ( .A(n579), .B(KEYINPUT41), .ZN(n560) );
  XNOR2_X1 U340 ( .A(n323), .B(n322), .ZN(n576) );
  XNOR2_X1 U341 ( .A(KEYINPUT92), .B(n483), .ZN(n526) );
  XNOR2_X1 U342 ( .A(n461), .B(G190GAT), .ZN(n462) );
  XNOR2_X1 U343 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U345 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n292) );
  XNOR2_X1 U346 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U347 ( .A(n294), .B(G183GAT), .Z(n296) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(G176GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n406) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n297), .B(G120GAT), .ZN(n430) );
  XOR2_X1 U352 ( .A(KEYINPUT80), .B(n430), .Z(n299) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U355 ( .A(G127GAT), .B(KEYINPUT20), .Z(n301) );
  XNOR2_X1 U356 ( .A(G15GAT), .B(KEYINPUT79), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U358 ( .A(n303), .B(n302), .Z(n305) );
  XOR2_X1 U359 ( .A(G43GAT), .B(G134GAT), .Z(n329) );
  XOR2_X1 U360 ( .A(G99GAT), .B(G71GAT), .Z(n375) );
  XNOR2_X1 U361 ( .A(n329), .B(n375), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n406), .B(n306), .ZN(n540) );
  XOR2_X1 U364 ( .A(G197GAT), .B(G141GAT), .Z(n308) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G113GAT), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U367 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n310) );
  XNOR2_X1 U368 ( .A(G8GAT), .B(G1GAT), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n323) );
  XOR2_X1 U371 ( .A(G50GAT), .B(G22GAT), .Z(n446) );
  XOR2_X1 U372 ( .A(G15GAT), .B(G36GAT), .Z(n314) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(G43GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U375 ( .A(n446), .B(n315), .Z(n317) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U378 ( .A(n318), .B(KEYINPUT29), .Z(n321) );
  XNOR2_X1 U379 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n319), .B(KEYINPUT65), .ZN(n340) );
  XNOR2_X1 U381 ( .A(n340), .B(KEYINPUT64), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U383 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n325) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G162GAT), .ZN(n324) );
  XOR2_X1 U385 ( .A(n325), .B(n324), .Z(n344) );
  XOR2_X1 U386 ( .A(G29GAT), .B(G85GAT), .Z(n418) );
  XNOR2_X1 U387 ( .A(G106GAT), .B(KEYINPUT68), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n326), .B(KEYINPUT69), .ZN(n372) );
  XNOR2_X1 U389 ( .A(G50GAT), .B(n328), .ZN(n335) );
  XOR2_X1 U390 ( .A(G92GAT), .B(n398), .Z(n331) );
  XNOR2_X1 U391 ( .A(G190GAT), .B(n329), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n333) );
  INV_X1 U393 ( .A(KEYINPUT10), .ZN(n336) );
  NAND2_X1 U394 ( .A1(n337), .A2(n336), .ZN(n339) );
  OR2_X1 U395 ( .A1(n337), .A2(n336), .ZN(n338) );
  NAND2_X1 U396 ( .A1(n339), .A2(n338), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n340), .B(KEYINPUT11), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n460) );
  XNOR2_X1 U400 ( .A(n460), .B(n345), .ZN(n587) );
  XOR2_X1 U401 ( .A(G78GAT), .B(G71GAT), .Z(n347) );
  XNOR2_X1 U402 ( .A(G15GAT), .B(G183GAT), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U404 ( .A(G8GAT), .B(KEYINPUT74), .Z(n402) );
  XOR2_X1 U405 ( .A(n348), .B(n402), .Z(n350) );
  XNOR2_X1 U406 ( .A(G22GAT), .B(G211GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n356) );
  XOR2_X1 U408 ( .A(G57GAT), .B(G155GAT), .Z(n352) );
  XNOR2_X1 U409 ( .A(G1GAT), .B(G127GAT), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n429) );
  XOR2_X1 U411 ( .A(G64GAT), .B(n429), .Z(n354) );
  NAND2_X1 U412 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U414 ( .A(n356), .B(n355), .Z(n364) );
  XOR2_X1 U415 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n358) );
  XNOR2_X1 U416 ( .A(KEYINPUT78), .B(KEYINPUT76), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U418 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n360) );
  XNOR2_X1 U419 ( .A(KEYINPUT13), .B(KEYINPUT12), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n565) );
  NOR2_X1 U423 ( .A1(n587), .A2(n565), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n365), .B(KEYINPUT45), .ZN(n384) );
  XOR2_X1 U425 ( .A(KEYINPUT67), .B(KEYINPUT31), .Z(n367) );
  XNOR2_X1 U426 ( .A(G57GAT), .B(KEYINPUT32), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n383) );
  XOR2_X1 U428 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n369) );
  NAND2_X1 U429 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U431 ( .A(n370), .B(KEYINPUT71), .Z(n374) );
  XNOR2_X1 U432 ( .A(G204GAT), .B(G92GAT), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n371), .B(G64GAT), .ZN(n399) );
  XNOR2_X1 U434 ( .A(n372), .B(n399), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n379) );
  XOR2_X1 U436 ( .A(G148GAT), .B(G78GAT), .Z(n440) );
  XOR2_X1 U437 ( .A(G85GAT), .B(n440), .Z(n377) );
  XNOR2_X1 U438 ( .A(n375), .B(G120GAT), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U440 ( .A(n379), .B(n378), .Z(n381) );
  XNOR2_X1 U441 ( .A(G176GAT), .B(KEYINPUT13), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  NAND2_X1 U443 ( .A1(n384), .A2(n579), .ZN(n385) );
  INV_X1 U444 ( .A(KEYINPUT109), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n395) );
  XOR2_X1 U446 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n389) );
  NAND2_X1 U447 ( .A1(n576), .A2(n560), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U449 ( .A(n565), .B(KEYINPUT106), .Z(n548) );
  NOR2_X1 U450 ( .A1(n460), .A2(n548), .ZN(n390) );
  NAND2_X1 U451 ( .A1(n391), .A2(n390), .ZN(n393) );
  NOR2_X1 U452 ( .A1(n395), .A2(n394), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n539) );
  XOR2_X1 U454 ( .A(n399), .B(n398), .Z(n401) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U457 ( .A(n403), .B(n402), .Z(n408) );
  XOR2_X1 U458 ( .A(G211GAT), .B(KEYINPUT83), .Z(n405) );
  XNOR2_X1 U459 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n442) );
  XNOR2_X1 U461 ( .A(n406), .B(n442), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n528) );
  XOR2_X1 U463 ( .A(KEYINPUT118), .B(n528), .Z(n409) );
  NOR2_X1 U464 ( .A1(n539), .A2(n409), .ZN(n411) );
  INV_X1 U465 ( .A(KEYINPUT54), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n435) );
  XOR2_X1 U467 ( .A(KEYINPUT84), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U468 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U470 ( .A(G141GAT), .B(n414), .ZN(n452) );
  INV_X1 U471 ( .A(n452), .ZN(n422) );
  XOR2_X1 U472 ( .A(KEYINPUT86), .B(KEYINPUT88), .Z(n416) );
  XNOR2_X1 U473 ( .A(G134GAT), .B(G148GAT), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U475 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n434) );
  XOR2_X1 U479 ( .A(KEYINPUT87), .B(KEYINPUT90), .Z(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U482 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n426) );
  XNOR2_X1 U483 ( .A(KEYINPUT91), .B(KEYINPUT6), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U485 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n483) );
  NOR2_X2 U489 ( .A1(n435), .A2(n526), .ZN(n575) );
  XOR2_X1 U490 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n437) );
  XNOR2_X1 U491 ( .A(G155GAT), .B(KEYINPUT85), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n450) );
  XOR2_X1 U493 ( .A(G204GAT), .B(KEYINPUT24), .Z(n439) );
  XNOR2_X1 U494 ( .A(G218GAT), .B(G106GAT), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U496 ( .A(n441), .B(n440), .Z(n448) );
  XOR2_X1 U497 ( .A(n442), .B(KEYINPUT82), .Z(n444) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U502 ( .A(n450), .B(n449), .Z(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n477) );
  NAND2_X1 U504 ( .A1(n575), .A2(n477), .ZN(n453) );
  NAND2_X1 U505 ( .A1(n453), .A2(KEYINPUT55), .ZN(n457) );
  INV_X1 U506 ( .A(KEYINPUT55), .ZN(n454) );
  NAND2_X1 U507 ( .A1(n575), .A2(n455), .ZN(n456) );
  NAND2_X1 U508 ( .A1(n457), .A2(n456), .ZN(n458) );
  NAND2_X1 U509 ( .A1(n570), .A2(n460), .ZN(n463) );
  XOR2_X1 U510 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n461) );
  NAND2_X1 U511 ( .A1(n570), .A2(n548), .ZN(n466) );
  XOR2_X1 U512 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n464) );
  XNOR2_X1 U513 ( .A(n464), .B(G183GAT), .ZN(n465) );
  XNOR2_X1 U514 ( .A(n466), .B(n465), .ZN(G1350GAT) );
  NAND2_X1 U515 ( .A1(n570), .A2(n560), .ZN(n470) );
  XOR2_X1 U516 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n468) );
  XNOR2_X1 U517 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n467) );
  XNOR2_X1 U518 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U519 ( .A(n470), .B(n469), .ZN(G1349GAT) );
  NAND2_X1 U520 ( .A1(n576), .A2(n579), .ZN(n504) );
  NOR2_X1 U521 ( .A1(n460), .A2(n565), .ZN(n471) );
  XNOR2_X1 U522 ( .A(n471), .B(KEYINPUT16), .ZN(n487) );
  XOR2_X1 U523 ( .A(n528), .B(KEYINPUT93), .Z(n472) );
  XNOR2_X1 U524 ( .A(KEYINPUT27), .B(n472), .ZN(n479) );
  NAND2_X1 U525 ( .A1(n479), .A2(n526), .ZN(n473) );
  XOR2_X1 U526 ( .A(KEYINPUT94), .B(n473), .Z(n555) );
  XNOR2_X1 U527 ( .A(n477), .B(KEYINPUT28), .ZN(n497) );
  NAND2_X1 U528 ( .A1(n555), .A2(n497), .ZN(n542) );
  XNOR2_X1 U529 ( .A(KEYINPUT81), .B(n540), .ZN(n474) );
  NOR2_X1 U530 ( .A1(n542), .A2(n474), .ZN(n485) );
  INV_X1 U531 ( .A(n540), .ZN(n531) );
  NAND2_X1 U532 ( .A1(n531), .A2(n528), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n477), .A2(n475), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(KEYINPUT25), .ZN(n481) );
  NOR2_X1 U535 ( .A1(n531), .A2(n477), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT26), .B(n478), .ZN(n574) );
  AND2_X1 U537 ( .A1(n574), .A2(n479), .ZN(n480) );
  NOR2_X1 U538 ( .A1(n481), .A2(n480), .ZN(n482) );
  NOR2_X1 U539 ( .A1(n483), .A2(n482), .ZN(n484) );
  NOR2_X1 U540 ( .A1(n485), .A2(n484), .ZN(n500) );
  INV_X1 U541 ( .A(n500), .ZN(n486) );
  NAND2_X1 U542 ( .A1(n487), .A2(n486), .ZN(n516) );
  NOR2_X1 U543 ( .A1(n504), .A2(n516), .ZN(n498) );
  NAND2_X1 U544 ( .A1(n526), .A2(n498), .ZN(n490) );
  XOR2_X1 U545 ( .A(G1GAT), .B(KEYINPUT34), .Z(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT95), .B(n488), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n490), .B(n489), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n498), .A2(n528), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n491), .B(KEYINPUT96), .ZN(n492) );
  XNOR2_X1 U550 ( .A(G8GAT), .B(n492), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n494) );
  NAND2_X1 U552 ( .A1(n498), .A2(n531), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n496) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT97), .Z(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  INV_X1 U556 ( .A(n497), .ZN(n533) );
  NAND2_X1 U557 ( .A1(n498), .A2(n533), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n499), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .Z(n507) );
  NOR2_X1 U560 ( .A1(n587), .A2(n500), .ZN(n501) );
  NAND2_X1 U561 ( .A1(n565), .A2(n501), .ZN(n502) );
  XNOR2_X1 U562 ( .A(KEYINPUT100), .B(n502), .ZN(n503) );
  XOR2_X1 U563 ( .A(KEYINPUT37), .B(n503), .Z(n525) );
  NOR2_X1 U564 ( .A1(n504), .A2(n525), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n505), .B(KEYINPUT38), .ZN(n513) );
  NAND2_X1 U566 ( .A1(n513), .A2(n526), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  XOR2_X1 U568 ( .A(G36GAT), .B(KEYINPUT101), .Z(n509) );
  NAND2_X1 U569 ( .A1(n528), .A2(n513), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(G1329GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT102), .B(KEYINPUT40), .Z(n511) );
  NAND2_X1 U572 ( .A1(n531), .A2(n513), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U574 ( .A(G43GAT), .B(n512), .Z(G1330GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n533), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n518) );
  INV_X1 U578 ( .A(n576), .ZN(n515) );
  NAND2_X1 U579 ( .A1(n515), .A2(n560), .ZN(n524) );
  NOR2_X1 U580 ( .A1(n524), .A2(n516), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n521), .A2(n526), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n528), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n531), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U588 ( .A1(n521), .A2(n533), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NOR2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n534), .A2(n526), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G85GAT), .B(n527), .ZN(G1336GAT) );
  XOR2_X1 U593 ( .A(G92GAT), .B(KEYINPUT103), .Z(n530) );
  NAND2_X1 U594 ( .A1(n534), .A2(n528), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n534), .A2(n531), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(KEYINPUT104), .ZN(n538) );
  XOR2_X1 U599 ( .A(KEYINPUT44), .B(KEYINPUT105), .Z(n536) );
  NAND2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1339GAT) );
  XOR2_X1 U603 ( .A(G113GAT), .B(KEYINPUT111), .Z(n544) );
  OR2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n542), .A2(n541), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n552), .A2(n576), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U609 ( .A1(n552), .A2(n560), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(n547), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n550) );
  NAND2_X1 U613 ( .A1(n552), .A2(n548), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n554) );
  NAND2_X1 U617 ( .A1(n552), .A2(n460), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1343GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n558) );
  NAND2_X1 U620 ( .A1(n574), .A2(n555), .ZN(n556) );
  NOR2_X1 U621 ( .A1(n539), .A2(n556), .ZN(n568) );
  NAND2_X1 U622 ( .A1(n568), .A2(n576), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(n559), .ZN(G1344GAT) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n562) );
  NAND2_X1 U627 ( .A1(n568), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  XOR2_X1 U630 ( .A(G155GAT), .B(KEYINPUT117), .Z(n567) );
  INV_X1 U631 ( .A(n565), .ZN(n583) );
  NAND2_X1 U632 ( .A1(n568), .A2(n583), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n460), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n576), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G169GAT), .B(n571), .ZN(G1348GAT) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT59), .ZN(n573) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(n573), .Z(n578) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n586) );
  INV_X1 U642 ( .A(n586), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n584), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n581) );
  OR2_X1 U646 ( .A1(n586), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n582), .Z(G1353GAT) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(G218GAT), .B(n590), .Z(G1355GAT) );
endmodule

