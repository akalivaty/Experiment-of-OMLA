

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788;

  AND2_X1 U382 ( .A1(n405), .A2(n406), .ZN(n369) );
  AND2_X1 U383 ( .A1(n770), .A2(n589), .ZN(n407) );
  XNOR2_X1 U384 ( .A(n399), .B(KEYINPUT42), .ZN(n788) );
  AND2_X1 U385 ( .A1(n651), .A2(n362), .ZN(n361) );
  INV_X1 U386 ( .A(n649), .ZN(n362) );
  BUF_X1 U387 ( .A(n629), .Z(n364) );
  XNOR2_X1 U388 ( .A(n629), .B(KEYINPUT38), .ZN(n621) );
  OR2_X1 U389 ( .A1(n622), .A2(n623), .ZN(n422) );
  AND2_X1 U390 ( .A1(G217), .A2(n541), .ZN(n542) );
  BUF_X1 U391 ( .A(n771), .Z(n365) );
  XNOR2_X1 U392 ( .A(n513), .B(n512), .ZN(n515) );
  INV_X1 U393 ( .A(G953), .ZN(n771) );
  NAND2_X1 U394 ( .A1(n363), .A2(n361), .ZN(n653) );
  INV_X1 U395 ( .A(n650), .ZN(n363) );
  XNOR2_X2 U396 ( .A(n422), .B(KEYINPUT106), .ZN(n704) );
  AND2_X2 U397 ( .A1(n402), .A2(n403), .ZN(n397) );
  XNOR2_X2 U398 ( .A(n729), .B(n486), .ZN(n402) );
  NOR2_X2 U399 ( .A1(n650), .A2(n663), .ZN(n483) );
  XNOR2_X1 U400 ( .A(G143), .B(G104), .ZN(n524) );
  INV_X1 U401 ( .A(G146), .ZN(n574) );
  XNOR2_X1 U402 ( .A(n517), .B(KEYINPUT10), .ZN(n767) );
  NOR2_X1 U403 ( .A1(n665), .A2(n658), .ZN(n414) );
  XNOR2_X1 U404 ( .A(n495), .B(G472), .ZN(n607) );
  INV_X1 U405 ( .A(n648), .ZN(n714) );
  XNOR2_X2 U406 ( .A(n468), .B(n388), .ZN(n498) );
  NAND2_X2 U407 ( .A1(n554), .A2(n553), .ZN(n388) );
  NOR2_X2 U408 ( .A1(n498), .A2(G902), .ZN(n555) );
  NAND2_X2 U409 ( .A1(n369), .A2(n404), .ZN(n403) );
  XNOR2_X2 U410 ( .A(n434), .B(n370), .ZN(n648) );
  XNOR2_X2 U411 ( .A(n582), .B(G134), .ZN(n550) );
  XOR2_X2 U412 ( .A(G146), .B(G125), .Z(n584) );
  OR2_X1 U413 ( .A1(n770), .A2(n412), .ZN(n411) );
  AND2_X2 U414 ( .A1(n487), .A2(n508), .ZN(n770) );
  XNOR2_X1 U415 ( .A(n442), .B(n441), .ZN(n782) );
  XNOR2_X1 U416 ( .A(n664), .B(KEYINPUT108), .ZN(n783) );
  XNOR2_X1 U417 ( .A(n393), .B(n615), .ZN(n785) );
  XNOR2_X1 U418 ( .A(n653), .B(n652), .ZN(n779) );
  XNOR2_X1 U419 ( .A(n398), .B(KEYINPUT40), .ZN(n787) );
  XNOR2_X1 U420 ( .A(n414), .B(n376), .ZN(n438) );
  XNOR2_X1 U421 ( .A(n545), .B(n544), .ZN(n622) );
  XNOR2_X1 U422 ( .A(n533), .B(n532), .ZN(n623) );
  XNOR2_X1 U423 ( .A(n747), .B(n509), .ZN(n748) );
  XNOR2_X1 U424 ( .A(n447), .B(n446), .ZN(n563) );
  XNOR2_X1 U425 ( .A(n459), .B(n539), .ZN(n752) );
  XNOR2_X1 U426 ( .A(n450), .B(n760), .ZN(n740) );
  OR2_X1 U427 ( .A1(n372), .A2(n552), .ZN(n554) );
  XNOR2_X1 U428 ( .A(n452), .B(n451), .ZN(n450) );
  XNOR2_X1 U429 ( .A(n421), .B(n415), .ZN(n452) );
  XNOR2_X1 U430 ( .A(n585), .B(n588), .ZN(n451) );
  XNOR2_X1 U431 ( .A(G119), .B(KEYINPUT71), .ZN(n566) );
  XNOR2_X1 U432 ( .A(n582), .B(KEYINPUT4), .ZN(n415) );
  OR2_X1 U433 ( .A1(n607), .A2(n665), .ZN(n721) );
  NOR2_X1 U434 ( .A1(n608), .A2(n658), .ZN(n609) );
  AND2_X1 U435 ( .A1(n630), .A2(n697), .ZN(n508) );
  XNOR2_X1 U436 ( .A(n428), .B(n465), .ZN(n487) );
  XNOR2_X1 U437 ( .A(n433), .B(KEYINPUT70), .ZN(n608) );
  NOR2_X1 U438 ( .A1(G953), .A2(G237), .ZN(n571) );
  NOR2_X1 U439 ( .A1(n387), .A2(n783), .ZN(n383) );
  NOR2_X1 U440 ( .A1(n673), .A2(n706), .ZN(n387) );
  NOR2_X1 U441 ( .A1(n678), .A2(G902), .ZN(n495) );
  INV_X1 U442 ( .A(KEYINPUT2), .ZN(n486) );
  NAND2_X1 U443 ( .A1(n436), .A2(n374), .ZN(n435) );
  AND2_X1 U444 ( .A1(n616), .A2(n489), .ZN(n436) );
  NAND2_X1 U445 ( .A1(n392), .A2(n423), .ZN(n432) );
  AND2_X1 U446 ( .A1(n368), .A2(n599), .ZN(n423) );
  INV_X1 U447 ( .A(n785), .ZN(n392) );
  NAND2_X1 U448 ( .A1(n676), .A2(n413), .ZN(n412) );
  INV_X1 U449 ( .A(KEYINPUT86), .ZN(n413) );
  XNOR2_X1 U450 ( .A(n655), .B(KEYINPUT91), .ZN(n485) );
  XNOR2_X1 U451 ( .A(G101), .B(G113), .ZN(n568) );
  XNOR2_X1 U452 ( .A(n607), .B(n606), .ZN(n658) );
  OR2_X1 U453 ( .A1(n607), .A2(n470), .ZN(n401) );
  INV_X1 U454 ( .A(KEYINPUT30), .ZN(n457) );
  XNOR2_X1 U455 ( .A(n591), .B(n590), .ZN(n592) );
  INV_X1 U456 ( .A(KEYINPUT81), .ZN(n590) );
  XNOR2_X1 U457 ( .A(n578), .B(KEYINPUT28), .ZN(n491) );
  NOR2_X1 U458 ( .A1(n608), .A2(n607), .ZN(n578) );
  XNOR2_X1 U459 ( .A(n543), .B(KEYINPUT104), .ZN(n544) );
  NOR2_X1 U460 ( .A1(G902), .A2(n752), .ZN(n545) );
  XNOR2_X1 U461 ( .A(G119), .B(G137), .ZN(n518) );
  XNOR2_X1 U462 ( .A(KEYINPUT96), .B(KEYINPUT72), .ZN(n510) );
  XOR2_X1 U463 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n511) );
  XNOR2_X1 U464 ( .A(G107), .B(KEYINPUT101), .ZN(n534) );
  XOR2_X1 U465 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n535) );
  XNOR2_X1 U466 ( .A(n529), .B(n527), .ZN(n475) );
  XNOR2_X1 U467 ( .A(G113), .B(G122), .ZN(n521) );
  AND2_X1 U468 ( .A1(n411), .A2(n408), .ZN(n404) );
  NAND2_X1 U469 ( .A1(n589), .A2(KEYINPUT86), .ZN(n408) );
  INV_X1 U470 ( .A(KEYINPUT64), .ZN(n507) );
  XNOR2_X1 U471 ( .A(n628), .B(n445), .ZN(n444) );
  INV_X1 U472 ( .A(KEYINPUT43), .ZN(n445) );
  NOR2_X1 U473 ( .A1(n663), .A2(n627), .ZN(n628) );
  XNOR2_X1 U474 ( .A(n494), .B(n493), .ZN(n631) );
  INV_X1 U475 ( .A(KEYINPUT39), .ZN(n493) );
  NOR2_X1 U476 ( .A1(n620), .A2(n621), .ZN(n494) );
  BUF_X1 U477 ( .A(n602), .Z(n629) );
  INV_X1 U478 ( .A(KEYINPUT0), .ZN(n462) );
  INV_X1 U479 ( .A(KEYINPUT89), .ZN(n660) );
  OR2_X1 U480 ( .A1(n563), .A2(G902), .ZN(n434) );
  INV_X1 U481 ( .A(KEYINPUT25), .ZN(n488) );
  XNOR2_X1 U482 ( .A(n388), .B(n496), .ZN(n678) );
  XNOR2_X1 U483 ( .A(n497), .B(n577), .ZN(n496) );
  INV_X1 U484 ( .A(n580), .ZN(n497) );
  XNOR2_X1 U485 ( .A(n460), .B(n461), .ZN(n468) );
  XNOR2_X1 U486 ( .A(n549), .B(G146), .ZN(n460) );
  OR2_X1 U487 ( .A1(G237), .A2(G902), .ZN(n594) );
  NOR2_X1 U488 ( .A1(n432), .A2(n619), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n430), .B(n625), .ZN(n429) );
  INV_X1 U490 ( .A(KEYINPUT48), .ZN(n465) );
  XOR2_X1 U491 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n522) );
  INV_X1 U492 ( .A(n412), .ZN(n409) );
  NAND2_X1 U493 ( .A1(n390), .A2(n389), .ZN(n626) );
  NAND2_X1 U494 ( .A1(n391), .A2(n371), .ZN(n390) );
  XNOR2_X1 U495 ( .A(n569), .B(n570), .ZN(n580) );
  XNOR2_X1 U496 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U497 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n573) );
  INV_X1 U498 ( .A(G107), .ZN(n492) );
  XNOR2_X1 U499 ( .A(n453), .B(n548), .ZN(n549) );
  XOR2_X1 U500 ( .A(G101), .B(G140), .Z(n548) );
  XNOR2_X1 U501 ( .A(n547), .B(n454), .ZN(n453) );
  INV_X1 U502 ( .A(KEYINPUT77), .ZN(n454) );
  XNOR2_X1 U503 ( .A(n580), .B(n449), .ZN(n760) );
  XNOR2_X1 U504 ( .A(n581), .B(n579), .ZN(n449) );
  INV_X1 U505 ( .A(KEYINPUT16), .ZN(n579) );
  NAND2_X1 U506 ( .A1(G234), .A2(G237), .ZN(n558) );
  NAND2_X1 U507 ( .A1(n366), .A2(n400), .ZN(n620) );
  XNOR2_X1 U508 ( .A(n401), .B(n457), .ZN(n400) );
  NAND2_X1 U509 ( .A1(n425), .A2(n491), .ZN(n600) );
  NOR2_X1 U510 ( .A1(n466), .A2(n426), .ZN(n425) );
  INV_X1 U511 ( .A(n490), .ZN(n426) );
  XNOR2_X1 U512 ( .A(n520), .B(n516), .ZN(n446) );
  XNOR2_X1 U513 ( .A(n448), .B(n767), .ZN(n447) );
  XNOR2_X1 U514 ( .A(n542), .B(n540), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n581), .B(n537), .ZN(n538) );
  XNOR2_X1 U516 ( .A(n528), .B(n475), .ZN(n531) );
  INV_X1 U517 ( .A(KEYINPUT112), .ZN(n441) );
  NAND2_X1 U518 ( .A1(n444), .A2(n443), .ZN(n442) );
  INV_X1 U519 ( .A(n364), .ZN(n443) );
  INV_X1 U520 ( .A(n659), .ZN(n499) );
  INV_X1 U521 ( .A(KEYINPUT31), .ZN(n666) );
  INV_X1 U522 ( .A(n600), .ZN(n690) );
  NOR2_X1 U523 ( .A1(n718), .A2(n714), .ZN(n480) );
  INV_X1 U524 ( .A(KEYINPUT109), .ZN(n482) );
  AND2_X1 U525 ( .A1(n662), .A2(n456), .ZN(n664) );
  NOR2_X1 U526 ( .A1(n663), .A2(n648), .ZN(n456) );
  NAND2_X1 U527 ( .A1(n505), .A2(n504), .ZN(n503) );
  XNOR2_X1 U528 ( .A(n506), .B(n377), .ZN(n505) );
  XNOR2_X1 U529 ( .A(n744), .B(n476), .ZN(n746) );
  AND2_X1 U530 ( .A1(n604), .A2(n603), .ZN(n366) );
  NOR2_X1 U531 ( .A1(n710), .A2(n419), .ZN(n367) );
  NOR2_X1 U532 ( .A1(n601), .A2(n424), .ZN(n368) );
  XOR2_X1 U533 ( .A(n565), .B(n488), .Z(n370) );
  AND2_X1 U534 ( .A1(n469), .A2(n610), .ZN(n371) );
  XNOR2_X1 U535 ( .A(G137), .B(n551), .ZN(n372) );
  INV_X1 U536 ( .A(n489), .ZN(n466) );
  AND2_X1 U537 ( .A1(n469), .A2(KEYINPUT110), .ZN(n373) );
  AND2_X1 U538 ( .A1(n491), .A2(n490), .ZN(n374) );
  NOR2_X1 U539 ( .A1(n724), .A2(n437), .ZN(n375) );
  XNOR2_X1 U540 ( .A(KEYINPUT93), .B(KEYINPUT33), .ZN(n376) );
  NAND2_X1 U541 ( .A1(G214), .A2(n594), .ZN(n700) );
  INV_X1 U542 ( .A(n700), .ZN(n470) );
  XOR2_X1 U543 ( .A(n678), .B(KEYINPUT62), .Z(n377) );
  XOR2_X1 U544 ( .A(G902), .B(KEYINPUT15), .Z(n589) );
  XOR2_X1 U545 ( .A(n563), .B(KEYINPUT122), .Z(n378) );
  XOR2_X1 U546 ( .A(n507), .B(KEYINPUT45), .Z(n379) );
  XNOR2_X1 U547 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n380) );
  NOR2_X1 U548 ( .A1(G952), .A2(n365), .ZN(n754) );
  INV_X1 U549 ( .A(n754), .ZN(n504) );
  BUF_X1 U550 ( .A(n712), .Z(n477) );
  XNOR2_X1 U551 ( .A(n657), .B(n656), .ZN(n665) );
  XNOR2_X1 U552 ( .A(n677), .B(n378), .ZN(n472) );
  NAND2_X1 U553 ( .A1(n472), .A2(n504), .ZN(n467) );
  NAND2_X1 U554 ( .A1(n439), .A2(n374), .ZN(n399) );
  NOR2_X1 U555 ( .A1(n650), .A2(n649), .ZN(n381) );
  XNOR2_X2 U556 ( .A(n382), .B(n379), .ZN(n755) );
  NAND2_X1 U557 ( .A1(n384), .A2(n383), .ZN(n382) );
  NAND2_X1 U558 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U559 ( .A1(n674), .A2(n675), .ZN(n385) );
  NAND2_X1 U560 ( .A1(n484), .A2(n780), .ZN(n386) );
  NAND2_X1 U561 ( .A1(n685), .A2(n779), .ZN(n654) );
  AND2_X2 U562 ( .A1(n755), .A2(n770), .ZN(n729) );
  XNOR2_X1 U563 ( .A(n388), .B(n767), .ZN(n768) );
  NAND2_X1 U564 ( .A1(n609), .A2(n373), .ZN(n389) );
  INV_X1 U565 ( .A(n609), .ZN(n391) );
  NAND2_X1 U566 ( .A1(n614), .A2(n663), .ZN(n393) );
  XNOR2_X1 U567 ( .A(n550), .B(n394), .ZN(n552) );
  INV_X1 U568 ( .A(KEYINPUT4), .ZN(n394) );
  NAND2_X1 U569 ( .A1(n395), .A2(n403), .ZN(n749) );
  AND2_X1 U570 ( .A1(n402), .A2(G475), .ZN(n395) );
  NAND2_X1 U571 ( .A1(n396), .A2(n403), .ZN(n742) );
  AND2_X1 U572 ( .A1(n402), .A2(G210), .ZN(n396) );
  NAND2_X1 U573 ( .A1(n397), .A2(G217), .ZN(n677) );
  NAND2_X1 U574 ( .A1(n397), .A2(G472), .ZN(n506) );
  NAND2_X1 U575 ( .A1(n397), .A2(G478), .ZN(n751) );
  NAND2_X1 U576 ( .A1(n397), .A2(G469), .ZN(n744) );
  NAND2_X1 U577 ( .A1(n788), .A2(n787), .ZN(n430) );
  NAND2_X1 U578 ( .A1(n631), .A2(n692), .ZN(n398) );
  XNOR2_X1 U579 ( .A(n624), .B(n440), .ZN(n439) );
  INV_X1 U580 ( .A(n607), .ZN(n718) );
  NAND2_X1 U581 ( .A1(n407), .A2(n755), .ZN(n405) );
  NAND2_X1 U582 ( .A1(n410), .A2(n409), .ZN(n406) );
  INV_X1 U583 ( .A(n755), .ZN(n410) );
  NAND2_X1 U584 ( .A1(n438), .A2(n418), .ZN(n502) );
  XNOR2_X2 U585 ( .A(n416), .B(n536), .ZN(n582) );
  XNOR2_X2 U586 ( .A(G143), .B(G128), .ZN(n416) );
  XNOR2_X2 U587 ( .A(n761), .B(KEYINPUT73), .ZN(n421) );
  XNOR2_X2 U588 ( .A(n417), .B(n492), .ZN(n761) );
  XNOR2_X2 U589 ( .A(G110), .B(G104), .ZN(n417) );
  INV_X1 U590 ( .A(n420), .ZN(n418) );
  INV_X1 U591 ( .A(n438), .ZN(n419) );
  NOR2_X2 U592 ( .A1(n420), .A2(n474), .ZN(n647) );
  NOR2_X1 U593 ( .A1(n420), .A2(n711), .ZN(n670) );
  NOR2_X1 U594 ( .A1(n721), .A2(n420), .ZN(n667) );
  XNOR2_X2 U595 ( .A(n463), .B(n462), .ZN(n420) );
  XNOR2_X1 U596 ( .A(n421), .B(KEYINPUT78), .ZN(n461) );
  NAND2_X1 U597 ( .A1(n689), .A2(n598), .ZN(n424) );
  NAND2_X1 U598 ( .A1(n600), .A2(KEYINPUT82), .ZN(n427) );
  NAND2_X1 U599 ( .A1(n597), .A2(n427), .ZN(n464) );
  NAND2_X1 U600 ( .A1(n431), .A2(n429), .ZN(n428) );
  NAND2_X1 U601 ( .A1(n648), .A2(n603), .ZN(n433) );
  NAND2_X1 U602 ( .A1(n435), .A2(KEYINPUT82), .ZN(n617) );
  INV_X1 U603 ( .A(n439), .ZN(n437) );
  AND2_X1 U604 ( .A1(n439), .A2(n438), .ZN(n698) );
  INV_X1 U605 ( .A(KEYINPUT41), .ZN(n440) );
  INV_X1 U606 ( .A(n782), .ZN(n630) );
  AND2_X1 U607 ( .A1(n541), .A2(G221), .ZN(n448) );
  XNOR2_X1 U608 ( .A(n596), .B(n595), .ZN(n644) );
  INV_X1 U609 ( .A(n455), .ZN(n528) );
  XNOR2_X1 U610 ( .A(n551), .B(n526), .ZN(n455) );
  XNOR2_X1 U611 ( .A(n483), .B(n482), .ZN(n481) );
  XNOR2_X1 U612 ( .A(n471), .B(KEYINPUT113), .ZN(n705) );
  XNOR2_X1 U613 ( .A(n458), .B(KEYINPUT107), .ZN(n474) );
  NOR2_X1 U614 ( .A1(n704), .A2(n645), .ZN(n458) );
  NOR2_X2 U615 ( .A1(n644), .A2(n643), .ZN(n463) );
  INV_X1 U616 ( .A(n780), .ZN(n674) );
  XNOR2_X2 U617 ( .A(n473), .B(n380), .ZN(n780) );
  NAND2_X1 U618 ( .A1(n464), .A2(KEYINPUT47), .ZN(n599) );
  XNOR2_X1 U619 ( .A(n515), .B(n514), .ZN(n541) );
  XNOR2_X1 U620 ( .A(n668), .B(KEYINPUT1), .ZN(n712) );
  XNOR2_X1 U621 ( .A(n467), .B(KEYINPUT123), .ZN(G66) );
  XNOR2_X2 U622 ( .A(n647), .B(n646), .ZN(n650) );
  NOR2_X1 U623 ( .A1(n611), .A2(n470), .ZN(n469) );
  NOR2_X1 U624 ( .A1(n621), .A2(n470), .ZN(n471) );
  NAND2_X1 U625 ( .A1(n500), .A2(n499), .ZN(n473) );
  XNOR2_X1 U626 ( .A(n498), .B(n745), .ZN(n476) );
  XNOR2_X1 U627 ( .A(n478), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U628 ( .A1(n750), .A2(n754), .ZN(n478) );
  XNOR2_X1 U629 ( .A(n479), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U630 ( .A1(n743), .A2(n754), .ZN(n479) );
  NAND2_X1 U631 ( .A1(n481), .A2(n480), .ZN(n685) );
  XNOR2_X1 U632 ( .A(n654), .B(n485), .ZN(n484) );
  INV_X1 U633 ( .A(n644), .ZN(n489) );
  INV_X1 U634 ( .A(n668), .ZN(n490) );
  INV_X1 U635 ( .A(n621), .ZN(n701) );
  NOR2_X1 U636 ( .A1(n705), .A2(n704), .ZN(n624) );
  XNOR2_X1 U637 ( .A(n502), .B(n501), .ZN(n500) );
  INV_X1 U638 ( .A(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U639 ( .A(n503), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U640 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U641 ( .A(n550), .B(n538), .ZN(n539) );
  XNOR2_X1 U642 ( .A(n593), .B(n592), .ZN(n602) );
  XNOR2_X1 U643 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n509) );
  XNOR2_X1 U644 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U645 ( .A(n574), .B(G116), .ZN(n575) );
  INV_X1 U646 ( .A(KEYINPUT65), .ZN(n536) );
  XNOR2_X1 U647 ( .A(n576), .B(n575), .ZN(n577) );
  INV_X1 U648 ( .A(KEYINPUT84), .ZN(n512) );
  INV_X1 U649 ( .A(KEYINPUT74), .ZN(n656) );
  INV_X1 U650 ( .A(n658), .ZN(n649) );
  XNOR2_X1 U651 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U652 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n652) );
  XNOR2_X1 U653 ( .A(n511), .B(n510), .ZN(n516) );
  NAND2_X1 U654 ( .A1(G234), .A2(n771), .ZN(n513) );
  XOR2_X1 U655 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n514) );
  XNOR2_X1 U656 ( .A(n584), .B(G140), .ZN(n517) );
  XOR2_X1 U657 ( .A(G110), .B(G128), .Z(n519) );
  XNOR2_X1 U658 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U659 ( .A(n522), .B(n521), .ZN(n529) );
  XNOR2_X1 U660 ( .A(G131), .B(KEYINPUT69), .ZN(n523) );
  XNOR2_X1 U661 ( .A(n523), .B(KEYINPUT68), .ZN(n551) );
  XOR2_X1 U662 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n525) );
  XNOR2_X1 U663 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U664 ( .A1(G214), .A2(n571), .ZN(n527) );
  INV_X1 U665 ( .A(n767), .ZN(n530) );
  XNOR2_X1 U666 ( .A(n531), .B(n530), .ZN(n747) );
  NOR2_X1 U667 ( .A1(G902), .A2(n747), .ZN(n533) );
  XNOR2_X1 U668 ( .A(KEYINPUT13), .B(G475), .ZN(n532) );
  XNOR2_X1 U669 ( .A(n535), .B(n534), .ZN(n540) );
  XOR2_X1 U670 ( .A(G116), .B(G122), .Z(n581) );
  XOR2_X1 U671 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n537) );
  INV_X1 U672 ( .A(G478), .ZN(n543) );
  INV_X1 U673 ( .A(n622), .ZN(n546) );
  NAND2_X1 U674 ( .A1(n623), .A2(n546), .ZN(n611) );
  INV_X1 U675 ( .A(n611), .ZN(n692) );
  NOR2_X1 U676 ( .A1(n623), .A2(n546), .ZN(n694) );
  NOR2_X1 U677 ( .A1(n692), .A2(n694), .ZN(n706) );
  INV_X1 U678 ( .A(n706), .ZN(n616) );
  OR2_X1 U679 ( .A1(KEYINPUT83), .A2(n616), .ZN(n597) );
  NAND2_X1 U680 ( .A1(G227), .A2(n771), .ZN(n547) );
  NAND2_X1 U681 ( .A1(n552), .A2(n372), .ZN(n553) );
  XNOR2_X2 U682 ( .A(n555), .B(G469), .ZN(n668) );
  NAND2_X1 U683 ( .A1(G952), .A2(n365), .ZN(n634) );
  INV_X1 U684 ( .A(n634), .ZN(n557) );
  NAND2_X1 U685 ( .A1(G953), .A2(G902), .ZN(n632) );
  NOR2_X1 U686 ( .A1(G900), .A2(n632), .ZN(n556) );
  NOR2_X1 U687 ( .A1(n557), .A2(n556), .ZN(n562) );
  XNOR2_X1 U688 ( .A(n558), .B(KEYINPUT14), .ZN(n699) );
  INV_X1 U689 ( .A(n589), .ZN(n676) );
  NAND2_X1 U690 ( .A1(n676), .A2(G234), .ZN(n559) );
  XNOR2_X1 U691 ( .A(n559), .B(KEYINPUT20), .ZN(n564) );
  NAND2_X1 U692 ( .A1(G221), .A2(n564), .ZN(n560) );
  XNOR2_X1 U693 ( .A(KEYINPUT21), .B(n560), .ZN(n645) );
  INV_X1 U694 ( .A(n645), .ZN(n715) );
  NAND2_X1 U695 ( .A1(n699), .A2(n715), .ZN(n561) );
  NOR2_X1 U696 ( .A1(n562), .A2(n561), .ZN(n603) );
  NAND2_X1 U697 ( .A1(n564), .A2(G217), .ZN(n565) );
  XNOR2_X1 U698 ( .A(n566), .B(KEYINPUT94), .ZN(n570) );
  INV_X1 U699 ( .A(KEYINPUT3), .ZN(n567) );
  NAND2_X1 U700 ( .A1(n571), .A2(G210), .ZN(n572) );
  XNOR2_X1 U701 ( .A(n573), .B(n572), .ZN(n576) );
  XOR2_X1 U702 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n583) );
  XOR2_X1 U703 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n587) );
  NAND2_X1 U704 ( .A1(G224), .A2(n771), .ZN(n586) );
  XNOR2_X1 U705 ( .A(n587), .B(n586), .ZN(n588) );
  NOR2_X1 U706 ( .A1(n740), .A2(n589), .ZN(n593) );
  NAND2_X1 U707 ( .A1(G210), .A2(n594), .ZN(n591) );
  NAND2_X1 U708 ( .A1(n602), .A2(n700), .ZN(n596) );
  XOR2_X1 U709 ( .A(KEYINPUT76), .B(KEYINPUT19), .Z(n595) );
  NAND2_X1 U710 ( .A1(n616), .A2(KEYINPUT83), .ZN(n598) );
  NOR2_X1 U711 ( .A1(KEYINPUT82), .A2(n600), .ZN(n601) );
  NOR2_X1 U712 ( .A1(n648), .A2(n668), .ZN(n604) );
  NAND2_X1 U713 ( .A1(n623), .A2(n622), .ZN(n659) );
  NOR2_X1 U714 ( .A1(n620), .A2(n659), .ZN(n605) );
  NAND2_X1 U715 ( .A1(n364), .A2(n605), .ZN(n689) );
  INV_X1 U716 ( .A(KEYINPUT114), .ZN(n615) );
  INV_X1 U717 ( .A(n477), .ZN(n663) );
  XNOR2_X1 U718 ( .A(KEYINPUT6), .B(KEYINPUT105), .ZN(n606) );
  INV_X1 U719 ( .A(KEYINPUT110), .ZN(n610) );
  NAND2_X1 U720 ( .A1(n626), .A2(n364), .ZN(n613) );
  XOR2_X1 U721 ( .A(KEYINPUT92), .B(KEYINPUT36), .Z(n612) );
  XNOR2_X1 U722 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X1 U723 ( .A1(KEYINPUT83), .A2(n617), .ZN(n618) );
  NOR2_X1 U724 ( .A1(KEYINPUT47), .A2(n618), .ZN(n619) );
  XOR2_X1 U725 ( .A(KEYINPUT46), .B(KEYINPUT88), .Z(n625) );
  XNOR2_X1 U726 ( .A(KEYINPUT111), .B(n626), .ZN(n627) );
  NAND2_X1 U727 ( .A1(n694), .A2(n631), .ZN(n697) );
  OR2_X1 U728 ( .A1(n632), .A2(G898), .ZN(n633) );
  NAND2_X1 U729 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U730 ( .A1(n635), .A2(n699), .ZN(n637) );
  INV_X1 U731 ( .A(KEYINPUT95), .ZN(n636) );
  NAND2_X1 U732 ( .A1(n637), .A2(n636), .ZN(n642) );
  INV_X1 U733 ( .A(G902), .ZN(n639) );
  NOR2_X1 U734 ( .A1(G898), .A2(n365), .ZN(n763) );
  NAND2_X1 U735 ( .A1(n763), .A2(KEYINPUT95), .ZN(n638) );
  NOR2_X1 U736 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U737 ( .A1(n640), .A2(n699), .ZN(n641) );
  NAND2_X1 U738 ( .A1(n642), .A2(n641), .ZN(n643) );
  INV_X1 U739 ( .A(KEYINPUT22), .ZN(n646) );
  NOR2_X1 U740 ( .A1(n714), .A2(n477), .ZN(n651) );
  INV_X1 U741 ( .A(KEYINPUT44), .ZN(n675) );
  NAND2_X1 U742 ( .A1(n675), .A2(KEYINPUT90), .ZN(n655) );
  NAND2_X1 U743 ( .A1(n714), .A2(n715), .ZN(n711) );
  NOR2_X1 U744 ( .A1(n712), .A2(n711), .ZN(n657) );
  XNOR2_X1 U745 ( .A(n381), .B(n660), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n667), .B(n666), .ZN(n695) );
  NOR2_X1 U747 ( .A1(n426), .A2(n718), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U749 ( .A(KEYINPUT97), .B(n671), .ZN(n681) );
  NOR2_X1 U750 ( .A1(n695), .A2(n681), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n672), .B(KEYINPUT98), .ZN(n673) );
  XOR2_X1 U752 ( .A(G104), .B(KEYINPUT115), .Z(n680) );
  NAND2_X1 U753 ( .A1(n681), .A2(n692), .ZN(n679) );
  XNOR2_X1 U754 ( .A(n680), .B(n679), .ZN(G6) );
  XOR2_X1 U755 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n683) );
  NAND2_X1 U756 ( .A1(n681), .A2(n694), .ZN(n682) );
  XNOR2_X1 U757 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U758 ( .A(G107), .B(n684), .ZN(G9) );
  XNOR2_X1 U759 ( .A(G110), .B(KEYINPUT116), .ZN(n686) );
  XNOR2_X1 U760 ( .A(n686), .B(n685), .ZN(G12) );
  XOR2_X1 U761 ( .A(G128), .B(KEYINPUT29), .Z(n688) );
  NAND2_X1 U762 ( .A1(n690), .A2(n694), .ZN(n687) );
  XNOR2_X1 U763 ( .A(n688), .B(n687), .ZN(G30) );
  XNOR2_X1 U764 ( .A(G143), .B(n689), .ZN(G45) );
  NAND2_X1 U765 ( .A1(n690), .A2(n692), .ZN(n691) );
  XNOR2_X1 U766 ( .A(n691), .B(G146), .ZN(G48) );
  NAND2_X1 U767 ( .A1(n695), .A2(n692), .ZN(n693) );
  XNOR2_X1 U768 ( .A(n693), .B(G113), .ZN(G15) );
  NAND2_X1 U769 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U770 ( .A(n696), .B(G116), .ZN(G18) );
  XNOR2_X1 U771 ( .A(G134), .B(n697), .ZN(G36) );
  NOR2_X1 U772 ( .A1(G953), .A2(n698), .ZN(n737) );
  NAND2_X1 U773 ( .A1(G952), .A2(n699), .ZN(n727) );
  NOR2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U775 ( .A(KEYINPUT119), .B(n702), .Z(n703) );
  NOR2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n709) );
  NOR2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U778 ( .A(n707), .B(KEYINPUT120), .ZN(n708) );
  NOR2_X1 U779 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U780 ( .A1(n477), .A2(n711), .ZN(n713) );
  XNOR2_X1 U781 ( .A(n713), .B(KEYINPUT50), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U783 ( .A(KEYINPUT49), .B(n716), .Z(n717) );
  NOR2_X1 U784 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U787 ( .A(KEYINPUT51), .B(n723), .ZN(n724) );
  NOR2_X1 U788 ( .A1(n367), .A2(n375), .ZN(n725) );
  XNOR2_X1 U789 ( .A(n725), .B(KEYINPUT52), .ZN(n726) );
  NOR2_X1 U790 ( .A1(n727), .A2(n726), .ZN(n735) );
  NOR2_X1 U791 ( .A1(KEYINPUT2), .A2(n770), .ZN(n728) );
  XNOR2_X1 U792 ( .A(n728), .B(KEYINPUT85), .ZN(n731) );
  NAND2_X1 U793 ( .A1(KEYINPUT2), .A2(n729), .ZN(n730) );
  NAND2_X1 U794 ( .A1(n731), .A2(n730), .ZN(n733) );
  NOR2_X1 U795 ( .A1(n755), .A2(KEYINPUT2), .ZN(n732) );
  NOR2_X1 U796 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U797 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U798 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U799 ( .A(KEYINPUT53), .B(n738), .Z(G75) );
  XOR2_X1 U800 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n739) );
  XNOR2_X1 U801 ( .A(n740), .B(n739), .ZN(n741) );
  XOR2_X1 U802 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n745) );
  NOR2_X1 U803 ( .A1(n754), .A2(n746), .ZN(G54) );
  XNOR2_X1 U804 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U805 ( .A1(n754), .A2(n753), .ZN(G63) );
  NAND2_X1 U806 ( .A1(n365), .A2(n755), .ZN(n759) );
  NAND2_X1 U807 ( .A1(G953), .A2(G224), .ZN(n756) );
  XNOR2_X1 U808 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U809 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U810 ( .A1(n759), .A2(n758), .ZN(n765) );
  XOR2_X1 U811 ( .A(n761), .B(n760), .Z(n762) );
  NOR2_X1 U812 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U813 ( .A(n765), .B(n764), .ZN(n766) );
  XNOR2_X1 U814 ( .A(KEYINPUT124), .B(n766), .ZN(G69) );
  XOR2_X1 U815 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n769) );
  XNOR2_X1 U816 ( .A(n769), .B(n768), .ZN(n773) );
  XOR2_X1 U817 ( .A(n770), .B(n773), .Z(n772) );
  NAND2_X1 U818 ( .A1(n772), .A2(n365), .ZN(n777) );
  XNOR2_X1 U819 ( .A(G227), .B(n773), .ZN(n774) );
  NAND2_X1 U820 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U821 ( .A1(n775), .A2(G953), .ZN(n776) );
  NAND2_X1 U822 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U823 ( .A(G119), .B(KEYINPUT127), .Z(n778) );
  XNOR2_X1 U824 ( .A(n779), .B(n778), .ZN(G21) );
  XNOR2_X1 U825 ( .A(n780), .B(G122), .ZN(G24) );
  XOR2_X1 U826 ( .A(G140), .B(KEYINPUT118), .Z(n781) );
  XNOR2_X1 U827 ( .A(n782), .B(n781), .ZN(G42) );
  XOR2_X1 U828 ( .A(G101), .B(n783), .Z(G3) );
  XOR2_X1 U829 ( .A(KEYINPUT117), .B(KEYINPUT37), .Z(n784) );
  XNOR2_X1 U830 ( .A(n785), .B(n784), .ZN(n786) );
  XNOR2_X1 U831 ( .A(G125), .B(n786), .ZN(G27) );
  XNOR2_X1 U832 ( .A(G131), .B(n787), .ZN(G33) );
  XNOR2_X1 U833 ( .A(n788), .B(G137), .ZN(G39) );
endmodule

