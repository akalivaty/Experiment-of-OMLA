//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT69), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT64), .A3(G134), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n192), .B1(new_n190), .B2(G134), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G137), .ZN(new_n195));
  OAI211_X1 g009(.A(G131), .B(new_n191), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n199), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n205), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT11), .B1(new_n190), .B2(G134), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n190), .A2(G134), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n190), .A2(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n194), .A2(G137), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(new_n192), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n219), .A2(KEYINPUT65), .A3(G131), .A4(new_n191), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n198), .A2(new_n210), .A3(new_n216), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  OAI22_X1  g038(.A1(new_n201), .A2(new_n203), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n222), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n214), .B1(new_n213), .B2(new_n215), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n194), .B2(G137), .ZN(new_n231));
  AND4_X1   g045(.A1(new_n214), .A2(new_n231), .A3(new_n215), .A4(new_n218), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n228), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G116), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT2), .B(G113), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n221), .A2(new_n233), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n221), .A2(new_n233), .A3(new_n241), .A4(KEYINPUT66), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n221), .A2(new_n233), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n221), .A2(new_n233), .A3(KEYINPUT30), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n240), .A3(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(G101), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n246), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT31), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n241), .B1(new_n247), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT68), .B1(new_n221), .B2(new_n233), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n244), .A2(new_n245), .B1(new_n240), .B2(new_n247), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n261), .ZN(new_n267));
  INV_X1    g081(.A(new_n256), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n260), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n246), .A2(new_n251), .A3(new_n271), .A4(new_n256), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n259), .B1(new_n258), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n189), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n258), .A2(new_n272), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n258), .A2(new_n259), .B1(new_n267), .B2(new_n268), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT32), .A3(new_n189), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n265), .B(new_n256), .C1(new_n266), .C2(new_n261), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n246), .A2(new_n251), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n268), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n282), .A2(new_n283), .ZN(new_n289));
  OAI21_X1  g103(.A(G472), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n276), .A2(new_n281), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G217), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(G234), .B2(new_n287), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n295));
  XNOR2_X1  g109(.A(G125), .B(G140), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n202), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n300), .A2(KEYINPUT16), .A3(G140), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n296), .A2(KEYINPUT16), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT16), .ZN(new_n304));
  INV_X1    g118(.A(G140), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G125), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(G146), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n199), .A2(G119), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT23), .ZN(new_n311));
  INV_X1    g125(.A(G110), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n199), .A2(G119), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n311), .B(new_n312), .C1(new_n315), .C2(new_n310), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT24), .B(G110), .Z(new_n318));
  OR2_X1    g132(.A1(new_n309), .A2(KEYINPUT70), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n309), .B1(new_n313), .B2(KEYINPUT70), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n299), .B(new_n308), .C1(new_n317), .C2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n311), .B1(new_n315), .B2(new_n310), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G110), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n296), .A2(KEYINPUT16), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n301), .A2(new_n302), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n307), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(new_n202), .ZN(new_n328));
  AOI21_X1  g142(.A(G146), .B1(new_n303), .B2(new_n307), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n319), .A2(new_n320), .A3(new_n318), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT71), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n319), .A2(new_n320), .A3(new_n333), .A4(new_n318), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n295), .B(new_n322), .C1(new_n330), .C2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G137), .ZN(new_n337));
  INV_X1    g151(.A(G953), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n338), .A2(G221), .A3(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n337), .B(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n327), .A2(new_n202), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n308), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n343), .A2(new_n324), .A3(new_n332), .A4(new_n334), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n295), .B1(new_n344), .B2(new_n322), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n295), .B(new_n340), .C1(new_n344), .C2(new_n322), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n287), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(new_n322), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT74), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(new_n336), .A3(new_n340), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n341), .A2(new_n345), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n287), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n294), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n293), .A2(G902), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n291), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G221), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT9), .B(G234), .Z(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(new_n366), .B2(new_n287), .ZN(new_n367));
  XOR2_X1   g181(.A(new_n367), .B(KEYINPUT76), .Z(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n370));
  AOI21_X1  g184(.A(G128), .B1(new_n206), .B2(new_n207), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n207), .A2(new_n208), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n205), .B(KEYINPUT78), .C1(new_n226), .C2(G128), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n209), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT77), .A3(G104), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(G101), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G107), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n382), .A2(new_n376), .A3(KEYINPUT77), .A4(G104), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n379), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n381), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n380), .A2(G107), .ZN(new_n386));
  OAI21_X1  g200(.A(G101), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n375), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n229), .A2(new_n232), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G101), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n396), .A3(G101), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n228), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n388), .A2(KEYINPUT10), .A3(new_n210), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n391), .A2(new_n392), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G110), .B(G140), .ZN(new_n401));
  INV_X1    g215(.A(G227), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G953), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n401), .B(new_n403), .Z(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n384), .A2(new_n387), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n371), .A2(new_n372), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n209), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n389), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n392), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT12), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT12), .ZN(new_n414));
  AOI211_X1 g228(.A(new_n414), .B(new_n392), .C1(new_n389), .C2(new_n410), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n400), .A2(KEYINPUT79), .A3(new_n404), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n391), .A2(new_n398), .A3(new_n399), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n412), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n404), .B1(new_n420), .B2(new_n400), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G469), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n287), .ZN(new_n425));
  INV_X1    g239(.A(new_n404), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n400), .B1(new_n413), .B2(new_n415), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n400), .A2(new_n404), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n426), .A2(new_n427), .B1(new_n428), .B2(new_n420), .ZN(new_n429));
  OAI21_X1  g243(.A(G469), .B1(new_n429), .B2(G902), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n369), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n299), .B1(new_n202), .B2(new_n296), .ZN(new_n432));
  INV_X1    g246(.A(G237), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n338), .A3(G214), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n200), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n252), .A2(G143), .A3(G214), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(KEYINPUT18), .A2(G131), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(G131), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT17), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n435), .A2(new_n214), .A3(new_n436), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n437), .A2(KEYINPUT17), .A3(G131), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n444), .A2(new_n342), .A3(new_n308), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G113), .B(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT84), .B(G104), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n448), .B(new_n449), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n440), .A2(new_n450), .A3(new_n446), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G475), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n441), .A2(new_n443), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT19), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n297), .B2(new_n298), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n296), .A2(new_n459), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n308), .B(new_n458), .C1(new_n462), .C2(G146), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n450), .B1(new_n463), .B2(new_n440), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n455), .A4(new_n287), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n455), .B(new_n287), .C1(new_n457), .C2(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT20), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n456), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G952), .ZN(new_n471));
  AOI211_X1 g285(.A(G953), .B(new_n471), .C1(G234), .C2(G237), .ZN(new_n472));
  XOR2_X1   g286(.A(KEYINPUT21), .B(G898), .Z(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI211_X1 g288(.A(new_n287), .B(new_n338), .C1(G234), .C2(G237), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n366), .A2(G217), .A3(new_n338), .ZN(new_n478));
  INV_X1    g292(.A(G122), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(G116), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n236), .A2(G122), .ZN(new_n481));
  OAI21_X1  g295(.A(G107), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n236), .A2(G122), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(G116), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n376), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n482), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n482), .B2(new_n486), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT87), .B1(new_n200), .B2(G128), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n199), .A3(G143), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT13), .ZN(new_n494));
  OAI211_X1 g308(.A(KEYINPUT86), .B(new_n494), .C1(new_n199), .C2(G143), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n200), .A2(G128), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT86), .B1(new_n497), .B2(new_n494), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n493), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n200), .A2(KEYINPUT13), .A3(G128), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G134), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(new_n194), .A3(new_n497), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n493), .A2(KEYINPUT89), .A3(new_n194), .A4(new_n497), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n489), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT90), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n236), .B2(G122), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n512), .B2(new_n481), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT90), .B(new_n485), .C1(new_n480), .C2(new_n511), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(new_n514), .C1(KEYINPUT14), .C2(new_n484), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G107), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n493), .A2(new_n497), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G134), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n504), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n519), .A3(new_n486), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n509), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n521), .B1(new_n509), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n478), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n509), .A2(new_n520), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT91), .ZN(new_n526));
  INV_X1    g340(.A(new_n478), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n509), .A2(new_n520), .A3(new_n521), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(G902), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G478), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n530), .B1(KEYINPUT15), .B2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n522), .A2(new_n523), .A3(new_n478), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n287), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n531), .A2(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n431), .A2(new_n470), .A3(new_n477), .A4(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT83), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT80), .B1(new_n235), .B2(KEYINPUT5), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n235), .A2(new_n237), .A3(KEYINPUT5), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT80), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT5), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n234), .A4(G116), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n542), .A2(new_n543), .A3(G113), .A4(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n238), .A2(new_n239), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n408), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT81), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n547), .A2(new_n548), .A3(new_n387), .A4(new_n384), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n388), .A2(KEYINPUT81), .A3(new_n548), .A4(new_n547), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G122), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(G125), .B1(new_n409), .B2(new_n209), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n300), .B1(new_n225), .B2(new_n227), .ZN(new_n559));
  OAI211_X1 g373(.A(G224), .B(new_n338), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n338), .A2(G224), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n210), .A2(new_n300), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n395), .A2(new_n240), .A3(new_n397), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n552), .A3(new_n555), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n561), .A2(new_n563), .A3(new_n565), .A4(new_n562), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n557), .A2(new_n567), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n571), .A2(new_n287), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n552), .ZN(new_n573));
  INV_X1    g387(.A(new_n555), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT6), .A3(new_n569), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n560), .A2(new_n564), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT6), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(new_n578), .A3(new_n574), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G210), .B1(G237), .B2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT82), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n572), .A2(new_n580), .A3(new_n582), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n572), .A2(new_n580), .A3(KEYINPUT82), .A4(new_n582), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G214), .B1(G237), .B2(G902), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n541), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n587), .A2(KEYINPUT83), .A3(new_n590), .A4(new_n588), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n540), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n291), .A2(KEYINPUT75), .A3(new_n361), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n364), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT92), .B(G101), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G3));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  OAI22_X1  g413(.A1(new_n533), .A2(new_n534), .B1(KEYINPUT94), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT94), .B(KEYINPUT33), .Z(new_n601));
  NAND3_X1  g415(.A1(new_n524), .A2(new_n529), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n600), .A2(G478), .A3(new_n287), .A4(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n535), .B2(new_n531), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n530), .A2(KEYINPUT95), .A3(G478), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n470), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n582), .B1(new_n572), .B2(new_n580), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n591), .B1(new_n609), .B2(KEYINPUT93), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT93), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n584), .A2(new_n611), .A3(new_n586), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n607), .A2(new_n608), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT96), .B1(new_n613), .B2(new_n476), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n581), .A2(KEYINPUT93), .A3(new_n583), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n586), .A2(new_n611), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n590), .B(new_n615), .C1(new_n616), .C2(new_n609), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n535), .A2(new_n604), .A3(new_n531), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT95), .B1(new_n530), .B2(G478), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n470), .B1(new_n621), .B2(new_n603), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n618), .A2(new_n622), .A3(new_n623), .A4(new_n477), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n614), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n278), .B2(new_n279), .ZN(new_n626));
  INV_X1    g440(.A(G472), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n274), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT25), .B1(new_n355), .B2(new_n287), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n349), .B(G902), .C1(new_n353), .C2(new_n354), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n293), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n359), .ZN(new_n632));
  AOI211_X1 g446(.A(G469), .B(G902), .C1(new_n418), .C2(new_n422), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n427), .A2(new_n426), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n428), .A2(new_n420), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n424), .B1(new_n636), .B2(new_n287), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n368), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n628), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n625), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  NAND2_X1  g456(.A1(new_n456), .A2(KEYINPUT97), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n454), .B2(new_n455), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n467), .A2(new_n469), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n647), .A3(new_n477), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n617), .A2(new_n648), .A3(new_n539), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n639), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  INV_X1    g466(.A(new_n628), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n340), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n351), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n358), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT98), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n655), .A2(new_n658), .A3(new_n358), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n631), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n594), .A2(new_n653), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  NOR2_X1   g478(.A1(new_n638), .A2(new_n617), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n472), .B1(new_n475), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n646), .A2(new_n647), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n291), .A2(new_n665), .A3(new_n538), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n657), .A2(new_n659), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n357), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n199), .ZN(G30));
  XOR2_X1   g488(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n667), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n431), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT40), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n589), .B(KEYINPUT38), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n661), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n608), .A2(new_n538), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT32), .B1(new_n280), .B2(new_n189), .ZN(new_n684));
  AOI211_X1 g498(.A(new_n275), .B(new_n188), .C1(new_n278), .C2(new_n279), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n284), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n268), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n266), .A2(new_n268), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n287), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n683), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n590), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n679), .B1(new_n682), .B2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n681), .A2(KEYINPUT99), .A3(new_n590), .A4(new_n692), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n678), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT101), .B(G143), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G45));
  AOI211_X1 g512(.A(new_n667), .B(new_n470), .C1(new_n621), .C2(new_n603), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n291), .A2(new_n665), .A3(new_n699), .A4(new_n661), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  AND3_X1   g515(.A1(new_n400), .A2(KEYINPUT79), .A3(new_n404), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT79), .B1(new_n400), .B2(new_n404), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n413), .A2(new_n415), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n287), .B1(new_n705), .B2(new_n421), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(KEYINPUT102), .A3(new_n425), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n706), .A2(new_n709), .A3(G469), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n367), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n711), .A2(new_n291), .A3(new_n361), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n625), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT41), .B(G113), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND4_X1  g529(.A1(new_n711), .A2(new_n649), .A3(new_n291), .A4(new_n361), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NOR3_X1   g531(.A1(new_n608), .A2(new_n538), .A3(new_n476), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n291), .A2(new_n718), .A3(new_n661), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n367), .B(new_n617), .C1(new_n708), .C2(new_n710), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  OAI21_X1  g536(.A(KEYINPUT104), .B1(new_n626), .B2(new_n627), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n267), .A2(new_n268), .B1(KEYINPUT31), .B2(new_n257), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n272), .B1(new_n724), .B2(new_n725), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n189), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n287), .B1(new_n270), .B2(new_n273), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(G472), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n723), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n357), .A2(new_n733), .A3(new_n360), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT105), .B1(new_n631), .B2(new_n359), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n608), .A2(new_n612), .A3(new_n538), .A4(new_n610), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n476), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n732), .A2(new_n711), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  NAND3_X1  g554(.A1(new_n711), .A2(new_n618), .A3(new_n699), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n723), .A2(new_n731), .A3(new_n728), .A4(new_n661), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n743), .A2(KEYINPUT106), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(KEYINPUT106), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT107), .B(G125), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G27));
  NAND2_X1  g562(.A1(new_n736), .A2(new_n291), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n591), .B1(new_n587), .B2(new_n588), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n367), .B1(new_n425), .B2(new_n430), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n699), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT42), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n362), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n622), .A2(new_n668), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(KEYINPUT42), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n755), .A2(new_n752), .A3(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  NAND4_X1  g574(.A1(new_n755), .A2(new_n538), .A3(new_n669), .A4(new_n752), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND2_X1  g576(.A1(new_n628), .A2(new_n661), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT108), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n607), .A2(new_n470), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(KEYINPUT43), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n607), .B2(new_n470), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n750), .B(KEYINPUT109), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n769), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n636), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n429), .A2(KEYINPUT45), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(G469), .ZN(new_n780));
  NAND2_X1  g594(.A1(G469), .A2(G902), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n781), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n425), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n367), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n676), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n776), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n425), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT46), .B1(new_n780), .B2(new_n781), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n786), .B2(new_n787), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n797), .B2(new_n794), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n686), .A2(new_n290), .A3(new_n632), .A4(new_n750), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n798), .A2(new_n756), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n305), .ZN(G42));
  NAND2_X1  g615(.A1(new_n361), .A2(KEYINPUT105), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n733), .B1(new_n357), .B2(new_n360), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n804), .A2(new_n591), .A3(new_n369), .A4(new_n765), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n686), .A2(new_n691), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n708), .A2(new_n710), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT49), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n805), .A2(new_n680), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n739), .A2(new_n716), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n625), .A2(new_n712), .B1(new_n719), .B2(new_n720), .ZN(new_n811));
  INV_X1    g625(.A(new_n753), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n744), .B2(new_n745), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n291), .A2(new_n669), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n672), .A2(new_n638), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(new_n539), .A3(new_n750), .A4(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n754), .A2(new_n761), .A3(new_n758), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n622), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n608), .B2(new_n539), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n592), .A2(new_n593), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n822), .A3(new_n477), .A4(new_n639), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n596), .A2(new_n662), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT111), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n596), .A2(new_n662), .A3(new_n826), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n700), .B1(new_n670), .B2(new_n672), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n743), .B(KEYINPUT106), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(new_n742), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n787), .B(new_n668), .C1(new_n633), .C2(new_n637), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(new_n661), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n672), .A2(new_n751), .A3(KEYINPUT113), .A4(new_n668), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n692), .A3(new_n618), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n831), .A2(new_n832), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n829), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n746), .A3(new_n838), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT52), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n819), .A2(new_n828), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n832), .B1(new_n831), .B2(new_n838), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n832), .A2(new_n840), .A3(new_n746), .A4(new_n838), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n828), .A4(new_n819), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n845), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT115), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n845), .A2(new_n849), .A3(new_n853), .A4(new_n850), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n819), .A2(new_n828), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n848), .B1(new_n856), .B2(KEYINPUT112), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(KEYINPUT112), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT53), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT114), .B1(new_n843), .B2(new_n844), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n819), .A2(new_n828), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT53), .A4(new_n848), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n855), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n861), .A2(new_n864), .ZN(new_n869));
  INV_X1    g683(.A(new_n859), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n844), .B1(new_n870), .B2(new_n857), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n850), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n852), .A2(new_n854), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT116), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n807), .A2(new_n369), .ZN(new_n875));
  INV_X1    g689(.A(new_n795), .ZN(new_n876));
  INV_X1    g690(.A(new_n796), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n794), .B1(new_n793), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n875), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n472), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n766), .A2(new_n880), .A3(new_n768), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n723), .A2(new_n728), .A3(new_n731), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n804), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n879), .A2(new_n774), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n711), .A2(new_n750), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n711), .A2(KEYINPUT117), .A3(new_n750), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n830), .A3(new_n881), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n591), .A2(new_n881), .A3(new_n883), .A4(new_n680), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT50), .B1(new_n892), .B2(new_n711), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n881), .A2(new_n883), .A3(new_n591), .A4(new_n680), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT50), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n807), .A2(new_n787), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n885), .B(new_n891), .C1(new_n893), .C2(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n888), .A2(new_n806), .A3(new_n889), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n632), .A2(new_n880), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n621), .A2(new_n470), .A3(new_n603), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n899), .A2(new_n900), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n888), .A2(new_n806), .A3(new_n889), .A4(new_n901), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT118), .B1(new_n905), .B2(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT51), .B1(new_n898), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n892), .A2(KEYINPUT50), .A3(new_n711), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n773), .B1(new_n798), .B2(new_n875), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n910), .A2(new_n911), .B1(new_n912), .B2(new_n884), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n907), .A4(new_n891), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n890), .A2(new_n291), .A3(new_n736), .A4(new_n881), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT48), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n899), .A2(new_n622), .A3(new_n901), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n471), .B(G953), .C1(new_n884), .C2(new_n720), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT119), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n868), .A2(new_n874), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(G952), .A2(G953), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n809), .B1(new_n923), .B2(new_n924), .ZN(G75));
  NAND2_X1  g739(.A1(new_n845), .A2(new_n849), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(G210), .A3(G902), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n576), .A2(new_n579), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(new_n577), .Z(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n338), .A2(G952), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n932), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n927), .A2(new_n928), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT120), .ZN(G51));
  XNOR2_X1  g753(.A(new_n781), .B(KEYINPUT121), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT57), .ZN(new_n941));
  INV_X1    g755(.A(new_n926), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n850), .ZN(new_n943));
  INV_X1    g757(.A(new_n851), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n423), .B(KEYINPUT122), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n942), .A2(new_n287), .A3(new_n780), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n934), .B1(new_n947), .B2(new_n948), .ZN(G54));
  NAND4_X1  g763(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n950));
  INV_X1    g764(.A(new_n465), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(new_n934), .ZN(G60));
  NAND2_X1  g768(.A1(new_n600), .A2(new_n602), .ZN(new_n955));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT59), .Z(new_n957));
  NOR2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n943), .B2(new_n944), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n935), .ZN(new_n960));
  INV_X1    g774(.A(new_n957), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n867), .B1(new_n855), .B2(new_n866), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT116), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n964), .B2(new_n955), .ZN(G63));
  XNOR2_X1  g779(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n292), .A2(new_n287), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n926), .A2(new_n655), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n935), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n355), .B1(new_n926), .B2(new_n968), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g787(.A(G224), .ZN(new_n974));
  OAI21_X1  g788(.A(G953), .B1(new_n474), .B2(new_n974), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n828), .A2(new_n810), .A3(new_n811), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n930), .B1(G898), .B2(new_n338), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G69));
  NAND2_X1  g793(.A1(new_n249), .A2(new_n250), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(new_n462), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  INV_X1    g797(.A(new_n831), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n696), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n696), .B2(new_n984), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n800), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n364), .A2(new_n595), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n677), .B1(new_n821), .B2(KEYINPUT124), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n821), .A2(KEYINPUT124), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n989), .A2(new_n750), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n789), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(KEYINPUT125), .B(new_n982), .C1(new_n994), .C2(G953), .ZN(new_n995));
  NAND2_X1  g809(.A1(G900), .A2(G953), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n776), .B1(new_n737), .B2(new_n749), .ZN(new_n997));
  INV_X1    g811(.A(new_n788), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n984), .A2(new_n800), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n999), .A2(new_n759), .A3(new_n761), .A4(new_n1000), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n981), .B(new_n996), .C1(new_n1001), .C2(G953), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT125), .ZN(new_n1003));
  AOI21_X1  g817(.A(G953), .B1(new_n987), .B2(new_n993), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n981), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n995), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(G953), .B1(new_n402), .B2(new_n666), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1008), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1010), .A2(new_n1011), .ZN(G72));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  INV_X1    g828(.A(new_n976), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1014), .B1(new_n1001), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n687), .A3(new_n268), .ZN(new_n1017));
  INV_X1    g831(.A(new_n688), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n987), .A2(new_n976), .A3(new_n993), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(new_n1014), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n935), .B(new_n1017), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g838(.A1(new_n869), .A2(new_n871), .B1(new_n257), .B2(new_n285), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1014), .B2(new_n1025), .ZN(G57));
endmodule


