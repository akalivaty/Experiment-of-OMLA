//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT71), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT71), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n193), .B2(G122), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(G122), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n187), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT71), .B(G116), .ZN(new_n197));
  INV_X1    g011(.A(G122), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n193), .A2(new_n188), .A3(G122), .ZN(new_n200));
  INV_X1    g014(.A(new_n195), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT93), .A4(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(new_n202), .A3(G107), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(G134), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n205), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n214), .B(new_n201), .C1(new_n197), .C2(new_n198), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT13), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n205), .B1(new_n207), .B2(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n219), .B(KEYINPUT91), .C1(new_n218), .C2(new_n205), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n220), .B(G134), .C1(KEYINPUT91), .C2(new_n219), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n201), .B1(new_n197), .B2(new_n198), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n215), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n212), .B(KEYINPUT92), .Z(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT9), .B(G234), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n228), .B(KEYINPUT84), .ZN(new_n229));
  INV_X1    g043(.A(G953), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(G217), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n217), .A2(new_n226), .A3(new_n231), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G478), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n233), .A2(new_n236), .A3(new_n234), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n237), .A3(G478), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT94), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G237), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n230), .A3(G214), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n246), .B(G143), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT18), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XOR2_X1   g064(.A(G125), .B(G140), .Z(new_n251));
  OR2_X1    g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n246), .B(new_n204), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G131), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n250), .B(new_n254), .C1(new_n248), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n247), .A2(new_n249), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n260), .A2(KEYINPUT16), .A3(G140), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT16), .ZN(new_n263));
  OAI211_X1 g077(.A(G146), .B(new_n262), .C1(new_n251), .C2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n251), .B(KEYINPUT19), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G146), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n257), .B1(new_n259), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G113), .B(G122), .ZN(new_n268));
  INV_X1    g082(.A(G104), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT17), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n256), .A2(new_n258), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G146), .ZN(new_n275));
  INV_X1    g089(.A(G140), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n260), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(G125), .A2(G140), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n263), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n275), .B1(new_n279), .B2(new_n261), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n255), .A2(KEYINPUT17), .A3(G131), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n274), .A2(new_n264), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n270), .B(KEYINPUT90), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n257), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n272), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G475), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n236), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT20), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n284), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n270), .B1(new_n282), .B2(new_n257), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n236), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G475), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n285), .A2(KEYINPUT20), .A3(new_n286), .A4(new_n236), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n289), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n230), .A2(G952), .ZN(new_n297));
  NAND2_X1  g111(.A1(G234), .A2(G237), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT21), .B(G898), .Z(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(G902), .A3(G953), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n244), .A2(KEYINPUT95), .A3(new_n296), .A4(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n242), .A2(new_n243), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT94), .B1(new_n239), .B2(new_n241), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n296), .B(new_n302), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT95), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(G110), .B(G122), .Z(new_n312));
  INV_X1    g126(.A(G119), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n197), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(KEYINPUT70), .A2(G119), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT70), .A2(G119), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n189), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT69), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT2), .B(G113), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT70), .B(G119), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G116), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n313), .B2(new_n197), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT69), .A3(new_n320), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT3), .B1(new_n269), .B2(G107), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(new_n214), .A3(G104), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G101), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n269), .A2(G107), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n332), .A2(KEYINPUT85), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n329), .A2(new_n331), .A3(new_n333), .A4(new_n334), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n329), .A2(new_n331), .A3(new_n334), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G101), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n328), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT4), .B1(new_n340), .B2(G101), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n327), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT88), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n324), .B(KEYINPUT5), .C1(new_n313), .C2(new_n197), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n346), .B(G113), .C1(KEYINPUT5), .C2(new_n324), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n214), .A2(G104), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n334), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n335), .A2(new_n338), .B1(G101), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n325), .A2(new_n320), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n344), .A2(new_n345), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n345), .B1(new_n344), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n312), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT89), .ZN(new_n357));
  INV_X1    g171(.A(new_n312), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n344), .A2(new_n358), .A3(new_n352), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT6), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n356), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n336), .A2(new_n337), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n336), .A2(new_n337), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n341), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n343), .B1(new_n365), .B2(KEYINPUT4), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n322), .A2(new_n326), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n352), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT88), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n358), .B1(new_n369), .B2(new_n353), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT89), .B1(new_n370), .B2(new_n360), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n275), .A2(G143), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n204), .A2(G146), .ZN(new_n375));
  NOR2_X1   g189(.A1(KEYINPUT0), .A2(G128), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n374), .A2(new_n375), .B1(new_n376), .B2(KEYINPUT64), .ZN(new_n377));
  OR2_X1    g191(.A1(KEYINPUT0), .A2(G128), .ZN(new_n378));
  AND2_X1   g192(.A1(KEYINPUT0), .A2(G128), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT64), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT65), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(KEYINPUT65), .A3(new_n381), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(new_n375), .A3(new_n379), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT66), .ZN(new_n387));
  XNOR2_X1  g201(.A(G143), .B(G146), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT66), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n379), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n384), .A2(new_n385), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G125), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n393));
  OAI22_X1  g207(.A1(new_n393), .A2(new_n375), .B1(new_n210), .B2(G146), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT68), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n374), .A2(new_n375), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT1), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G128), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n395), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n388), .A2(KEYINPUT68), .A3(new_n393), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n394), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n392), .B1(G125), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n230), .A2(G224), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n362), .A2(new_n371), .A3(new_n373), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n402), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n347), .A2(new_n351), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(new_n350), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n312), .B(KEYINPUT8), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n407), .B(new_n359), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(new_n236), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G210), .B1(G237), .B2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n405), .A2(new_n414), .A3(new_n412), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n311), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G221), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n229), .B2(new_n236), .ZN(new_n420));
  INV_X1    g234(.A(G469), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n394), .A2(KEYINPUT86), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n399), .A2(new_n400), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n394), .A2(KEYINPUT86), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n350), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT10), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n401), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n426), .A2(new_n427), .B1(new_n428), .B2(new_n350), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n391), .B1(new_n342), .B2(new_n343), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT11), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n211), .B2(G137), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n211), .A2(G137), .ZN(new_n433));
  INV_X1    g247(.A(G137), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(KEYINPUT11), .A3(G134), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G131), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n432), .A2(new_n435), .A3(new_n249), .A4(new_n433), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n429), .A2(new_n430), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G140), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n230), .A2(G227), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n442), .B(new_n443), .Z(new_n444));
  AND2_X1   g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT12), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n349), .A2(G101), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n363), .B2(new_n364), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n401), .ZN(new_n449));
  AOI211_X1 g263(.A(new_n446), .B(new_n440), .C1(new_n426), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n426), .A2(new_n449), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT12), .B1(new_n451), .B2(new_n439), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n445), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT87), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT87), .B1(new_n429), .B2(new_n430), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n439), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n444), .B1(new_n457), .B2(new_n441), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n421), .B(new_n236), .C1(new_n454), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n444), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n441), .B1(new_n452), .B2(new_n450), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n457), .A2(new_n445), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G469), .B1(new_n462), .B2(G902), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n420), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n309), .A2(new_n418), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT32), .ZN(new_n466));
  NOR2_X1   g280(.A1(G472), .A2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT76), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n387), .A2(new_n390), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n377), .A2(KEYINPUT65), .A3(new_n381), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT65), .B1(new_n377), .B2(new_n381), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n439), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n394), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT68), .B1(new_n388), .B2(new_n393), .ZN(new_n475));
  AND4_X1   g289(.A1(KEYINPUT68), .A2(new_n393), .A3(new_n374), .A4(new_n375), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n434), .A2(G134), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n211), .A2(G137), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n438), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n473), .A2(new_n483), .A3(new_n322), .A4(new_n326), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n438), .A2(new_n480), .A3(KEYINPUT67), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n477), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n488), .A2(new_n473), .B1(new_n322), .B2(new_n326), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n484), .B1(new_n489), .B2(KEYINPUT75), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n473), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n491), .A2(KEYINPUT75), .A3(new_n327), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT28), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n484), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT73), .B(KEYINPUT27), .Z(new_n497));
  NAND3_X1  g311(.A1(new_n245), .A2(new_n230), .A3(G210), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT26), .B(G101), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n499), .B(new_n500), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n469), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  AOI211_X1 g317(.A(KEYINPUT76), .B(new_n501), .C1(new_n493), .C2(new_n495), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT31), .ZN(new_n506));
  INV_X1    g320(.A(new_n484), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n473), .A2(KEYINPUT30), .A3(new_n483), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT72), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n473), .A2(new_n483), .A3(KEYINPUT72), .A4(KEYINPUT30), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n367), .B1(new_n491), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n507), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n506), .B1(new_n515), .B2(new_n501), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n514), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n517), .A2(new_n506), .A3(new_n484), .A4(new_n501), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT74), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n515), .A2(KEYINPUT74), .A3(new_n506), .A4(new_n501), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n468), .B1(new_n505), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT77), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n466), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n520), .A2(new_n521), .ZN(new_n526));
  INV_X1    g340(.A(new_n516), .ZN(new_n527));
  INV_X1    g341(.A(new_n495), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n491), .A2(new_n327), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n489), .A2(KEYINPUT75), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n484), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n528), .B1(new_n533), .B2(KEYINPUT28), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT76), .B1(new_n534), .B2(new_n501), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n496), .A2(new_n469), .A3(new_n502), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n526), .A2(new_n527), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n467), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT77), .A3(KEYINPUT32), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n525), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n484), .A2(KEYINPUT78), .A3(new_n494), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT78), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n495), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n473), .A2(new_n483), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n327), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n484), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n541), .B(new_n543), .C1(new_n547), .C2(new_n494), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT29), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n501), .C1(KEYINPUT29), .C2(new_n496), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n515), .A2(new_n502), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n550), .B(new_n236), .C1(KEYINPUT29), .C2(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n552), .A2(G472), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n540), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(G137), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n230), .A2(G221), .A3(G234), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT82), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT80), .ZN(new_n561));
  INV_X1    g375(.A(new_n317), .ZN(new_n562));
  NOR4_X1   g376(.A1(new_n562), .A2(new_n315), .A3(KEYINPUT23), .A4(G128), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n313), .A2(G128), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n323), .B2(G128), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n563), .B1(new_n565), .B2(KEYINPUT23), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT79), .B1(new_n566), .B2(G110), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT24), .B(G110), .Z(new_n568));
  OR2_X1    g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G128), .B1(new_n562), .B2(new_n315), .ZN(new_n570));
  INV_X1    g384(.A(new_n564), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(KEYINPUT23), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT23), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n316), .A2(new_n573), .A3(new_n209), .A4(new_n317), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT79), .ZN(new_n576));
  INV_X1    g390(.A(G110), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n567), .A2(new_n569), .A3(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n264), .A2(new_n252), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n264), .A2(new_n280), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n572), .A2(G110), .A3(new_n574), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n565), .A2(new_n568), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n561), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  AOI211_X1 g401(.A(KEYINPUT80), .B(new_n585), .C1(new_n579), .C2(new_n580), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n560), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n581), .A2(new_n586), .A3(new_n559), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n236), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT25), .ZN(new_n592));
  INV_X1    g406(.A(G217), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(G234), .B2(new_n236), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n589), .A2(new_n595), .A3(new_n236), .A4(new_n590), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n592), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n589), .A2(new_n590), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n594), .A2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT83), .B1(new_n555), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n553), .B1(new_n525), .B2(new_n539), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT83), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n604), .A2(new_n605), .A3(new_n601), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n465), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  NAND2_X1  g422(.A1(new_n537), .A2(new_n236), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n523), .B1(new_n609), .B2(G472), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n464), .A3(new_n602), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n405), .A2(new_n414), .A3(new_n412), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n414), .B1(new_n405), .B2(new_n412), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n310), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n302), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n235), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n231), .A2(KEYINPUT96), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n233), .A2(new_n234), .A3(new_n619), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n227), .A2(new_n619), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(KEYINPUT33), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(KEYINPUT97), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n625), .A2(G478), .A3(new_n236), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G478), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n240), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n295), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n615), .A2(new_n616), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n612), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n269), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n633), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(new_n244), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n418), .A2(new_n296), .A3(new_n637), .A4(new_n302), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n612), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n645));
  OR4_X1    g459(.A1(KEYINPUT36), .A2(new_n587), .A3(new_n588), .A4(new_n560), .ZN(new_n646));
  OAI22_X1  g460(.A1(new_n587), .A2(new_n588), .B1(KEYINPUT36), .B2(new_n560), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n599), .A3(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n597), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n645), .B1(new_n597), .B2(new_n648), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n644), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n597), .A2(new_n648), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT100), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n597), .A2(new_n645), .A3(new_n648), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(KEYINPUT101), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n309), .A2(new_n418), .A3(new_n610), .A4(new_n464), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n658), .B(new_n660), .ZN(G12));
  NAND2_X1  g475(.A1(new_n459), .A2(new_n463), .ZN(new_n662));
  INV_X1    g476(.A(new_n420), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n615), .B(new_n664), .C1(new_n651), .C2(new_n655), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n299), .B1(G900), .B2(new_n301), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n637), .A2(new_n296), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n604), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n209), .ZN(G30));
  OAI21_X1  g484(.A(KEYINPUT103), .B1(new_n613), .B2(new_n614), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT38), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n613), .A2(new_n614), .A3(KEYINPUT103), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n673), .B1(new_n672), .B2(new_n674), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n525), .A2(new_n539), .ZN(new_n679));
  INV_X1    g493(.A(G472), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n515), .A2(new_n502), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(G902), .B1(new_n547), .B2(new_n502), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n311), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n653), .A2(new_n654), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n244), .A2(new_n296), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n678), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n678), .A2(new_n686), .A3(new_n693), .A4(new_n690), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n666), .B(KEYINPUT39), .Z(new_n696));
  NOR2_X1   g510(.A1(new_n664), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n695), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT105), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  AOI21_X1  g517(.A(new_n664), .B1(new_n651), .B2(new_n655), .ZN(new_n704));
  INV_X1    g518(.A(new_n666), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n296), .B(new_n705), .C1(new_n627), .C2(new_n629), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n418), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n704), .A2(new_n555), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n604), .A2(new_n707), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n704), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  NOR2_X1   g529(.A1(new_n454), .A2(new_n458), .ZN(new_n716));
  OAI21_X1  g530(.A(G469), .B1(new_n716), .B2(G902), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n663), .A3(new_n459), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n555), .A2(new_n632), .A3(new_n602), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NOR3_X1   g536(.A1(new_n604), .A2(new_n601), .A3(new_n718), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n640), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NAND2_X1  g539(.A1(new_n651), .A2(new_n655), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n615), .A2(new_n718), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n555), .A2(new_n726), .A3(new_n309), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT107), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NAND2_X1  g544(.A1(new_n609), .A2(G472), .ZN(new_n731));
  AOI22_X1  g545(.A1(new_n546), .A2(KEYINPUT28), .B1(new_n495), .B2(new_n542), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n501), .B1(new_n732), .B2(new_n541), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n527), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT108), .B1(new_n516), .B2(new_n733), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n737), .A3(new_n526), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n467), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n731), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n601), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n302), .A3(new_n688), .A4(new_n727), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  AOI22_X1  g557(.A1(new_n609), .A2(G472), .B1(new_n467), .B2(new_n738), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n653), .A3(new_n706), .A4(new_n654), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n719), .A2(new_n418), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n260), .ZN(G27));
  XNOR2_X1  g562(.A(new_n523), .B(new_n466), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n601), .B1(new_n749), .B2(new_n554), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n664), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n613), .A2(new_n614), .A3(new_n311), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n464), .A2(KEYINPUT109), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n750), .A2(new_n755), .A3(new_n706), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n757));
  INV_X1    g571(.A(new_n706), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n604), .A2(new_n601), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n756), .A2(KEYINPUT42), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NAND3_X1  g576(.A1(new_n668), .A2(new_n602), .A3(new_n755), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  INV_X1    g578(.A(new_n753), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n630), .A2(new_n296), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n610), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(new_n653), .A4(new_n654), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n765), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n462), .A2(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n462), .A2(KEYINPUT45), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(G469), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(G469), .A2(G902), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT46), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n459), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n776), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n420), .A3(new_n696), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n772), .B(new_n782), .C1(new_n771), .C2(new_n770), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n781), .B2(new_n420), .ZN(new_n786));
  OAI211_X1 g600(.A(KEYINPUT47), .B(new_n663), .C1(new_n779), .C2(new_n780), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n758), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n604), .A3(new_n601), .A4(new_n753), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  OR2_X1    g604(.A1(new_n679), .A2(new_n684), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n601), .A2(new_n311), .A3(new_n420), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(KEYINPUT110), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n674), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT38), .B1(new_n795), .B2(new_n671), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n675), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n766), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n717), .A2(new_n459), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT49), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n794), .A2(new_n797), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n747), .B1(new_n665), .B2(new_n668), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n418), .A2(new_n688), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n652), .B2(new_n705), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n597), .A2(KEYINPUT112), .A3(new_n648), .A4(new_n666), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n664), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n791), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n711), .A2(new_n712), .A3(new_n704), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n712), .B1(new_n711), .B2(new_n704), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n803), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n714), .A2(KEYINPUT52), .A3(new_n803), .A4(new_n810), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n242), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n753), .A2(new_n818), .A3(new_n666), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n704), .A2(new_n819), .A3(new_n555), .A4(new_n296), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n740), .A2(new_n687), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n755), .A2(new_n706), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n763), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT111), .B1(new_n818), .B2(new_n295), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n296), .A2(new_n826), .A3(new_n242), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n631), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n418), .A3(new_n302), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n656), .A2(new_n657), .B1(new_n829), .B2(new_n611), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n555), .A2(KEYINPUT83), .A3(new_n602), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n605), .B1(new_n604), .B2(new_n601), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n830), .B1(new_n833), .B2(new_n465), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n824), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n728), .A2(new_n720), .A3(new_n742), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n761), .A2(new_n836), .A3(new_n724), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n817), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n817), .B2(new_n838), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT54), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n299), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n768), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n727), .A3(new_n741), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n839), .A2(new_n840), .ZN(new_n847));
  INV_X1    g661(.A(new_n830), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n607), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT113), .B1(new_n849), .B2(new_n823), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n824), .A2(new_n834), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n840), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n837), .B1(new_n815), .B2(new_n816), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n847), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(KEYINPUT50), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n797), .A2(new_n311), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n768), .A2(new_n741), .A3(new_n844), .A4(new_n719), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n861), .ZN(new_n863));
  INV_X1    g677(.A(new_n859), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n311), .A3(new_n797), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n768), .A2(new_n741), .A3(new_n844), .A4(new_n753), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n800), .A2(new_n420), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n786), .A2(new_n787), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n765), .A2(new_n718), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n685), .A2(new_n844), .A3(new_n602), .A4(new_n873), .ZN(new_n874));
  OR3_X1    g688(.A1(new_n874), .A2(new_n295), .A3(new_n630), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n845), .A2(new_n873), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n821), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n866), .A2(new_n872), .A3(new_n875), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n869), .A2(new_n871), .B1(new_n821), .B2(new_n876), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(KEYINPUT51), .A3(new_n875), .A4(new_n866), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n880), .A2(new_n297), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n843), .A2(new_n846), .A3(new_n857), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n874), .A2(new_n631), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n876), .A2(new_n750), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT48), .Z(new_n887));
  NOR3_X1   g701(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n802), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT116), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n892), .B(new_n802), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(G75));
  AOI21_X1  g708(.A(new_n236), .B1(new_n847), .B2(new_n855), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(G210), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n362), .A2(new_n371), .A3(new_n373), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n404), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n896), .A2(new_n899), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n230), .A2(G952), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G51));
  AND2_X1   g717(.A1(new_n853), .A2(new_n854), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT54), .B1(new_n904), .B2(new_n842), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(KEYINPUT117), .A3(new_n857), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT117), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n847), .A2(new_n855), .A3(new_n907), .A4(new_n856), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n776), .B(KEYINPUT57), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n716), .B(KEYINPUT118), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n895), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n775), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n917));
  INV_X1    g731(.A(new_n902), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n910), .B2(new_n911), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT119), .B1(new_n920), .B2(new_n902), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(G54));
  NAND3_X1  g736(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n923));
  INV_X1    g737(.A(new_n285), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n923), .A2(KEYINPUT120), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT120), .B1(new_n923), .B2(new_n924), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(G60));
  NAND2_X1  g742(.A1(new_n625), .A2(new_n626), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT59), .Z(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n906), .A2(new_n908), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n843), .A2(new_n857), .ZN(new_n936));
  INV_X1    g750(.A(new_n931), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n902), .B1(new_n938), .B2(new_n929), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n933), .A2(new_n934), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n935), .A2(new_n939), .A3(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n847), .B2(new_n855), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n646), .A3(new_n647), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n945), .B(new_n918), .C1(new_n598), .C2(new_n944), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT61), .Z(G66));
  NAND3_X1  g761(.A1(new_n834), .A2(new_n724), .A3(new_n836), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n230), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n230), .B1(new_n300), .B2(G224), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n897), .B1(G898), .B2(new_n230), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  NAND2_X1  g771(.A1(new_n491), .A2(new_n513), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n512), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT124), .Z(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n265), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(G900), .A2(G953), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n782), .A2(new_n750), .A3(new_n805), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n789), .A2(new_n783), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n714), .A2(new_n803), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n965), .A2(new_n761), .A3(new_n763), .A4(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n962), .B(new_n963), .C1(new_n967), .C2(G953), .ZN(new_n968));
  NAND2_X1  g782(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n789), .A2(new_n783), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n701), .A2(new_n966), .ZN(new_n971));
  NOR2_X1   g785(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n701), .B(new_n966), .C1(KEYINPUT125), .C2(KEYINPUT62), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n833), .A2(new_n697), .A3(new_n753), .A4(new_n828), .ZN(new_n976));
  AOI21_X1  g790(.A(G953), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n968), .B1(new_n977), .B2(new_n962), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n230), .B1(G227), .B2(G900), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT126), .Z(new_n981));
  OR3_X1    g795(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n978), .B2(new_n980), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n978), .A2(new_n981), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n975), .A2(new_n976), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(new_n948), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n902), .B1(new_n989), .B2(new_n681), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n987), .B1(new_n967), .B2(new_n948), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n515), .A3(new_n502), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n841), .A2(new_n842), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n993), .A2(new_n551), .A3(new_n682), .A4(new_n987), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n990), .A2(new_n992), .A3(new_n994), .ZN(G57));
endmodule


