

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791;

  AND2_X1 U383 ( .A1(n607), .A2(n606), .ZN(n733) );
  INV_X1 U384 ( .A(n720), .ZN(n717) );
  NAND2_X1 U385 ( .A1(n580), .A2(n581), .ZN(n720) );
  XNOR2_X1 U386 ( .A(n440), .B(n427), .ZN(n673) );
  XNOR2_X2 U387 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X2 U388 ( .A(n635), .B(KEYINPUT6), .ZN(n620) );
  XNOR2_X2 U389 ( .A(n429), .B(n428), .ZN(n635) );
  XNOR2_X2 U390 ( .A(n563), .B(G146), .ZN(n440) );
  AND2_X2 U391 ( .A1(n398), .A2(n397), .ZN(n366) );
  BUF_X2 U392 ( .A(n372), .Z(n692) );
  OR2_X1 U393 ( .A1(n566), .A2(n431), .ZN(n386) );
  INV_X2 U394 ( .A(G953), .ZN(n774) );
  AND2_X2 U395 ( .A1(n407), .A2(n406), .ZN(n405) );
  XNOR2_X2 U396 ( .A(n508), .B(n412), .ZN(n563) );
  AND2_X1 U397 ( .A1(n390), .A2(n389), .ZN(n388) );
  INV_X1 U398 ( .A(KEYINPUT35), .ZN(n375) );
  NAND2_X1 U399 ( .A1(n388), .A2(n391), .ZN(n414) );
  NOR2_X1 U400 ( .A1(n572), .A2(n791), .ZN(n573) );
  XNOR2_X1 U401 ( .A(n579), .B(KEYINPUT114), .ZN(n789) );
  AND2_X1 U402 ( .A1(n394), .A2(n627), .ZN(n390) );
  XNOR2_X1 U403 ( .A(n381), .B(n554), .ZN(n572) );
  NAND2_X1 U404 ( .A1(n392), .A2(n393), .ZN(n391) );
  XNOR2_X1 U405 ( .A(n541), .B(n540), .ZN(n624) );
  OR2_X1 U406 ( .A1(n570), .A2(n569), .ZN(n588) );
  AND2_X1 U407 ( .A1(n555), .A2(n615), .ZN(n376) );
  NAND2_X1 U408 ( .A1(n387), .A2(n364), .ZN(n541) );
  XNOR2_X1 U409 ( .A(n386), .B(n432), .ZN(n385) );
  OR2_X1 U410 ( .A1(n699), .A2(G902), .ZN(n441) );
  AND2_X1 U411 ( .A1(n556), .A2(n555), .ZN(n616) );
  NAND2_X1 U412 ( .A1(n556), .A2(n376), .ZN(n395) );
  INV_X1 U413 ( .A(n557), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n640), .B(KEYINPUT1), .ZN(n738) );
  NAND2_X1 U415 ( .A1(n405), .A2(n402), .ZN(n363) );
  NAND2_X1 U416 ( .A1(n405), .A2(n402), .ZN(n495) );
  XOR2_X1 U417 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n462) );
  XNOR2_X1 U418 ( .A(KEYINPUT72), .B(G131), .ZN(n518) );
  NAND2_X1 U419 ( .A1(n494), .A2(n659), .ZN(n406) );
  XNOR2_X1 U420 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n656) );
  XNOR2_X1 U421 ( .A(G101), .B(G116), .ZN(n422) );
  XNOR2_X1 U422 ( .A(n458), .B(KEYINPUT98), .ZN(n459) );
  INV_X1 U423 ( .A(KEYINPUT24), .ZN(n458) );
  XNOR2_X1 U424 ( .A(G119), .B(G137), .ZN(n455) );
  XOR2_X1 U425 ( .A(G110), .B(G128), .Z(n456) );
  XNOR2_X1 U426 ( .A(n503), .B(n502), .ZN(n506) );
  INV_X1 U427 ( .A(KEYINPUT7), .ZN(n502) );
  XNOR2_X1 U428 ( .A(n514), .B(n513), .ZN(n580) );
  XNOR2_X1 U429 ( .A(n512), .B(n511), .ZN(n513) );
  INV_X1 U430 ( .A(KEYINPUT104), .ZN(n511) );
  NOR2_X1 U431 ( .A1(G953), .A2(G237), .ZN(n523) );
  XOR2_X1 U432 ( .A(G104), .B(G143), .Z(n517) );
  XNOR2_X1 U433 ( .A(G113), .B(G122), .ZN(n519) );
  XNOR2_X1 U434 ( .A(n420), .B(n518), .ZN(n412) );
  INV_X1 U435 ( .A(G237), .ZN(n430) );
  NAND2_X1 U436 ( .A1(n754), .A2(n753), .ZN(n757) );
  NAND2_X1 U437 ( .A1(n404), .A2(n491), .ZN(n403) );
  XNOR2_X1 U438 ( .A(G119), .B(G113), .ZN(n425) );
  XNOR2_X1 U439 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n424) );
  XNOR2_X1 U440 ( .A(G104), .B(KEYINPUT93), .ZN(n434) );
  XNOR2_X1 U441 ( .A(G107), .B(G101), .ZN(n433) );
  NOR2_X1 U442 ( .A1(n729), .A2(KEYINPUT2), .ZN(n730) );
  XNOR2_X1 U443 ( .A(n411), .B(n409), .ZN(n752) );
  XNOR2_X1 U444 ( .A(n564), .B(n410), .ZN(n409) );
  NOR2_X1 U445 ( .A1(n757), .A2(n756), .ZN(n411) );
  INV_X1 U446 ( .A(KEYINPUT111), .ZN(n410) );
  BUF_X1 U447 ( .A(n635), .Z(n641) );
  XNOR2_X1 U448 ( .A(n472), .B(n471), .ZN(n619) );
  XNOR2_X1 U449 ( .A(n468), .B(KEYINPUT78), .ZN(n469) );
  XOR2_X1 U450 ( .A(KEYINPUT62), .B(n673), .Z(n674) );
  XNOR2_X1 U451 ( .A(n460), .B(n459), .ZN(n464) );
  INV_X1 U452 ( .A(G107), .ZN(n507) );
  XNOR2_X1 U453 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U454 ( .A1(n367), .A2(n717), .ZN(n381) );
  NAND2_X1 U455 ( .A1(n416), .A2(n387), .ZN(n589) );
  INV_X1 U456 ( .A(n588), .ZN(n416) );
  AND2_X1 U457 ( .A1(n539), .A2(n737), .ZN(n364) );
  XOR2_X1 U458 ( .A(n533), .B(n532), .Z(n365) );
  XOR2_X1 U459 ( .A(n500), .B(n499), .Z(n367) );
  AND2_X1 U460 ( .A1(n370), .A2(n631), .ZN(n368) );
  NAND2_X1 U461 ( .A1(n654), .A2(n653), .ZN(n369) );
  NAND2_X1 U462 ( .A1(n398), .A2(n397), .ZN(n370) );
  NAND2_X1 U463 ( .A1(n401), .A2(n732), .ZN(n371) );
  NAND2_X1 U464 ( .A1(n401), .A2(n732), .ZN(n399) );
  NAND2_X1 U465 ( .A1(n624), .A2(n543), .ZN(n415) );
  XNOR2_X2 U466 ( .A(n399), .B(KEYINPUT67), .ZN(n372) );
  XOR2_X1 U467 ( .A(G140), .B(KEYINPUT10), .Z(n454) );
  XNOR2_X1 U468 ( .A(n470), .B(n469), .ZN(n472) );
  NAND2_X1 U469 ( .A1(n396), .A2(n368), .ZN(n633) );
  BUF_X1 U470 ( .A(n632), .Z(n787) );
  INV_X1 U471 ( .A(n632), .ZN(n396) );
  INV_X1 U472 ( .A(n374), .ZN(n632) );
  XNOR2_X1 U473 ( .A(n614), .B(KEYINPUT107), .ZN(n615) );
  AND2_X2 U474 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X2 U475 ( .A1(n550), .A2(n565), .ZN(n574) );
  OR2_X1 U476 ( .A1(n560), .A2(n742), .ZN(n373) );
  XNOR2_X2 U477 ( .A(n414), .B(n375), .ZN(n374) );
  XNOR2_X2 U478 ( .A(n589), .B(KEYINPUT81), .ZN(n718) );
  OR2_X2 U479 ( .A1(n560), .A2(n742), .ZN(n648) );
  NAND2_X1 U480 ( .A1(n400), .A2(KEYINPUT2), .ZN(n732) );
  NAND2_X1 U481 ( .A1(n663), .A2(n380), .ZN(n377) );
  AND2_X2 U482 ( .A1(n377), .A2(n378), .ZN(n401) );
  OR2_X1 U483 ( .A1(n379), .A2(n418), .ZN(n378) );
  INV_X1 U484 ( .A(n662), .ZN(n379) );
  AND2_X1 U485 ( .A1(n658), .A2(n662), .ZN(n380) );
  INV_X1 U486 ( .A(n617), .ZN(n397) );
  XNOR2_X2 U487 ( .A(n395), .B(KEYINPUT32), .ZN(n398) );
  NAND2_X1 U488 ( .A1(n413), .A2(KEYINPUT34), .ZN(n394) );
  AND2_X1 U489 ( .A1(n385), .A2(n474), .ZN(n585) );
  NAND2_X1 U490 ( .A1(n385), .A2(n382), .ZN(n500) );
  NOR2_X1 U491 ( .A1(n384), .A2(n383), .ZN(n382) );
  INV_X1 U492 ( .A(n754), .ZN(n383) );
  INV_X1 U493 ( .A(n474), .ZN(n384) );
  XNOR2_X2 U494 ( .A(n575), .B(n365), .ZN(n387) );
  NAND2_X1 U495 ( .A1(n725), .A2(KEYINPUT34), .ZN(n389) );
  INV_X1 U496 ( .A(n725), .ZN(n392) );
  AND2_X1 U497 ( .A1(n637), .A2(n625), .ZN(n393) );
  INV_X1 U498 ( .A(n398), .ZN(n618) );
  XNOR2_X2 U499 ( .A(n408), .B(G134), .ZN(n508) );
  XNOR2_X1 U500 ( .A(n408), .B(n477), .ZN(n484) );
  NAND2_X1 U501 ( .A1(n495), .A2(n753), .ZN(n575) );
  XNOR2_X2 U502 ( .A(n371), .B(KEYINPUT67), .ZN(n696) );
  INV_X1 U503 ( .A(n663), .ZN(n400) );
  OR2_X1 U504 ( .A1(n679), .A2(n403), .ZN(n402) );
  INV_X1 U505 ( .A(n494), .ZN(n404) );
  NAND2_X1 U506 ( .A1(n679), .A2(n494), .ZN(n407) );
  XNOR2_X1 U507 ( .A(n490), .B(n489), .ZN(n679) );
  XNOR2_X2 U508 ( .A(n419), .B(G143), .ZN(n408) );
  INV_X1 U509 ( .A(n637), .ZN(n413) );
  XNOR2_X2 U510 ( .A(n415), .B(n544), .ZN(n556) );
  XNOR2_X1 U511 ( .A(n657), .B(n656), .ZN(n728) );
  NAND2_X1 U512 ( .A1(n728), .A2(n733), .ZN(n663) );
  OR2_X1 U513 ( .A1(G902), .A2(n666), .ZN(n417) );
  AND2_X1 U514 ( .A1(n659), .A2(KEYINPUT70), .ZN(n418) );
  INV_X1 U515 ( .A(KEYINPUT90), .ZN(n651) );
  INV_X1 U516 ( .A(KEYINPUT34), .ZN(n625) );
  INV_X1 U517 ( .A(n626), .ZN(n627) );
  INV_X1 U518 ( .A(KEYINPUT0), .ZN(n540) );
  XNOR2_X1 U519 ( .A(n506), .B(n505), .ZN(n510) );
  XNOR2_X2 U520 ( .A(G128), .B(KEYINPUT66), .ZN(n419) );
  XNOR2_X2 U521 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n475) );
  XNOR2_X1 U522 ( .A(n475), .B(G137), .ZN(n420) );
  NAND2_X1 U523 ( .A1(n523), .A2(G210), .ZN(n421) );
  XNOR2_X1 U524 ( .A(n421), .B(KEYINPUT5), .ZN(n423) );
  XNOR2_X1 U525 ( .A(n423), .B(n422), .ZN(n426) );
  XNOR2_X1 U526 ( .A(n425), .B(n424), .ZN(n486) );
  XNOR2_X1 U527 ( .A(n426), .B(n486), .ZN(n427) );
  OR2_X2 U528 ( .A1(n673), .A2(G902), .ZN(n429) );
  INV_X1 U529 ( .A(G472), .ZN(n428) );
  XNOR2_X1 U530 ( .A(n635), .B(KEYINPUT108), .ZN(n566) );
  INV_X1 U531 ( .A(G902), .ZN(n536) );
  NAND2_X1 U532 ( .A1(n536), .A2(n430), .ZN(n492) );
  NAND2_X1 U533 ( .A1(n492), .A2(G214), .ZN(n753) );
  INV_X1 U534 ( .A(n753), .ZN(n431) );
  INV_X1 U535 ( .A(KEYINPUT30), .ZN(n432) );
  XNOR2_X1 U536 ( .A(n433), .B(G110), .ZN(n435) );
  XNOR2_X1 U537 ( .A(n435), .B(n434), .ZN(n780) );
  XNOR2_X1 U538 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n436) );
  XNOR2_X1 U539 ( .A(n780), .B(n436), .ZN(n489) );
  NAND2_X1 U540 ( .A1(n774), .A2(G227), .ZN(n437) );
  XNOR2_X1 U541 ( .A(n437), .B(G140), .ZN(n438) );
  XNOR2_X1 U542 ( .A(n489), .B(n438), .ZN(n439) );
  XNOR2_X1 U543 ( .A(n440), .B(n439), .ZN(n699) );
  XNOR2_X2 U544 ( .A(n441), .B(G469), .ZN(n640) );
  XNOR2_X1 U545 ( .A(G902), .B(KEYINPUT15), .ZN(n491) );
  NAND2_X1 U546 ( .A1(n491), .A2(G234), .ZN(n442) );
  XNOR2_X1 U547 ( .A(n442), .B(KEYINPUT20), .ZN(n467) );
  AND2_X1 U548 ( .A1(n467), .A2(G221), .ZN(n444) );
  XNOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT21), .ZN(n443) );
  XNOR2_X1 U550 ( .A(n444), .B(n443), .ZN(n741) );
  NAND2_X1 U551 ( .A1(G237), .A2(G234), .ZN(n445) );
  XNOR2_X1 U552 ( .A(n445), .B(KEYINPUT14), .ZN(n737) );
  NAND2_X1 U553 ( .A1(G902), .A2(n737), .ZN(n446) );
  NOR2_X1 U554 ( .A1(G900), .A2(n446), .ZN(n447) );
  NAND2_X1 U555 ( .A1(G953), .A2(n447), .ZN(n448) );
  XNOR2_X1 U556 ( .A(n448), .B(KEYINPUT109), .ZN(n451) );
  NAND2_X1 U557 ( .A1(n774), .A2(G952), .ZN(n537) );
  INV_X1 U558 ( .A(n537), .ZN(n449) );
  AND2_X1 U559 ( .A1(n737), .A2(n449), .ZN(n450) );
  NOR2_X1 U560 ( .A1(n451), .A2(n450), .ZN(n452) );
  XNOR2_X1 U561 ( .A(n452), .B(KEYINPUT82), .ZN(n453) );
  NOR2_X1 U562 ( .A1(n741), .A2(n453), .ZN(n549) );
  XNOR2_X2 U563 ( .A(G146), .B(G125), .ZN(n476) );
  XNOR2_X1 U564 ( .A(n476), .B(n454), .ZN(n561) );
  XNOR2_X1 U565 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U566 ( .A(n561), .B(n457), .ZN(n466) );
  XNOR2_X1 U567 ( .A(KEYINPUT23), .B(KEYINPUT97), .ZN(n460) );
  NAND2_X1 U568 ( .A1(n774), .A2(G234), .ZN(n461) );
  XNOR2_X1 U569 ( .A(n462), .B(n461), .ZN(n501) );
  NAND2_X1 U570 ( .A1(G221), .A2(n501), .ZN(n463) );
  XNOR2_X1 U571 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U572 ( .A(n466), .B(n465), .ZN(n688) );
  NOR2_X1 U573 ( .A1(G902), .A2(n688), .ZN(n470) );
  NAND2_X1 U574 ( .A1(G217), .A2(n467), .ZN(n468) );
  INV_X1 U575 ( .A(KEYINPUT25), .ZN(n471) );
  INV_X1 U576 ( .A(n619), .ZN(n545) );
  AND2_X1 U577 ( .A1(n549), .A2(n545), .ZN(n473) );
  AND2_X1 U578 ( .A1(n640), .A2(n473), .ZN(n474) );
  XNOR2_X1 U579 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U580 ( .A1(n774), .A2(G224), .ZN(n478) );
  XNOR2_X1 U581 ( .A(n478), .B(KEYINPUT79), .ZN(n482) );
  XNOR2_X1 U582 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n480) );
  XNOR2_X1 U583 ( .A(KEYINPUT80), .B(KEYINPUT94), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U585 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U586 ( .A(n484), .B(n483), .ZN(n488) );
  INV_X1 U587 ( .A(G122), .ZN(n485) );
  XNOR2_X1 U588 ( .A(n485), .B(G116), .ZN(n504) );
  XNOR2_X1 U589 ( .A(n504), .B(KEYINPUT16), .ZN(n487) );
  XNOR2_X1 U590 ( .A(n487), .B(n486), .ZN(n781) );
  XNOR2_X1 U591 ( .A(n488), .B(n781), .ZN(n490) );
  INV_X1 U592 ( .A(n491), .ZN(n659) );
  NAND2_X1 U593 ( .A1(n492), .A2(G210), .ZN(n493) );
  XNOR2_X1 U594 ( .A(n493), .B(KEYINPUT95), .ZN(n494) );
  INV_X1 U595 ( .A(KEYINPUT76), .ZN(n496) );
  XNOR2_X1 U596 ( .A(n496), .B(KEYINPUT38), .ZN(n497) );
  XNOR2_X1 U597 ( .A(n363), .B(n497), .ZN(n754) );
  INV_X1 U598 ( .A(KEYINPUT88), .ZN(n498) );
  XNOR2_X1 U599 ( .A(n498), .B(KEYINPUT39), .ZN(n499) );
  NAND2_X1 U600 ( .A1(G217), .A2(n501), .ZN(n503) );
  XOR2_X1 U601 ( .A(n504), .B(KEYINPUT9), .Z(n505) );
  XNOR2_X1 U602 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U603 ( .A(n510), .B(n509), .ZN(n693) );
  NOR2_X1 U604 ( .A1(G902), .A2(n693), .ZN(n514) );
  INV_X1 U605 ( .A(G478), .ZN(n512) );
  XOR2_X1 U606 ( .A(KEYINPUT13), .B(KEYINPUT103), .Z(n516) );
  XNOR2_X1 U607 ( .A(KEYINPUT102), .B(G475), .ZN(n515) );
  XNOR2_X1 U608 ( .A(n516), .B(n515), .ZN(n529) );
  XNOR2_X1 U609 ( .A(n518), .B(n517), .ZN(n522) );
  XOR2_X1 U610 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n520) );
  XNOR2_X1 U611 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U612 ( .A(n522), .B(n521), .ZN(n527) );
  XOR2_X1 U613 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n525) );
  NAND2_X1 U614 ( .A1(G214), .A2(n523), .ZN(n524) );
  XNOR2_X1 U615 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U616 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U617 ( .A(n528), .B(n561), .ZN(n666) );
  XNOR2_X1 U618 ( .A(n529), .B(n417), .ZN(n542) );
  INV_X1 U619 ( .A(n542), .ZN(n581) );
  NOR2_X1 U620 ( .A1(n580), .A2(n581), .ZN(n531) );
  INV_X1 U621 ( .A(KEYINPUT105), .ZN(n530) );
  XNOR2_X1 U622 ( .A(n531), .B(n530), .ZN(n711) );
  NAND2_X1 U623 ( .A1(n367), .A2(n711), .ZN(n604) );
  XNOR2_X1 U624 ( .A(n604), .B(G134), .ZN(G36) );
  XNOR2_X1 U625 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n533) );
  INV_X1 U626 ( .A(KEYINPUT71), .ZN(n532) );
  INV_X1 U627 ( .A(G898), .ZN(n534) );
  NAND2_X1 U628 ( .A1(n534), .A2(G953), .ZN(n535) );
  XNOR2_X1 U629 ( .A(n535), .B(KEYINPUT96), .ZN(n783) );
  OR2_X1 U630 ( .A1(n783), .A2(n536), .ZN(n538) );
  NAND2_X1 U631 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U632 ( .A1(n580), .A2(n542), .ZN(n756) );
  NOR2_X1 U633 ( .A1(n756), .A2(n741), .ZN(n543) );
  INV_X1 U634 ( .A(KEYINPUT22), .ZN(n544) );
  INV_X1 U635 ( .A(n566), .ZN(n546) );
  OR2_X1 U636 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U637 ( .A1(n547), .A2(n362), .ZN(n548) );
  AND2_X1 U638 ( .A1(n556), .A2(n548), .ZN(n617) );
  XOR2_X1 U639 ( .A(G110), .B(n617), .Z(G12) );
  NAND2_X1 U640 ( .A1(n549), .A2(n619), .ZN(n565) );
  NAND2_X1 U641 ( .A1(n717), .A2(n620), .ZN(n550) );
  AND2_X1 U642 ( .A1(n574), .A2(n753), .ZN(n551) );
  INV_X1 U643 ( .A(n738), .ZN(n557) );
  NAND2_X1 U644 ( .A1(n551), .A2(n557), .ZN(n552) );
  XNOR2_X1 U645 ( .A(n552), .B(KEYINPUT43), .ZN(n553) );
  INV_X1 U646 ( .A(n363), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n553), .A2(n583), .ZN(n605) );
  XNOR2_X1 U648 ( .A(n605), .B(G140), .ZN(G42) );
  INV_X1 U649 ( .A(KEYINPUT40), .ZN(n554) );
  XOR2_X1 U650 ( .A(G131), .B(n572), .Z(G33) );
  INV_X1 U651 ( .A(n620), .ZN(n555) );
  NAND2_X1 U652 ( .A1(n616), .A2(n557), .ZN(n559) );
  INV_X1 U653 ( .A(KEYINPUT89), .ZN(n558) );
  XNOR2_X1 U654 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U655 ( .A(n619), .B(KEYINPUT106), .ZN(n742) );
  XNOR2_X1 U656 ( .A(n373), .B(G101), .ZN(G3) );
  XOR2_X1 U657 ( .A(KEYINPUT126), .B(n561), .Z(n562) );
  XNOR2_X1 U658 ( .A(n563), .B(n562), .ZN(n609) );
  XNOR2_X1 U659 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n564) );
  OR2_X1 U660 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U661 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n567) );
  XNOR2_X1 U662 ( .A(n568), .B(n567), .ZN(n570) );
  INV_X1 U663 ( .A(n640), .ZN(n569) );
  NOR2_X1 U664 ( .A1(n752), .A2(n588), .ZN(n571) );
  XNOR2_X1 U665 ( .A(n571), .B(KEYINPUT42), .ZN(n791) );
  XNOR2_X1 U666 ( .A(n573), .B(KEYINPUT46), .ZN(n601) );
  XNOR2_X1 U667 ( .A(n574), .B(KEYINPUT113), .ZN(n576) );
  NOR2_X1 U668 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U669 ( .A(n577), .B(KEYINPUT36), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n578), .A2(n362), .ZN(n579) );
  INV_X1 U671 ( .A(n580), .ZN(n582) );
  NAND2_X1 U672 ( .A1(n582), .A2(n581), .ZN(n626) );
  NOR2_X1 U673 ( .A1(n626), .A2(n583), .ZN(n584) );
  NAND2_X1 U674 ( .A1(n585), .A2(n584), .ZN(n715) );
  INV_X1 U675 ( .A(KEYINPUT83), .ZN(n590) );
  OR2_X1 U676 ( .A1(KEYINPUT47), .A2(n590), .ZN(n586) );
  AND2_X1 U677 ( .A1(n715), .A2(n586), .ZN(n587) );
  AND2_X1 U678 ( .A1(n789), .A2(n587), .ZN(n594) );
  OR2_X1 U679 ( .A1(n711), .A2(n717), .ZN(n645) );
  INV_X1 U680 ( .A(n645), .ZN(n758) );
  NAND2_X1 U681 ( .A1(n758), .A2(n590), .ZN(n591) );
  NAND2_X1 U682 ( .A1(n718), .A2(n591), .ZN(n592) );
  NAND2_X1 U683 ( .A1(n592), .A2(KEYINPUT47), .ZN(n593) );
  NAND2_X1 U684 ( .A1(n594), .A2(n593), .ZN(n599) );
  INV_X1 U685 ( .A(KEYINPUT47), .ZN(n595) );
  NAND2_X1 U686 ( .A1(n718), .A2(n595), .ZN(n596) );
  NAND2_X1 U687 ( .A1(n596), .A2(n590), .ZN(n597) );
  AND2_X1 U688 ( .A1(n597), .A2(n645), .ZN(n598) );
  NOR2_X1 U689 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U690 ( .A1(n601), .A2(n600), .ZN(n603) );
  INV_X1 U691 ( .A(KEYINPUT48), .ZN(n602) );
  XNOR2_X1 U692 ( .A(n603), .B(n602), .ZN(n607) );
  AND2_X1 U693 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U694 ( .A(n609), .B(n733), .Z(n608) );
  NAND2_X1 U695 ( .A1(n608), .A2(n774), .ZN(n613) );
  XNOR2_X1 U696 ( .A(G227), .B(n609), .ZN(n610) );
  NAND2_X1 U697 ( .A1(n610), .A2(G900), .ZN(n611) );
  NAND2_X1 U698 ( .A1(G953), .A2(n611), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n613), .A2(n612), .ZN(G72) );
  NAND2_X1 U700 ( .A1(n738), .A2(n742), .ZN(n614) );
  XOR2_X1 U701 ( .A(n618), .B(G119), .Z(G21) );
  NOR2_X1 U702 ( .A1(n741), .A2(n619), .ZN(n739) );
  AND2_X1 U703 ( .A1(n620), .A2(n739), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n621), .A2(n738), .ZN(n623) );
  INV_X1 U705 ( .A(KEYINPUT33), .ZN(n622) );
  XNOR2_X2 U706 ( .A(n623), .B(n622), .ZN(n725) );
  BUF_X2 U707 ( .A(n624), .Z(n637) );
  NAND2_X1 U708 ( .A1(n374), .A2(n366), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n628), .A2(KEYINPUT44), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n629), .A2(KEYINPUT68), .ZN(n634) );
  INV_X1 U711 ( .A(KEYINPUT68), .ZN(n630) );
  AND2_X1 U712 ( .A1(n630), .A2(KEYINPUT44), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n650) );
  AND2_X1 U714 ( .A1(n738), .A2(n739), .ZN(n636) );
  INV_X1 U715 ( .A(n641), .ZN(n744) );
  NAND2_X1 U716 ( .A1(n636), .A2(n744), .ZN(n748) );
  INV_X1 U717 ( .A(n637), .ZN(n644) );
  OR2_X1 U718 ( .A1(n748), .A2(n644), .ZN(n639) );
  INV_X1 U719 ( .A(KEYINPUT31), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n639), .B(n638), .ZN(n722) );
  AND2_X1 U721 ( .A1(n739), .A2(n640), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  OR2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n708) );
  NAND2_X1 U724 ( .A1(n722), .A2(n708), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(n655) );
  NOR2_X1 U728 ( .A1(n787), .A2(KEYINPUT44), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n370), .B(KEYINPUT91), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n655), .A2(n369), .ZN(n657) );
  INV_X1 U731 ( .A(KEYINPUT2), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n659), .A2(KEYINPUT2), .ZN(n661) );
  INV_X1 U733 ( .A(KEYINPUT70), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U735 ( .A1(n696), .A2(G475), .ZN(n668) );
  XNOR2_X1 U736 ( .A(KEYINPUT69), .B(KEYINPUT122), .ZN(n664) );
  XOR2_X1 U737 ( .A(n664), .B(KEYINPUT59), .Z(n665) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(n670) );
  INV_X1 U739 ( .A(G952), .ZN(n669) );
  NAND2_X1 U740 ( .A1(n669), .A2(G953), .ZN(n690) );
  NAND2_X1 U741 ( .A1(n670), .A2(n690), .ZN(n672) );
  XNOR2_X1 U742 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n671) );
  XNOR2_X1 U743 ( .A(n672), .B(n671), .ZN(G60) );
  NAND2_X1 U744 ( .A1(n696), .A2(G472), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U746 ( .A1(n676), .A2(n690), .ZN(n678) );
  XNOR2_X1 U747 ( .A(KEYINPUT92), .B(KEYINPUT63), .ZN(n677) );
  XNOR2_X1 U748 ( .A(n678), .B(n677), .ZN(G57) );
  NAND2_X1 U749 ( .A1(n372), .A2(G210), .ZN(n683) );
  BUF_X1 U750 ( .A(n679), .Z(n681) );
  XNOR2_X1 U751 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n683), .B(n682), .ZN(n684) );
  NAND2_X1 U753 ( .A1(n684), .A2(n690), .ZN(n687) );
  XNOR2_X1 U754 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n685), .B(KEYINPUT87), .ZN(n686) );
  XNOR2_X1 U756 ( .A(n687), .B(n686), .ZN(G51) );
  NAND2_X1 U757 ( .A1(n692), .A2(G217), .ZN(n689) );
  XNOR2_X1 U758 ( .A(n689), .B(n688), .ZN(n691) );
  INV_X1 U759 ( .A(n690), .ZN(n702) );
  NOR2_X1 U760 ( .A1(n691), .A2(n702), .ZN(G66) );
  NAND2_X1 U761 ( .A1(n692), .A2(G478), .ZN(n694) );
  XNOR2_X1 U762 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n695), .A2(n702), .ZN(G63) );
  NAND2_X1 U764 ( .A1(n692), .A2(G469), .ZN(n701) );
  XNOR2_X1 U765 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n697) );
  XNOR2_X1 U766 ( .A(n697), .B(KEYINPUT57), .ZN(n698) );
  XNOR2_X1 U767 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U768 ( .A(n701), .B(n700), .ZN(n703) );
  NOR2_X1 U769 ( .A1(n703), .A2(n702), .ZN(G54) );
  NOR2_X1 U770 ( .A1(n720), .A2(n708), .ZN(n705) );
  XNOR2_X1 U771 ( .A(G104), .B(KEYINPUT115), .ZN(n704) );
  XNOR2_X1 U772 ( .A(n705), .B(n704), .ZN(G6) );
  XOR2_X1 U773 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n707) );
  XNOR2_X1 U774 ( .A(G107), .B(KEYINPUT116), .ZN(n706) );
  XNOR2_X1 U775 ( .A(n707), .B(n706), .ZN(n710) );
  INV_X1 U776 ( .A(n711), .ZN(n723) );
  NOR2_X1 U777 ( .A1(n723), .A2(n708), .ZN(n709) );
  XOR2_X1 U778 ( .A(n710), .B(n709), .Z(G9) );
  XOR2_X1 U779 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n713) );
  NAND2_X1 U780 ( .A1(n718), .A2(n711), .ZN(n712) );
  XNOR2_X1 U781 ( .A(n713), .B(n712), .ZN(n714) );
  XOR2_X1 U782 ( .A(G128), .B(n714), .Z(G30) );
  XNOR2_X1 U783 ( .A(n715), .B(G143), .ZN(n716) );
  XNOR2_X1 U784 ( .A(KEYINPUT118), .B(n716), .ZN(G45) );
  NAND2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U786 ( .A(n719), .B(G146), .ZN(G48) );
  NOR2_X1 U787 ( .A1(n720), .A2(n722), .ZN(n721) );
  XOR2_X1 U788 ( .A(G113), .B(n721), .Z(G15) );
  NOR2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U790 ( .A(G116), .B(n724), .Z(G18) );
  BUF_X1 U791 ( .A(n725), .Z(n726) );
  NOR2_X1 U792 ( .A1(n752), .A2(n726), .ZN(n727) );
  NOR2_X1 U793 ( .A1(G953), .A2(n727), .ZN(n772) );
  BUF_X1 U794 ( .A(n728), .Z(n729) );
  XNOR2_X1 U795 ( .A(n730), .B(KEYINPUT85), .ZN(n731) );
  NAND2_X1 U796 ( .A1(n732), .A2(n731), .ZN(n736) );
  NOR2_X1 U797 ( .A1(n733), .A2(KEYINPUT2), .ZN(n734) );
  XNOR2_X1 U798 ( .A(n734), .B(KEYINPUT86), .ZN(n735) );
  NOR2_X1 U799 ( .A1(n736), .A2(n735), .ZN(n770) );
  INV_X1 U800 ( .A(n737), .ZN(n768) );
  NOR2_X1 U801 ( .A1(n739), .A2(n362), .ZN(n740) );
  XOR2_X1 U802 ( .A(KEYINPUT50), .B(n740), .Z(n747) );
  NAND2_X1 U803 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U804 ( .A(n743), .B(KEYINPUT49), .ZN(n745) );
  NOR2_X1 U805 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U806 ( .A1(n747), .A2(n746), .ZN(n749) );
  AND2_X1 U807 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U808 ( .A(KEYINPUT51), .B(n750), .Z(n751) );
  NOR2_X1 U809 ( .A1(n752), .A2(n751), .ZN(n763) );
  NOR2_X1 U810 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U811 ( .A1(n756), .A2(n755), .ZN(n760) );
  NOR2_X1 U812 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U813 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U814 ( .A1(n761), .A2(n726), .ZN(n762) );
  NOR2_X1 U815 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U816 ( .A(n764), .B(KEYINPUT119), .ZN(n765) );
  XNOR2_X1 U817 ( .A(n765), .B(KEYINPUT52), .ZN(n766) );
  NAND2_X1 U818 ( .A1(n766), .A2(G952), .ZN(n767) );
  NOR2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U820 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U821 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U822 ( .A(KEYINPUT53), .B(n773), .Z(G75) );
  NAND2_X1 U823 ( .A1(n729), .A2(n774), .ZN(n778) );
  NAND2_X1 U824 ( .A1(G953), .A2(G224), .ZN(n775) );
  XNOR2_X1 U825 ( .A(KEYINPUT61), .B(n775), .ZN(n776) );
  NAND2_X1 U826 ( .A1(n776), .A2(G898), .ZN(n777) );
  NAND2_X1 U827 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U828 ( .A(n779), .B(KEYINPUT125), .ZN(n786) );
  XNOR2_X1 U829 ( .A(n780), .B(KEYINPUT124), .ZN(n782) );
  XNOR2_X1 U830 ( .A(n782), .B(n781), .ZN(n784) );
  AND2_X1 U831 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U832 ( .A(n786), .B(n785), .Z(G69) );
  XNOR2_X1 U833 ( .A(n787), .B(G122), .ZN(n788) );
  XNOR2_X1 U834 ( .A(n788), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U835 ( .A(G125), .B(n789), .Z(n790) );
  XNOR2_X1 U836 ( .A(KEYINPUT37), .B(n790), .ZN(G27) );
  XOR2_X1 U837 ( .A(G137), .B(n791), .Z(G39) );
endmodule

