//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n561, new_n562, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT66), .A2(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT67), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n470), .B2(KEYINPUT67), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n465), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n466), .A2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n464), .ZN(new_n481));
  INV_X1    g056(.A(G137), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n475), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n465), .A2(new_n480), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n468), .A2(G2105), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n488), .A2(G124), .B1(G136), .B2(new_n489), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n464), .C2(G112), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT68), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n476), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n480), .A2(G138), .A3(new_n464), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n480), .A2(new_n501), .A3(G138), .A4(new_n464), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT69), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(G543), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n509), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n520), .A2(new_n504), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n513), .A2(new_n519), .A3(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND2_X1  g098(.A1(new_n518), .A2(G89), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n512), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(new_n528), .B1(new_n516), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n524), .A2(new_n525), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n518), .A2(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n512), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n504), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND4_X1  g113(.A1(new_n509), .A2(G43), .A3(G543), .A4(new_n510), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n509), .A2(G81), .A3(new_n510), .A4(new_n516), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n514), .B2(new_n515), .ZN(new_n544));
  INV_X1    g119(.A(G68), .ZN(new_n545));
  INV_X1    g120(.A(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT70), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  AND2_X1   g125(.A1(KEYINPUT5), .A2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(KEYINPUT5), .A2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g128(.A(new_n549), .B(new_n550), .C1(new_n553), .C2(new_n543), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n548), .A2(new_n554), .A3(G651), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n541), .A2(new_n542), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n542), .B1(new_n541), .B2(new_n555), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  AND2_X1   g138(.A1(G53), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n506), .B1(new_n507), .B2(G651), .ZN(new_n565));
  NOR3_X1   g140(.A1(new_n504), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n510), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n505), .A2(new_n508), .B1(KEYINPUT6), .B2(new_n504), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n570), .A2(KEYINPUT72), .A3(new_n564), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(KEYINPUT9), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n509), .A2(new_n573), .A3(new_n510), .A4(new_n564), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n574), .A2(KEYINPUT73), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n569), .A2(new_n571), .A3(new_n577), .A4(KEYINPUT9), .ZN(new_n578));
  AND4_X1   g153(.A1(G91), .A2(new_n509), .A3(new_n510), .A4(new_n516), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n514), .B2(new_n515), .ZN(new_n581));
  AND2_X1   g156(.A1(G78), .A2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g160(.A(KEYINPUT74), .B(G651), .C1(new_n581), .C2(new_n582), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n579), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n576), .A2(new_n578), .A3(new_n587), .ZN(G299));
  NAND2_X1  g163(.A1(new_n512), .A2(G49), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n518), .A2(G87), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n512), .A2(G48), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n518), .A2(G86), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n504), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(KEYINPUT75), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(KEYINPUT75), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n518), .A2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n512), .A2(G47), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(new_n504), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(G290));
  XNOR2_X1  g181(.A(KEYINPUT76), .B(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n517), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n516), .A2(G66), .ZN(new_n610));
  AND2_X1   g185(.A1(G79), .A2(G543), .ZN(new_n611));
  OAI21_X1  g186(.A(G651), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n607), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n570), .A2(G92), .A3(new_n516), .A4(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n570), .A2(G54), .A3(G543), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n609), .A2(new_n612), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G171), .B2(new_n617), .ZN(G284));
  OAI21_X1  g194(.A(new_n618), .B1(G171), .B2(new_n617), .ZN(G321));
  NOR2_X1   g195(.A1(G286), .A2(new_n617), .ZN(new_n621));
  XNOR2_X1  g196(.A(G299), .B(KEYINPUT77), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n617), .ZN(G297));
  AOI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n617), .ZN(G280));
  INV_X1    g199(.A(new_n616), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT78), .B(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(G860), .B2(new_n626), .ZN(G148));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n558), .B2(G868), .ZN(G323));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n631));
  XNOR2_X1  g206(.A(G323), .B(new_n631), .ZN(G282));
  NAND2_X1  g207(.A1(new_n480), .A2(new_n478), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n489), .A2(G135), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT80), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n488), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n464), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n638), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n636), .A2(G2100), .B1(new_n642), .B2(G2096), .ZN(new_n643));
  INV_X1    g218(.A(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n643), .B(new_n645), .C1(G2096), .C2(new_n642), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT81), .Z(G156));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n651), .B(new_n657), .Z(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n661), .A3(G14), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT82), .ZN(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(new_n644), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(G2096), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT83), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n677), .A2(new_n679), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n682), .A3(new_n680), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n684), .B(new_n687), .C1(new_n682), .C2(new_n686), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1981), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT84), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(G229));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G6), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n600), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n696), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n696), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n696), .A2(G23), .ZN(new_n706));
  INV_X1    g281(.A(G288), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(new_n696), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n700), .A2(new_n701), .A3(new_n705), .A4(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n488), .A2(G119), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT85), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n464), .A2(G107), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n718), .A2(new_n720), .B1(new_n489), .B2(G131), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n715), .B1(new_n723), .B2(new_n714), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n696), .A2(G24), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT86), .Z(new_n728));
  INV_X1    g303(.A(G290), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n696), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT87), .B(G1986), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n712), .A2(new_n713), .A3(new_n726), .A4(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT36), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n714), .A2(G35), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G162), .B2(new_n714), .ZN(new_n736));
  INV_X1    g311(.A(G2090), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  NOR2_X1   g316(.A1(new_n642), .A2(new_n714), .ZN(new_n742));
  INV_X1    g317(.A(G28), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n743), .B2(KEYINPUT30), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n741), .B(new_n742), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n714), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n488), .A2(G128), .ZN(new_n750));
  NOR2_X1   g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT89), .Z(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n489), .A2(G140), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n749), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2067), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(G29), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n758), .B2(new_n759), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G160), .B2(new_n714), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n746), .B(new_n757), .C1(G2084), .C2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G32), .ZN(new_n764));
  AOI21_X1  g339(.A(KEYINPUT92), .B1(new_n714), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n489), .A2(G141), .ZN(new_n766));
  INV_X1    g341(.A(G105), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n477), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT26), .Z(new_n770));
  INV_X1    g345(.A(G129), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n487), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  MUX2_X1   g349(.A(KEYINPUT92), .B(new_n765), .S(new_n774), .Z(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  NOR2_X1   g352(.A1(G27), .A2(G29), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G164), .B2(G29), .ZN(new_n779));
  OAI22_X1  g354(.A1(new_n775), .A2(new_n777), .B1(new_n779), .B2(G2078), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n775), .A2(new_n777), .ZN(new_n781));
  INV_X1    g356(.A(G2078), .ZN(new_n782));
  INV_X1    g357(.A(new_n779), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G4), .A2(G16), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n625), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT88), .B(G1348), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n763), .A2(new_n780), .A3(new_n784), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n714), .A2(G33), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT25), .Z(new_n792));
  AOI22_X1  g367(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(new_n464), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n489), .A2(G139), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT91), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n790), .B1(new_n800), .B2(new_n714), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G2072), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n696), .A2(G21), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G168), .B2(new_n696), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT94), .B(G1966), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G2084), .B2(new_n762), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n804), .A2(new_n806), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n740), .A2(new_n789), .A3(new_n802), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n696), .A2(G5), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G171), .B2(new_n696), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT95), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G1341), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n558), .A2(new_n696), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n696), .B2(G19), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n815), .A2(G1961), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n696), .A2(G20), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT23), .Z(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G299), .B2(G16), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1956), .ZN(new_n823));
  INV_X1    g398(.A(new_n818), .ZN(new_n824));
  INV_X1    g399(.A(G1961), .ZN(new_n825));
  AOI22_X1  g400(.A1(G1341), .A2(new_n824), .B1(new_n814), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n819), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n734), .A2(new_n811), .A3(new_n827), .ZN(G311));
  INV_X1    g403(.A(G311), .ZN(G150));
  NAND2_X1  g404(.A1(new_n541), .A2(new_n555), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT71), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n832));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  AND2_X1   g408(.A1(G80), .A2(G543), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n516), .B2(G67), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n511), .A2(new_n833), .B1(new_n835), .B2(new_n504), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n517), .A2(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n541), .A2(new_n555), .A3(new_n542), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n831), .A2(new_n832), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n836), .A2(new_n838), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n556), .A2(new_n557), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n830), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT98), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n841), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n625), .A2(G559), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n846), .B(new_n847), .Z(new_n848));
  XOR2_X1   g423(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  INV_X1    g426(.A(G860), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n842), .A2(new_n852), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n642), .B(G160), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n493), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n722), .B(new_n634), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n488), .A2(G130), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT100), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n489), .A2(G142), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n464), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n863), .B(new_n864), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n861), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G164), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n871));
  INV_X1    g446(.A(new_n773), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n800), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n798), .A2(new_n871), .A3(new_n799), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n773), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n755), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n755), .B1(new_n873), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n870), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(G164), .A3(new_n876), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n869), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n881), .A3(new_n869), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(KEYINPUT101), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n885));
  AOI211_X1 g460(.A(new_n885), .B(new_n869), .C1(new_n879), .C2(new_n881), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n860), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n882), .A2(new_n860), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n888), .B2(new_n883), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n889), .A3(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(G395));
  NAND4_X1  g470(.A1(new_n576), .A2(new_n616), .A3(new_n587), .A4(new_n578), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n896), .A2(KEYINPUT41), .ZN(new_n897));
  AND3_X1   g472(.A1(G299), .A2(KEYINPUT103), .A3(new_n625), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT103), .B1(G299), .B2(new_n625), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT105), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n897), .B(new_n905), .C1(new_n898), .C2(new_n899), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n846), .B(new_n628), .Z(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n902), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(KEYINPUT104), .B(new_n896), .C1(new_n898), .C2(new_n899), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(new_n908), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n909), .A2(new_n914), .A3(KEYINPUT42), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT42), .B1(new_n909), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G303), .B(G288), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n600), .A2(new_n729), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G290), .B1(new_n598), .B2(new_n599), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n918), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n919), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n917), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n617), .B1(new_n917), .B2(new_n926), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(KEYINPUT106), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT106), .B1(new_n842), .B2(G868), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n927), .B2(new_n928), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n930), .A2(new_n932), .ZN(G295));
  NOR2_X1   g508(.A1(new_n930), .A2(new_n932), .ZN(G331));
  NAND3_X1  g509(.A1(new_n831), .A2(new_n840), .A3(new_n839), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n832), .B1(new_n842), .B2(new_n830), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n937), .A2(G301), .A3(new_n841), .ZN(new_n938));
  AOI21_X1  g513(.A(G301), .B1(new_n937), .B2(new_n841), .ZN(new_n939));
  OAI21_X1  g514(.A(G286), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n846), .A2(G171), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(G301), .A3(new_n841), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(G168), .A3(new_n942), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n940), .A2(new_n943), .B1(new_n911), .B2(new_n912), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n926), .B1(new_n944), .B2(KEYINPUT109), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n911), .A2(new_n912), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n938), .A2(new_n939), .A3(G286), .ZN(new_n947));
  AOI21_X1  g522(.A(G168), .B1(new_n941), .B2(new_n942), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n904), .A2(new_n900), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n943), .A3(new_n940), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n907), .A2(new_n943), .A3(new_n940), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n902), .B1(new_n947), .B2(new_n948), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n926), .A3(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n956), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n964), .A2(KEYINPUT110), .A3(new_n955), .A4(new_n954), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n957), .A2(new_n958), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n926), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n957), .A2(KEYINPUT107), .A3(new_n958), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n963), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n967), .B1(new_n972), .B2(new_n955), .ZN(new_n973));
  INV_X1    g548(.A(new_n971), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT107), .B1(new_n957), .B2(new_n958), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n974), .A2(new_n975), .A3(new_n926), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT108), .B(KEYINPUT43), .C1(new_n976), .C2(new_n963), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n966), .A2(new_n973), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n964), .A2(KEYINPUT43), .A3(new_n954), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT44), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(G397));
  NOR2_X1   g559(.A1(G164), .A2(G1384), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n475), .A2(G40), .A3(new_n484), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n722), .B(new_n725), .Z(new_n989));
  INV_X1    g564(.A(G2067), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n755), .B(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n773), .B(G1996), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(G290), .B(G1986), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n988), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G303), .A2(G8), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT55), .ZN(new_n999));
  OR2_X1    g574(.A1(G164), .A2(G1384), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n987), .B1(new_n1000), .B2(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n985), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G2090), .B1(new_n1004), .B2(KEYINPUT116), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1001), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1007));
  INV_X1    g582(.A(new_n987), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n986), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1005), .A2(new_n1007), .B1(new_n704), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n1012));
  OAI21_X1  g587(.A(G8), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1010), .A2(new_n704), .ZN(new_n1014));
  AOI211_X1 g589(.A(KEYINPUT117), .B(new_n1014), .C1(new_n1007), .C2(new_n1005), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n999), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1000), .A2(new_n987), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n707), .A2(G1976), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT113), .B(G1976), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n1026));
  INV_X1    g601(.A(new_n597), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n597), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n1029), .A2(new_n1030), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1019), .B1(new_n1032), .B2(KEYINPUT49), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1022), .B(new_n1025), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n999), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n985), .A2(KEYINPUT111), .A3(new_n1002), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT111), .B1(new_n985), .B2(new_n1002), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1001), .B(new_n737), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1041), .A2(KEYINPUT112), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1041), .A2(KEYINPUT112), .B1(new_n704), .B2(new_n1010), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1018), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1036), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1010), .A2(new_n805), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1001), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(G2084), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G286), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1016), .A2(new_n1045), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT63), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1044), .A2(new_n1037), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1045), .A2(new_n1054), .A3(KEYINPUT63), .A4(new_n1050), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1016), .A2(new_n1045), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT124), .B(G1961), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n986), .A2(new_n782), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1047), .A2(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(G2078), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n986), .A2(new_n1008), .A3(new_n1009), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(G301), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G168), .A2(new_n1018), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT51), .B1(new_n1065), .B2(KEYINPUT123), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1049), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1067), .ZN(new_n1069));
  OAI211_X1 g644(.A(G8), .B(new_n1069), .C1(new_n1048), .C2(G286), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1048), .A2(new_n1065), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT62), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1071), .A2(KEYINPUT62), .A3(new_n1072), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1057), .B(new_n1064), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1076));
  OR2_X1    g651(.A1(G288), .A2(G1976), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1019), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1036), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1081), .A2(new_n1044), .A3(new_n1037), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1080), .A2(new_n1082), .A3(KEYINPUT115), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1056), .A2(new_n1075), .A3(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n483), .A2(KEYINPUT125), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1062), .A2(G40), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n483), .B2(KEYINPUT125), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1089), .A2(new_n475), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n986), .A2(new_n1009), .A3(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT126), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n1061), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(G171), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1061), .A2(G301), .A3(new_n1063), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(KEYINPUT54), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT127), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1096), .A2(KEYINPUT127), .A3(KEYINPUT54), .A4(new_n1097), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1095), .A2(G171), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1064), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1102), .A2(new_n1057), .A3(new_n1103), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1956), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1004), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n986), .A2(new_n1008), .A3(new_n1009), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G299), .B(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(KEYINPUT119), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1112), .A2(new_n1117), .A3(new_n1114), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1120));
  INV_X1    g695(.A(G1348), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1047), .A2(new_n1121), .B1(new_n990), .B2(new_n1017), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1120), .B1(new_n625), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1120), .A2(KEYINPUT61), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT61), .B1(new_n1120), .B2(new_n1115), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1122), .A2(KEYINPUT60), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(new_n625), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1123), .A2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1127), .A2(new_n1128), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n1134));
  INV_X1    g709(.A(new_n558), .ZN(new_n1135));
  INV_X1    g710(.A(G1996), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n986), .A2(new_n1136), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT58), .B(G1341), .Z(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1000), .B2(new_n987), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1137), .A2(KEYINPUT120), .A3(new_n1139), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1135), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1134), .B1(new_n1145), .B2(KEYINPUT59), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n1147));
  OR3_X1    g722(.A1(new_n1144), .A2(KEYINPUT121), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(KEYINPUT122), .A3(new_n1147), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1146), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1125), .B1(new_n1133), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1107), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n997), .B1(new_n1088), .B2(new_n1153), .ZN(new_n1154));
  NOR4_X1   g729(.A1(new_n986), .A2(G1986), .A3(G290), .A4(new_n987), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n995), .A2(new_n988), .B1(KEYINPUT48), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(KEYINPUT48), .B2(new_n1155), .ZN(new_n1157));
  INV_X1    g732(.A(new_n991), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n988), .B1(new_n1158), .B2(new_n872), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT46), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(new_n988), .B2(new_n1136), .ZN(new_n1161));
  NOR4_X1   g736(.A1(new_n986), .A2(KEYINPUT46), .A3(G1996), .A4(new_n987), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT47), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n723), .A2(new_n725), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1165), .A2(new_n993), .B1(G2067), .B2(new_n755), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n988), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1157), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1154), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g744(.A(new_n662), .ZN(new_n1171));
  OR4_X1    g745(.A1(new_n460), .A2(G229), .A3(new_n1171), .A4(G227), .ZN(new_n1172));
  AOI21_X1  g746(.A(new_n1172), .B1(new_n887), .B2(new_n889), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n1173), .A2(new_n978), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


