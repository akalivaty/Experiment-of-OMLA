//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G58), .A2(G232), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n205), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n208), .B1(new_n212), .B2(new_n213), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n214), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n210), .A3(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n209), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(G50), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n250), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n256), .B1(G50), .B2(new_n257), .ZN(new_n258));
  XOR2_X1   g0058(.A(new_n258), .B(KEYINPUT69), .Z(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n260), .A2(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(new_n267), .B2(new_n268), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n252), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n259), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT9), .ZN(new_n274));
  INV_X1    g0074(.A(G200), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  AND2_X1   g0076(.A1(G1), .A2(G13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(new_n278), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n280), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n290));
  OAI21_X1  g0090(.A(KEYINPUT66), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT66), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n287), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n294), .B1(new_n292), .B2(new_n293), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n296), .A2(G223), .B1(new_n299), .B2(G77), .ZN(new_n300));
  INV_X1    g0100(.A(G222), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n291), .A2(new_n295), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT67), .B(G1698), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n300), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n286), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G190), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n308), .A2(KEYINPUT73), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(KEYINPUT73), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n274), .B1(new_n275), .B2(new_n307), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT10), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n273), .B1(new_n307), .B2(G169), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n283), .A2(G232), .A3(new_n280), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n282), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G87), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n303), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n288), .A2(KEYINPUT78), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT78), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n325), .A3(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n292), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n321), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n320), .B1(new_n328), .B2(new_n306), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT79), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT79), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n289), .B1(new_n332), .B2(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT67), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n336), .A3(G223), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G226), .A2(G1698), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n283), .B1(new_n340), .B2(new_n321), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n331), .B1(new_n341), .B2(new_n320), .ZN(new_n342));
  AOI21_X1  g0142(.A(G169), .B1(new_n330), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n329), .A2(new_n314), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT80), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n252), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n201), .B1(new_n218), .B2(G58), .ZN(new_n348));
  INV_X1    g0148(.A(G159), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n348), .A2(new_n210), .B1(new_n349), .B2(new_n266), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n327), .A2(new_n210), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT7), .ZN(new_n352));
  AOI21_X1  g0152(.A(G20), .B1(new_n326), .B2(new_n292), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n214), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n350), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n347), .B1(new_n356), .B2(KEYINPUT16), .ZN(new_n357));
  INV_X1    g0157(.A(new_n350), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n291), .A2(new_n210), .A3(new_n295), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n293), .B1(new_n332), .B2(G33), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n354), .A2(G20), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n359), .A2(new_n354), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n358), .B1(new_n362), .B2(new_n219), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT16), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n357), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n253), .ZN(new_n367));
  INV_X1    g0167(.A(new_n260), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n255), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n367), .A2(new_n369), .B1(new_n257), .B2(new_n368), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G169), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n328), .A2(new_n306), .ZN(new_n374));
  INV_X1    g0174(.A(new_n320), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT79), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI211_X1 g0176(.A(new_n331), .B(new_n320), .C1(new_n328), .C2(new_n306), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT80), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n344), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n346), .A2(new_n372), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT18), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n346), .A2(new_n372), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(G200), .B1(new_n330), .B2(new_n342), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n341), .A2(G190), .A3(new_n320), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n366), .B(new_n371), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT17), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n370), .B1(new_n357), .B2(new_n365), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n390), .B(KEYINPUT17), .C1(new_n385), .C2(new_n386), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n382), .A2(new_n384), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT81), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT71), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n260), .B1(new_n394), .B2(new_n266), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n394), .B2(new_n266), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT15), .B(G87), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n347), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n253), .A2(G77), .A3(new_n255), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(G77), .B2(new_n257), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n302), .A2(G238), .A3(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n299), .A2(G107), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n404), .B(new_n405), .C1(new_n304), .C2(new_n231), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n306), .ZN(new_n407));
  INV_X1    g0207(.A(G244), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n282), .B1(new_n284), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT70), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n282), .B(KEYINPUT70), .C1(new_n284), .C2(new_n408), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n403), .B1(new_n415), .B2(new_n373), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n416), .A2(KEYINPUT72), .ZN(new_n417));
  INV_X1    g0217(.A(new_n403), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n413), .B1(new_n406), .B2(new_n306), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n418), .B(KEYINPUT72), .C1(new_n419), .C2(G169), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n314), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n418), .B1(new_n415), .B2(G200), .ZN(new_n424));
  INV_X1    g0224(.A(G190), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n415), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n318), .A2(new_n393), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n218), .A2(new_n210), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n249), .A2(G1), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(KEYINPUT12), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n253), .A2(G68), .A3(new_n255), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n257), .A2(G68), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n431), .B(new_n432), .C1(KEYINPUT12), .C2(new_n433), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n434), .A2(KEYINPUT76), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(KEYINPUT76), .ZN(new_n436));
  INV_X1    g0236(.A(G77), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n263), .A2(new_n437), .B1(new_n242), .B2(new_n266), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n252), .B1(new_n438), .B2(new_n429), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT11), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT13), .ZN(new_n443));
  OAI211_X1 g0243(.A(G226), .B(new_n303), .C1(new_n297), .C2(new_n298), .ZN(new_n444));
  OAI211_X1 g0244(.A(G232), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G97), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT74), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n306), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n282), .B1(new_n284), .B2(new_n220), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n443), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  AOI211_X1 g0253(.A(KEYINPUT13), .B(new_n451), .C1(new_n449), .C2(new_n306), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n442), .B(G169), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n447), .B1(new_n296), .B2(G232), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n283), .B1(new_n456), .B2(new_n444), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT13), .B1(new_n457), .B2(new_n451), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n450), .A2(new_n443), .A3(new_n452), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(G179), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n459), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n442), .B1(new_n462), .B2(G169), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n441), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n441), .B1(new_n462), .B2(G200), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT75), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n453), .A2(new_n454), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n467), .B2(G190), .ZN(new_n468));
  NOR4_X1   g0268(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT75), .A4(new_n425), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g0271(.A(new_n471), .B(KEYINPUT77), .Z(new_n472));
  NAND2_X1  g0272(.A1(new_n428), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT89), .A2(KEYINPUT21), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n254), .A2(G33), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n253), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT87), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n257), .B2(G116), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n250), .A2(KEYINPUT87), .A3(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n476), .A2(G116), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(G20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n252), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT88), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT88), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n252), .A2(new_n485), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n210), .C1(G33), .C2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT20), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n252), .A2(new_n485), .A3(new_n482), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n485), .B1(new_n252), .B2(new_n482), .ZN(new_n493));
  OAI211_X1 g0293(.A(KEYINPUT20), .B(new_n490), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n481), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G169), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT83), .B1(new_n498), .B2(G41), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT83), .ZN(new_n500));
  INV_X1    g0300(.A(G41), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT5), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n254), .B(G45), .C1(new_n501), .C2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n306), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G270), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n504), .B1(new_n499), .B2(new_n502), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT84), .B1(new_n508), .B2(new_n279), .ZN(new_n509));
  AND4_X1   g0309(.A1(KEYINPUT84), .A2(new_n503), .A3(new_n505), .A4(new_n279), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT86), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n303), .A2(G257), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n327), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n334), .A2(new_n336), .A3(G257), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(KEYINPUT86), .A3(new_n292), .A4(new_n326), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n291), .A2(G303), .A3(new_n295), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n326), .A2(G264), .A3(G1698), .A4(new_n292), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n511), .B1(new_n306), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n474), .B1(new_n497), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n478), .A2(new_n480), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n253), .A2(new_n475), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n479), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n491), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n494), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT86), .B1(new_n333), .B2(new_n515), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n306), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n503), .A2(new_n505), .ZN(new_n531));
  INV_X1    g0331(.A(new_n279), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n508), .A2(KEYINPUT84), .A3(new_n279), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(G270), .B2(new_n506), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n529), .A2(G190), .A3(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n526), .B(new_n536), .C1(new_n520), .C2(new_n275), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n529), .A2(G179), .A3(new_n535), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n496), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n529), .A2(new_n535), .ZN(new_n540));
  INV_X1    g0340(.A(new_n474), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n540), .A2(G169), .A3(new_n541), .A4(new_n496), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n521), .A2(new_n537), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n334), .A2(new_n336), .A3(G250), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G257), .A2(G1698), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G294), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n546), .A2(new_n327), .B1(new_n261), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(new_n306), .B1(G264), .B2(new_n506), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n533), .A2(new_n534), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n425), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n506), .A2(G264), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n544), .A2(new_n545), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n333), .A2(new_n553), .B1(G33), .B2(G294), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n554), .B2(new_n283), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n509), .A2(new_n510), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n551), .B1(new_n557), .B2(G200), .ZN(new_n558));
  INV_X1    g0358(.A(G87), .ZN(new_n559));
  OR2_X1    g0359(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n560));
  NAND2_X1  g0360(.A1(KEYINPUT90), .A2(KEYINPUT22), .ZN(new_n561));
  AOI211_X1 g0361(.A(G20), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n302), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n326), .A2(new_n210), .A3(G87), .A4(new_n292), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT22), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT24), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n262), .A2(G116), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n210), .A2(G107), .ZN(new_n569));
  OR3_X1    g0369(.A1(new_n569), .A2(KEYINPUT91), .A3(KEYINPUT23), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT23), .B1(new_n569), .B2(KEYINPUT91), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n302), .A2(new_n562), .B1(new_n564), .B2(KEYINPUT22), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n568), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT24), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n252), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT92), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n430), .B(new_n569), .C1(new_n579), .C2(KEYINPUT25), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(KEYINPUT25), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n581), .ZN(new_n583));
  AOI22_X1  g0383(.A1(G107), .A2(new_n476), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n558), .A2(new_n578), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n557), .A2(new_n314), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n373), .B1(new_n555), .B2(new_n556), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n347), .B1(new_n573), .B2(new_n576), .ZN(new_n588));
  INV_X1    g0388(.A(new_n584), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT93), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT93), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n585), .A2(new_n593), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g0395(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n446), .A2(KEYINPUT74), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n446), .A2(KEYINPUT74), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT19), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(new_n210), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n326), .A2(new_n210), .A3(G68), .A4(new_n292), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n263), .B2(new_n489), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n252), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n398), .A2(new_n257), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n607), .C1(new_n397), .C2(new_n523), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G116), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n303), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n327), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n306), .ZN(new_n612));
  INV_X1    g0412(.A(G45), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(G1), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT85), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n254), .A2(G45), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n615), .A2(new_n618), .A3(new_n283), .A4(G250), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n279), .A2(new_n614), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n612), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n373), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n611), .B2(new_n306), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n314), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n608), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(G20), .B1(new_n447), .B2(KEYINPUT19), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n601), .B(new_n603), .C1(new_n628), .C2(new_n596), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n606), .B1(new_n629), .B2(new_n252), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n625), .A2(G190), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n334), .A2(new_n336), .A3(G238), .ZN(new_n632));
  NAND2_X1  g0432(.A1(G244), .A2(G1698), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n333), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n283), .B1(new_n635), .B2(new_n609), .ZN(new_n636));
  OAI21_X1  g0436(.A(G200), .B1(new_n636), .B2(new_n621), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n476), .A2(G87), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n630), .A2(new_n631), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT4), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n303), .A2(G244), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n327), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n641), .A2(new_n408), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n303), .B(new_n644), .C1(new_n297), .C2(new_n298), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n643), .A2(new_n488), .A3(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(G250), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT82), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT82), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n302), .A2(new_n649), .A3(G250), .A4(G1698), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n283), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n506), .A2(G257), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n550), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(G200), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n654), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n643), .A2(new_n488), .A3(new_n645), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n650), .B2(new_n648), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n656), .B(G190), .C1(new_n658), .C2(new_n283), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n257), .A2(G97), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n476), .B2(G97), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT6), .ZN(new_n663));
  INV_X1    g0463(.A(G107), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n489), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(G97), .A2(G107), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(KEYINPUT6), .A3(G97), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G20), .ZN(new_n670));
  OAI221_X1 g0470(.A(new_n670), .B1(new_n437), .B2(new_n266), .C1(new_n362), .C2(new_n664), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n662), .B1(new_n671), .B2(new_n252), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n655), .A2(new_n659), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n373), .B1(new_n652), .B2(new_n654), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n656), .B(new_n314), .C1(new_n658), .C2(new_n283), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n670), .B1(new_n437), .B2(new_n266), .ZN(new_n676));
  INV_X1    g0476(.A(new_n362), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(G107), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n661), .B1(new_n678), .B2(new_n347), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n674), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n640), .A2(new_n673), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n595), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n473), .A2(new_n543), .A3(new_n682), .ZN(G372));
  INV_X1    g0483(.A(new_n473), .ZN(new_n684));
  INV_X1    g0484(.A(new_n627), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n630), .A2(new_n637), .A3(new_n638), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n686), .A2(new_n687), .B1(G190), .B2(new_n625), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n585), .A3(new_n680), .A4(new_n673), .ZN(new_n691));
  INV_X1    g0491(.A(new_n590), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n521), .A2(new_n539), .A3(new_n542), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n627), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n640), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT26), .B1(new_n696), .B2(new_n680), .ZN(new_n697));
  INV_X1    g0497(.A(new_n680), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n690), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n699), .B2(KEYINPUT26), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n684), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n382), .A2(new_n384), .ZN(new_n703));
  INV_X1    g0503(.A(new_n464), .ZN(new_n704));
  INV_X1    g0504(.A(new_n423), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n704), .B1(new_n470), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n389), .A2(new_n391), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n703), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n316), .B1(new_n312), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n702), .A2(new_n710), .ZN(G369));
  NAND2_X1  g0511(.A1(new_n430), .A2(new_n210), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT95), .Z(new_n714));
  INV_X1    g0514(.A(G213), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n712), .B2(KEYINPUT27), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G343), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n693), .A2(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n595), .A2(new_n720), .B1(new_n692), .B2(new_n719), .ZN(new_n721));
  INV_X1    g0521(.A(new_n719), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n588), .B2(new_n589), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n595), .A2(new_n723), .B1(new_n692), .B2(new_n722), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n719), .A2(new_n526), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n693), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n543), .B2(new_n725), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n721), .B1(new_n724), .B2(new_n728), .ZN(G399));
  INV_X1    g0529(.A(new_n206), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G41), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n596), .A2(new_n479), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n731), .A2(new_n732), .A3(new_n254), .ZN(new_n733));
  INV_X1    g0533(.A(new_n213), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(new_n731), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT28), .Z(new_n736));
  NAND2_X1  g0536(.A1(new_n699), .A2(KEYINPUT26), .ZN(new_n737));
  OR3_X1    g0537(.A1(new_n696), .A2(KEYINPUT26), .A3(new_n680), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n695), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT29), .B1(new_n740), .B2(new_n722), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n701), .A2(new_n719), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(KEYINPUT29), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G330), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n543), .A2(new_n722), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n585), .A2(new_n593), .A3(new_n590), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n593), .B1(new_n585), .B2(new_n590), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n681), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT97), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n595), .A2(KEYINPUT97), .A3(new_n681), .A4(new_n745), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT30), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n656), .B1(new_n658), .B2(new_n283), .ZN(new_n754));
  AOI221_X4 g0554(.A(new_n314), .B1(new_n506), .B2(G270), .C1(new_n533), .C2(new_n534), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n755), .A2(new_n529), .A3(new_n549), .A4(new_n625), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n646), .A2(new_n651), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n654), .B1(new_n758), .B2(new_n306), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n623), .A2(new_n555), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n759), .A2(KEYINPUT30), .A3(new_n538), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n314), .B1(new_n636), .B2(new_n621), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n557), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n754), .A2(new_n540), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n757), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT96), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n719), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n757), .A2(new_n761), .A3(new_n764), .A4(KEYINPUT96), .ZN(new_n768));
  AOI21_X1  g0568(.A(KEYINPUT31), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT31), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n719), .A2(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n744), .B1(new_n752), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n743), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n736), .B1(new_n775), .B2(G1), .ZN(G364));
  NOR2_X1   g0576(.A1(new_n249), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n254), .B1(new_n777), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n731), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n727), .B2(G330), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G330), .B2(new_n727), .ZN(new_n782));
  INV_X1    g0582(.A(new_n780), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n209), .B1(G20), .B2(new_n373), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n210), .A2(G179), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(new_n425), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n664), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n210), .A2(new_n314), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n790), .A2(new_n275), .A3(G190), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n425), .A2(new_n275), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n792), .A2(new_n214), .B1(new_n794), .B2(new_n242), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G190), .A2(G200), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n789), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n788), .B(new_n795), .C1(G77), .C2(new_n798), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n425), .A2(G179), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n210), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G97), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n793), .A2(new_n786), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n559), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n790), .A2(new_n425), .A3(G200), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n805), .B(new_n299), .C1(G58), .C2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n786), .A2(new_n796), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n349), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT32), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n799), .A2(new_n803), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n794), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G326), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT33), .B(G317), .Z(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n792), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G303), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n804), .B1(new_n797), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n299), .B1(new_n547), .B2(new_n801), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n815), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n808), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n806), .A2(G322), .B1(G329), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n820), .B(new_n822), .C1(new_n823), .C2(new_n787), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n785), .B1(new_n811), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(G13), .A2(G33), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G20), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n784), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n247), .A2(new_n613), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n333), .A2(new_n730), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n613), .B2(new_n734), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT98), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n299), .A2(new_n730), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G355), .B1(new_n479), .B2(new_n730), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n783), .B(new_n825), .C1(new_n829), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n828), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n727), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n782), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  NOR2_X1   g0644(.A1(new_n787), .A2(new_n559), .ZN(new_n845));
  XOR2_X1   g0645(.A(KEYINPUT99), .B(G283), .Z(new_n846));
  OAI22_X1  g0646(.A1(new_n792), .A2(new_n846), .B1(new_n804), .B2(new_n664), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(G116), .C2(new_n798), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n794), .A2(new_n816), .B1(new_n808), .B2(new_n817), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G294), .B2(new_n806), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n848), .A2(new_n299), .A3(new_n803), .A4(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n791), .A2(G150), .B1(G159), .B2(new_n798), .ZN(new_n854));
  INV_X1    g0654(.A(G137), .ZN(new_n855));
  INV_X1    g0655(.A(new_n806), .ZN(new_n856));
  XNOR2_X1  g0656(.A(KEYINPUT101), .B(G143), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n854), .B1(new_n855), .B2(new_n794), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT34), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n808), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n787), .A2(new_n214), .ZN(new_n864));
  INV_X1    g0664(.A(new_n804), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n863), .B(new_n864), .C1(G50), .C2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n327), .B1(new_n802), .B2(G58), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n861), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n853), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n851), .A2(new_n852), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n784), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n784), .A2(new_n826), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n783), .B1(new_n437), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n416), .A2(KEYINPUT72), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n420), .A2(new_n421), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n426), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n722), .A2(new_n418), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(KEYINPUT102), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n877), .A2(new_n878), .B1(new_n423), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n871), .B(new_n873), .C1(new_n880), .C2(new_n827), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n701), .B2(new_n719), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n719), .B(new_n880), .C1(new_n695), .C2(new_n700), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT103), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n882), .B(new_n884), .Z(new_n885));
  INV_X1    g0685(.A(new_n774), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n780), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n885), .A2(new_n886), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n881), .B1(new_n888), .B2(new_n889), .ZN(G384));
  NOR2_X1   g0690(.A1(new_n212), .A2(new_n479), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n669), .B(KEYINPUT104), .Z(new_n892));
  INV_X1    g0692(.A(KEYINPUT35), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT36), .ZN(new_n896));
  INV_X1    g0696(.A(G58), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n734), .B(G77), .C1(new_n219), .C2(new_n897), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n254), .B(G13), .C1(new_n898), .C2(new_n243), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(G68), .B1(new_n351), .B2(KEYINPUT7), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n353), .A2(new_n354), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n358), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT106), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n356), .A2(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n364), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n370), .B1(new_n907), .B2(new_n357), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n717), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n392), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n364), .B1(new_n356), .B2(KEYINPUT106), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n904), .B(new_n350), .C1(new_n352), .C2(new_n355), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n357), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n371), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n914), .A2(new_n380), .A3(new_n346), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n387), .B1(new_n908), .B2(new_n717), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n372), .A2(new_n718), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n381), .A2(new_n918), .A3(new_n387), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n910), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n910), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n722), .A2(new_n441), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n464), .A2(new_n470), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(new_n464), .B2(new_n470), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n880), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n765), .A2(new_n766), .ZN(new_n931));
  AND4_X1   g0731(.A1(KEYINPUT31), .A2(new_n931), .A3(new_n722), .A4(new_n768), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(new_n769), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n930), .B1(new_n752), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT107), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT107), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n935), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n392), .A2(new_n372), .A3(new_n718), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n381), .A2(new_n387), .A3(new_n919), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT37), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n920), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT38), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n936), .B1(new_n947), .B2(new_n925), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n934), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n752), .A2(new_n933), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n684), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n952), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(G330), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n428), .A2(new_n472), .A3(new_n743), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n710), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT39), .ZN(new_n958));
  INV_X1    g0758(.A(new_n925), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n946), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n925), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n704), .A2(new_n719), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n703), .A2(new_n718), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n928), .A2(new_n929), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n423), .A2(new_n722), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT105), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n966), .B1(new_n883), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n965), .B1(new_n969), .B2(new_n926), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n964), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n957), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n955), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT109), .Z(new_n974));
  OAI22_X1  g0774(.A1(new_n955), .A2(new_n972), .B1(new_n254), .B2(new_n777), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT108), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(KEYINPUT108), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n900), .B1(new_n977), .B2(new_n978), .ZN(G367));
  OAI221_X1 g0779(.A(new_n829), .B1(new_n206), .B2(new_n397), .C1(new_n832), .C2(new_n237), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(new_n780), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n787), .A2(new_n437), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n792), .A2(new_n349), .B1(new_n808), .B2(new_n855), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(G58), .C2(new_n865), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n802), .A2(G68), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n302), .A3(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n806), .A2(G150), .B1(G50), .B2(new_n798), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n794), .B2(new_n857), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n865), .A2(G116), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT46), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n817), .A2(new_n794), .B1(new_n787), .B2(new_n489), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G317), .B2(new_n821), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G294), .A2(new_n791), .B1(new_n806), .B2(G303), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n992), .A3(new_n327), .A4(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n801), .A2(new_n664), .B1(new_n846), .B2(new_n797), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT113), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n986), .A2(new_n988), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  AOI21_X1  g0798(.A(new_n719), .B1(new_n630), .B2(new_n638), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT110), .Z(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n690), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n627), .B2(new_n1000), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n981), .B1(new_n785), .B2(new_n998), .C1(new_n1002), .C2(new_n841), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n673), .B(new_n680), .C1(new_n672), .C2(new_n719), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(new_n590), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n722), .B1(new_n1005), .B2(new_n680), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1004), .B1(new_n680), .B2(new_n719), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(new_n595), .A3(new_n720), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1006), .B1(new_n1008), .B2(KEYINPUT42), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(KEYINPUT42), .B2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT111), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n724), .A2(new_n728), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n1007), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1015), .B(new_n1017), .Z(new_n1018));
  XOR2_X1   g0818(.A(new_n731), .B(KEYINPUT41), .Z(new_n1019));
  NAND2_X1  g0819(.A1(new_n721), .A2(new_n1007), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT45), .Z(new_n1021));
  NOR2_X1   g0821(.A1(new_n721), .A2(new_n1007), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(KEYINPUT112), .B(KEYINPUT44), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(new_n1016), .ZN(new_n1026));
  MUX2_X1   g0826(.A(new_n724), .B(new_n595), .S(new_n720), .Z(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(new_n728), .Z(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n775), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1019), .B1(new_n1030), .B2(new_n775), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(new_n779), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1003), .B1(new_n1018), .B2(new_n1032), .ZN(G387));
  OAI22_X1  g0833(.A1(new_n856), .A2(new_n242), .B1(new_n794), .B2(new_n349), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G68), .B2(new_n798), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n787), .ZN(new_n1036));
  XOR2_X1   g0836(.A(KEYINPUT115), .B(G150), .Z(new_n1037));
  AOI22_X1  g0837(.A1(new_n1036), .A2(G97), .B1(new_n821), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n791), .A2(new_n368), .B1(G77), .B2(new_n865), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n327), .B1(new_n802), .B2(new_n398), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1036), .A2(G116), .B1(new_n821), .B2(G326), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n801), .A2(new_n846), .B1(new_n804), .B2(new_n547), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n806), .A2(G317), .B1(new_n812), .B2(G322), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n816), .B2(new_n797), .C1(new_n817), .C2(new_n792), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT49), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n327), .B(new_n1042), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1041), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n784), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n234), .A2(new_n613), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1054), .A2(new_n831), .B1(new_n732), .B2(new_n837), .ZN(new_n1055));
  XOR2_X1   g0855(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1056));
  AND3_X1   g0856(.A1(new_n368), .A2(new_n242), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1056), .B1(new_n368), .B2(new_n242), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n613), .B1(new_n214), .B2(new_n437), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n732), .A4(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1055), .A2(new_n1060), .B1(G107), .B2(new_n206), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n783), .B1(new_n1061), .B2(new_n829), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1053), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n724), .B2(new_n828), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n1028), .B2(new_n779), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1029), .A2(new_n731), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1028), .A2(new_n775), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(G393));
  NAND2_X1  g0868(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1030), .A2(new_n731), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1007), .A2(new_n841), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n829), .B1(new_n489), .B2(new_n206), .C1(new_n832), .C2(new_n241), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n821), .A2(G322), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n792), .B2(new_n816), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G294), .B2(new_n798), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n846), .A2(new_n804), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n302), .A2(new_n1076), .A3(new_n788), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1075), .B(new_n1077), .C1(new_n479), .C2(new_n801), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n806), .A2(G311), .B1(new_n812), .B2(G317), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n792), .A2(new_n242), .B1(new_n808), .B2(new_n857), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n368), .B2(new_n798), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n802), .A2(G77), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n327), .B(new_n845), .C1(new_n218), .C2(new_n865), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n806), .A2(G159), .B1(new_n812), .B2(G150), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT51), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1078), .A2(new_n1080), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT116), .Z(new_n1089));
  OAI211_X1 g0889(.A(new_n780), .B(new_n1072), .C1(new_n1089), .C2(new_n785), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1070), .B1(new_n778), .B2(new_n1026), .C1(new_n1071), .C2(new_n1090), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1091), .A2(KEYINPUT117), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(KEYINPUT117), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(G390));
  INV_X1    g0895(.A(new_n966), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n774), .A2(new_n880), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT119), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1097), .B(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n744), .B1(new_n752), .B2(new_n933), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1096), .B1(new_n1100), .B2(new_n880), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n719), .B(new_n880), .C1(new_n739), .C2(new_n695), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n967), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT118), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(KEYINPUT118), .A3(new_n1103), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1101), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1096), .B1(new_n774), .B2(new_n880), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n744), .B(new_n930), .C1(new_n752), .C2(new_n933), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n883), .A2(new_n968), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1099), .A2(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n428), .A2(new_n472), .A3(new_n1100), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n956), .A3(new_n710), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1106), .A2(new_n1096), .A3(new_n1107), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n947), .A2(new_n925), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n962), .A3(new_n1120), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n969), .A2(new_n963), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n960), .A2(new_n961), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1110), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1099), .A2(new_n1124), .A3(new_n1121), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1118), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1114), .A2(new_n1117), .A3(new_n1127), .A4(new_n1126), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n731), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1123), .A2(new_n826), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n856), .A2(new_n479), .B1(new_n794), .B2(new_n823), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G107), .B2(new_n791), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n797), .A2(new_n489), .B1(new_n808), .B2(new_n547), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1135), .A2(new_n864), .A3(new_n805), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1134), .A2(new_n299), .A3(new_n1083), .A4(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G137), .A2(new_n791), .B1(new_n802), .B2(G159), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT120), .Z(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1138), .B1(new_n1141), .B2(new_n797), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT121), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n794), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(G125), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n787), .A2(new_n242), .B1(new_n808), .B2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1145), .B(new_n1147), .C1(G132), .C2(new_n806), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n865), .A2(new_n1037), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n299), .B1(KEYINPUT53), .B2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(KEYINPUT53), .C2(new_n1149), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1137), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n784), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n783), .B1(new_n260), .B2(new_n872), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1132), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n1128), .B2(new_n778), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT122), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1131), .B1(new_n1158), .B2(new_n1159), .ZN(G378));
  AOI21_X1  g0960(.A(new_n744), .B1(new_n948), .B2(new_n934), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n939), .B1(new_n935), .B2(new_n936), .ZN(new_n1162));
  AOI211_X1 g0962(.A(KEYINPUT107), .B(KEYINPUT40), .C1(new_n926), .C2(new_n934), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n971), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n318), .A2(new_n273), .A3(new_n718), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n273), .A2(new_n718), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n312), .A2(new_n317), .A3(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n971), .B(new_n1161), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1166), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1173), .B1(new_n1166), .B2(new_n1174), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1117), .B1(new_n1128), .B2(new_n1113), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n1179), .A3(KEYINPUT57), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT124), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1173), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n971), .B1(new_n941), .B2(new_n1161), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1174), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1166), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(KEYINPUT124), .A3(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1182), .A2(new_n1188), .B1(new_n1117), .B2(new_n1130), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1180), .B(new_n731), .C1(new_n1189), .C2(KEYINPUT57), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n856), .A2(new_n1144), .B1(new_n797), .B2(new_n855), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n792), .A2(new_n862), .B1(new_n794), .B2(new_n1146), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(G150), .C2(new_n802), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n804), .B2(new_n1141), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(G33), .A2(G41), .ZN(new_n1197));
  INV_X1    g0997(.A(G124), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1197), .B1(new_n808), .B2(new_n1198), .C1(new_n349), .C2(new_n787), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1195), .B2(KEYINPUT59), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n806), .A2(G107), .B1(G77), .B2(new_n865), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n787), .A2(new_n897), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G283), .B2(new_n821), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1203), .A3(new_n985), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G116), .A2(new_n812), .B1(new_n798), .B2(new_n398), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n489), .B2(new_n792), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1204), .A2(new_n1206), .A3(G41), .A4(new_n333), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1196), .A2(new_n1200), .B1(KEYINPUT58), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1197), .A2(G50), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n333), .B2(G41), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1207), .B2(KEYINPUT58), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT123), .Z(new_n1212));
  AOI21_X1  g1012(.A(new_n785), .B1(new_n1208), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n872), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n780), .B1(G50), .B2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(new_n1173), .C2(new_n826), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1217), .B2(new_n779), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1191), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(G375));
  OAI22_X1  g1021(.A1(new_n792), .A2(new_n479), .B1(new_n794), .B2(new_n547), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G107), .B2(new_n798), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n982), .B1(G303), .B2(new_n821), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n806), .A2(G283), .B1(G97), .B2(new_n865), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n302), .B1(new_n398), .B2(new_n802), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n794), .A2(new_n862), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n264), .A2(new_n797), .B1(new_n804), .B2(new_n349), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(G137), .C2(new_n806), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n802), .A2(G50), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n327), .B(new_n1202), .C1(G128), .C2(new_n821), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1140), .A2(new_n791), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n785), .B1(new_n1227), .B2(new_n1234), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n783), .B(new_n1235), .C1(new_n214), .C2(new_n872), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1096), .B2(new_n827), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1113), .B2(new_n778), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1019), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1118), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1238), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G381));
  NOR4_X1   g1044(.A1(G387), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1245), .A2(new_n1094), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1156), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1131), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1220), .A3(new_n1243), .A4(new_n1249), .ZN(G407));
  NOR2_X1   g1050(.A1(new_n715), .A2(G343), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1220), .A2(new_n1249), .A3(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G407), .A2(G213), .A3(new_n1252), .ZN(G409));
  OR2_X1    g1053(.A1(new_n1094), .A2(G387), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(G393), .B(new_n843), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1094), .A2(G387), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT61), .ZN(new_n1261));
  INV_X1    g1061(.A(G384), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1118), .A2(new_n731), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1242), .A2(KEYINPUT126), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1242), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1263), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1262), .B1(new_n1268), .B2(new_n1238), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1238), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1267), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT60), .B1(new_n1242), .B2(KEYINPUT126), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G384), .B(new_n1270), .C1(new_n1273), .C2(new_n1263), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT127), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1251), .A2(G2897), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1269), .A2(new_n1274), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1269), .A2(new_n1274), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1276), .B1(new_n1279), .B2(KEYINPUT127), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1275), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1278), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1189), .A2(new_n1239), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1216), .B1(new_n1178), .B2(new_n779), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1248), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT57), .B1(new_n1217), .B2(new_n1179), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1179), .A2(KEYINPUT57), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n731), .B1(new_n1287), .B2(new_n1177), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1218), .C1(new_n1286), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1190), .A2(KEYINPUT125), .A3(G378), .A4(new_n1218), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1285), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1282), .B1(new_n1293), .B2(new_n1251), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1293), .A2(new_n1251), .A3(new_n1279), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1261), .B(new_n1294), .C1(new_n1295), .C2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1285), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1251), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1279), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1303), .A2(KEYINPUT62), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1260), .B1(new_n1297), .B2(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1294), .A2(new_n1261), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1303), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1295), .A2(KEYINPUT63), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1306), .A2(new_n1259), .A3(new_n1308), .A4(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1310), .ZN(G405));
  NAND2_X1  g1111(.A1(G375), .A2(new_n1249), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1298), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1302), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(new_n1279), .A3(new_n1298), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1260), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1259), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(G402));
endmodule


