

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759;

  BUF_X1 U382 ( .A(n718), .Z(n725) );
  AND2_X1 U383 ( .A1(n383), .A2(n427), .ZN(n370) );
  XNOR2_X1 U384 ( .A(n537), .B(KEYINPUT32), .ZN(n758) );
  AND2_X1 U385 ( .A1(n595), .A2(n593), .ZN(n383) );
  NAND2_X1 U386 ( .A1(n367), .A2(n545), .ZN(n546) );
  NOR2_X1 U387 ( .A1(n530), .A2(n678), .ZN(n401) );
  XNOR2_X1 U388 ( .A(n603), .B(n470), .ZN(n586) );
  BUF_X1 U389 ( .A(G113), .Z(n359) );
  XNOR2_X1 U390 ( .A(n454), .B(n453), .ZN(n456) );
  NAND2_X1 U391 ( .A1(n360), .A2(n667), .ZN(n552) );
  NAND2_X1 U392 ( .A1(n700), .A2(n714), .ZN(n360) );
  AND2_X1 U393 ( .A1(n361), .A2(n586), .ZN(n706) );
  INV_X1 U394 ( .A(n588), .ZN(n361) );
  INV_X1 U395 ( .A(G953), .ZN(n748) );
  AND2_X1 U396 ( .A1(n540), .A2(n536), .ZN(n537) );
  AND2_X2 U397 ( .A1(n417), .A2(n422), .ZN(n419) );
  NOR2_X2 U398 ( .A1(n596), .A2(n581), .ZN(n583) );
  NOR2_X2 U399 ( .A1(n755), .A2(n758), .ZN(n541) );
  XNOR2_X2 U400 ( .A(n399), .B(KEYINPUT35), .ZN(n755) );
  XNOR2_X2 U401 ( .A(n514), .B(n457), .ZN(n736) );
  XNOR2_X2 U402 ( .A(n456), .B(n455), .ZN(n514) );
  BUF_X2 U403 ( .A(n663), .Z(n362) );
  NOR2_X1 U404 ( .A1(n759), .A2(n757), .ZN(n585) );
  XNOR2_X1 U405 ( .A(KEYINPUT15), .B(G902), .ZN(n627) );
  NOR2_X1 U406 ( .A1(n525), .A2(n565), .ZN(n699) );
  NAND2_X1 U407 ( .A1(n599), .A2(n656), .ZN(n567) );
  NOR2_X1 U408 ( .A1(n650), .A2(n649), .ZN(n526) );
  NOR2_X1 U409 ( .A1(n733), .A2(n627), .ZN(n626) );
  XNOR2_X1 U410 ( .A(n558), .B(n557), .ZN(n733) );
  NOR2_X1 U411 ( .A1(n384), .A2(n699), .ZN(n556) );
  XNOR2_X1 U412 ( .A(n396), .B(KEYINPUT70), .ZN(n555) );
  XNOR2_X1 U413 ( .A(n709), .B(KEYINPUT83), .ZN(n408) );
  XNOR2_X1 U414 ( .A(n415), .B(n584), .ZN(n759) );
  XNOR2_X1 U415 ( .A(n413), .B(n372), .ZN(n540) );
  NOR2_X1 U416 ( .A1(n577), .A2(n576), .ZN(n580) );
  XNOR2_X1 U417 ( .A(n737), .B(n509), .ZN(n520) );
  XNOR2_X1 U418 ( .A(G107), .B(n368), .ZN(n737) );
  INV_X1 U419 ( .A(KEYINPUT3), .ZN(n453) );
  XOR2_X1 U420 ( .A(G143), .B(G128), .Z(n480) );
  XNOR2_X1 U421 ( .A(n363), .B(KEYINPUT122), .ZN(n684) );
  AND2_X1 U422 ( .A1(n683), .A2(n682), .ZN(n363) );
  NOR2_X1 U423 ( .A1(n755), .A2(n758), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n568), .B(n523), .ZN(n650) );
  INV_X1 U425 ( .A(n641), .ZN(n365) );
  INV_X1 U426 ( .A(n379), .ZN(n366) );
  INV_X1 U427 ( .A(n366), .ZN(n367) );
  XNOR2_X2 U428 ( .A(n499), .B(n498), .ZN(n515) );
  XNOR2_X2 U429 ( .A(KEYINPUT66), .B(G131), .ZN(n499) );
  XNOR2_X1 U430 ( .A(n395), .B(n465), .ZN(n697) );
  XNOR2_X2 U431 ( .A(n746), .B(n432), .ZN(n522) );
  XNOR2_X2 U432 ( .A(n433), .B(n516), .ZN(n746) );
  XNOR2_X1 U433 ( .A(n450), .B(n449), .ZN(n646) );
  OR2_X1 U434 ( .A1(n726), .A2(G902), .ZN(n450) );
  INV_X1 U435 ( .A(G146), .ZN(n432) );
  NOR2_X1 U436 ( .A1(n425), .A2(n421), .ZN(n420) );
  NAND2_X1 U437 ( .A1(n624), .A2(n424), .ZN(n421) );
  INV_X1 U438 ( .A(KEYINPUT44), .ZN(n397) );
  XNOR2_X1 U439 ( .A(G128), .B(G110), .ZN(n442) );
  XNOR2_X1 U440 ( .A(n480), .B(n479), .ZN(n516) );
  INV_X1 U441 ( .A(G134), .ZN(n479) );
  XNOR2_X1 U442 ( .A(n359), .B(G143), .ZN(n491) );
  XNOR2_X1 U443 ( .A(n736), .B(n459), .ZN(n395) );
  XNOR2_X1 U444 ( .A(n407), .B(n406), .ZN(n405) );
  INV_X1 U445 ( .A(KEYINPUT90), .ZN(n406) );
  NAND2_X1 U446 ( .A1(n540), .A2(n600), .ZN(n407) );
  XNOR2_X1 U447 ( .A(n412), .B(n410), .ZN(n726) );
  XNOR2_X1 U448 ( .A(n411), .B(n439), .ZN(n410) );
  XNOR2_X1 U449 ( .A(n444), .B(n744), .ZN(n412) );
  XNOR2_X1 U450 ( .A(n522), .B(n430), .ZN(n720) );
  XNOR2_X1 U451 ( .A(n520), .B(n431), .ZN(n430) );
  XNOR2_X1 U452 ( .A(n521), .B(G140), .ZN(n431) );
  XNOR2_X1 U453 ( .A(n445), .B(KEYINPUT20), .ZN(n451) );
  NAND2_X1 U454 ( .A1(G234), .A2(G237), .ZN(n471) );
  INV_X1 U455 ( .A(KEYINPUT67), .ZN(n498) );
  XNOR2_X1 U456 ( .A(n394), .B(KEYINPUT4), .ZN(n509) );
  XNOR2_X1 U457 ( .A(G101), .B(KEYINPUT65), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n515), .B(G137), .ZN(n433) );
  XOR2_X1 U459 ( .A(KEYINPUT18), .B(KEYINPUT80), .Z(n461) );
  NAND2_X1 U460 ( .A1(n423), .A2(KEYINPUT86), .ZN(n422) );
  OR2_X1 U461 ( .A1(n425), .A2(n717), .ZN(n423) );
  NOR2_X1 U462 ( .A1(G237), .A2(G902), .ZN(n466) );
  INV_X1 U463 ( .A(KEYINPUT113), .ZN(n574) );
  OR2_X2 U464 ( .A1(n720), .A2(G902), .ZN(n402) );
  NAND2_X1 U465 ( .A1(n646), .A2(n647), .ZN(n649) );
  NOR2_X1 U466 ( .A1(G237), .A2(G953), .ZN(n500) );
  XNOR2_X1 U467 ( .A(n509), .B(n393), .ZN(n512) );
  INV_X1 U468 ( .A(KEYINPUT5), .ZN(n393) );
  XNOR2_X1 U469 ( .A(KEYINPUT16), .B(G122), .ZN(n457) );
  XNOR2_X1 U470 ( .A(n462), .B(n440), .ZN(n744) );
  XNOR2_X1 U471 ( .A(n443), .B(n438), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U473 ( .A(KEYINPUT79), .ZN(n441) );
  XNOR2_X1 U474 ( .A(G116), .B(G107), .ZN(n481) );
  NAND2_X1 U475 ( .A1(n468), .A2(G214), .ZN(n662) );
  XNOR2_X1 U476 ( .A(n527), .B(KEYINPUT33), .ZN(n528) );
  INV_X1 U477 ( .A(KEYINPUT95), .ZN(n527) );
  AND2_X1 U478 ( .A1(n570), .A2(n647), .ZN(n414) );
  INV_X1 U479 ( .A(G125), .ZN(n687) );
  AND2_X1 U480 ( .A1(n409), .A2(n598), .ZN(n709) );
  XNOR2_X1 U481 ( .A(n404), .B(n403), .ZN(n525) );
  INV_X1 U482 ( .A(KEYINPUT91), .ZN(n403) );
  XNOR2_X1 U483 ( .A(n728), .B(n727), .ZN(n380) );
  XNOR2_X1 U484 ( .A(n724), .B(n723), .ZN(n382) );
  INV_X1 U485 ( .A(KEYINPUT60), .ZN(n385) );
  XNOR2_X1 U486 ( .A(n722), .B(n721), .ZN(n381) );
  INV_X1 U487 ( .A(KEYINPUT56), .ZN(n387) );
  XOR2_X1 U488 ( .A(G104), .B(G110), .Z(n368) );
  AND2_X1 U489 ( .A1(n426), .A2(n624), .ZN(n369) );
  AND2_X1 U490 ( .A1(n704), .A2(n397), .ZN(n371) );
  XOR2_X1 U491 ( .A(KEYINPUT72), .B(KEYINPUT22), .Z(n372) );
  XOR2_X1 U492 ( .A(KEYINPUT94), .B(KEYINPUT0), .Z(n373) );
  XOR2_X1 U493 ( .A(n636), .B(KEYINPUT62), .Z(n374) );
  XOR2_X1 U494 ( .A(n694), .B(n693), .Z(n375) );
  XOR2_X1 U495 ( .A(n697), .B(n696), .Z(n376) );
  INV_X1 U496 ( .A(KEYINPUT86), .ZN(n424) );
  INV_X1 U497 ( .A(n729), .ZN(n389) );
  INV_X1 U498 ( .A(n608), .ZN(n524) );
  BUF_X1 U499 ( .A(n678), .Z(n377) );
  AND2_X1 U500 ( .A1(n419), .A2(n418), .ZN(n378) );
  NAND2_X1 U501 ( .A1(n416), .A2(KEYINPUT86), .ZN(n418) );
  NOR2_X1 U502 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X2 U503 ( .A1(n419), .A2(n418), .ZN(n747) );
  INV_X1 U504 ( .A(n379), .ZN(n530) );
  NAND2_X1 U505 ( .A1(n379), .A2(n414), .ZN(n413) );
  XNOR2_X2 U506 ( .A(n478), .B(n373), .ZN(n379) );
  NAND2_X1 U507 ( .A1(n367), .A2(n658), .ZN(n549) );
  NOR2_X1 U508 ( .A1(n380), .A2(n729), .ZN(G66) );
  NOR2_X1 U509 ( .A1(n381), .A2(n729), .ZN(G54) );
  NOR2_X1 U510 ( .A1(n382), .A2(n729), .ZN(G63) );
  NAND2_X1 U511 ( .A1(n554), .A2(n553), .ZN(n384) );
  XNOR2_X1 U512 ( .A(n386), .B(n385), .ZN(G60) );
  NAND2_X1 U513 ( .A1(n391), .A2(n389), .ZN(n386) );
  XNOR2_X1 U514 ( .A(n388), .B(n387), .ZN(G51) );
  NAND2_X1 U515 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U516 ( .A(n583), .B(n582), .ZN(n392) );
  XNOR2_X1 U517 ( .A(n698), .B(n376), .ZN(n390) );
  XNOR2_X1 U518 ( .A(n695), .B(n375), .ZN(n391) );
  NAND2_X1 U519 ( .A1(n392), .A2(n690), .ZN(n415) );
  NAND2_X1 U520 ( .A1(n392), .A2(n705), .ZN(n716) );
  NAND2_X1 U521 ( .A1(n541), .A2(n704), .ZN(n398) );
  NAND2_X1 U522 ( .A1(n364), .A2(n371), .ZN(n396) );
  NAND2_X1 U523 ( .A1(n398), .A2(KEYINPUT44), .ZN(n554) );
  NAND2_X1 U524 ( .A1(n400), .A2(n598), .ZN(n399) );
  XNOR2_X1 U525 ( .A(n401), .B(KEYINPUT34), .ZN(n400) );
  XNOR2_X2 U526 ( .A(n402), .B(G469), .ZN(n568) );
  NAND2_X1 U527 ( .A1(n405), .A2(n524), .ZN(n404) );
  NAND2_X1 U528 ( .A1(n370), .A2(n408), .ZN(n611) );
  XNOR2_X1 U529 ( .A(n597), .B(KEYINPUT114), .ZN(n409) );
  INV_X1 U530 ( .A(n649), .ZN(n544) );
  INV_X1 U531 ( .A(n646), .ZN(n565) );
  NAND2_X1 U532 ( .A1(n556), .A2(n555), .ZN(n558) );
  INV_X1 U533 ( .A(n426), .ZN(n416) );
  XNOR2_X2 U534 ( .A(n617), .B(n616), .ZN(n426) );
  NAND2_X1 U535 ( .A1(n426), .A2(n420), .ZN(n417) );
  INV_X1 U536 ( .A(n716), .ZN(n425) );
  NAND2_X1 U537 ( .A1(n428), .A2(n590), .ZN(n427) );
  NAND2_X1 U538 ( .A1(n594), .A2(n429), .ZN(n428) );
  AND2_X1 U539 ( .A1(n667), .A2(KEYINPUT82), .ZN(n429) );
  NAND2_X1 U540 ( .A1(n571), .A2(n662), .ZN(n469) );
  NAND2_X1 U541 ( .A1(n544), .A2(n568), .ZN(n575) );
  XNOR2_X1 U542 ( .A(n726), .B(KEYINPUT124), .ZN(n727) );
  AND2_X1 U543 ( .A1(n468), .A2(G210), .ZN(n434) );
  XNOR2_X1 U544 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U545 ( .A(n686), .B(n685), .ZN(G75) );
  NAND2_X1 U546 ( .A1(G234), .A2(n748), .ZN(n435) );
  XOR2_X1 U547 ( .A(KEYINPUT8), .B(n435), .Z(n484) );
  NAND2_X1 U548 ( .A1(n484), .A2(G221), .ZN(n444) );
  XOR2_X1 U549 ( .A(KEYINPUT23), .B(KEYINPUT101), .Z(n437) );
  XNOR2_X1 U550 ( .A(G119), .B(G137), .ZN(n436) );
  XNOR2_X1 U551 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U552 ( .A(KEYINPUT24), .B(KEYINPUT84), .Z(n438) );
  XNOR2_X1 U553 ( .A(n687), .B(G146), .ZN(n462) );
  XNOR2_X1 U554 ( .A(KEYINPUT10), .B(G140), .ZN(n440) );
  XOR2_X1 U555 ( .A(KEYINPUT102), .B(KEYINPUT78), .Z(n447) );
  NAND2_X1 U556 ( .A1(n627), .A2(G234), .ZN(n445) );
  NAND2_X1 U557 ( .A1(G217), .A2(n451), .ZN(n446) );
  XNOR2_X1 U558 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U559 ( .A(KEYINPUT25), .B(n448), .ZN(n449) );
  NAND2_X1 U560 ( .A1(n451), .A2(G221), .ZN(n452) );
  XNOR2_X1 U561 ( .A(KEYINPUT21), .B(n452), .ZN(n563) );
  XNOR2_X2 U562 ( .A(G116), .B(G113), .ZN(n454) );
  XOR2_X1 U563 ( .A(G119), .B(KEYINPUT69), .Z(n455) );
  XOR2_X1 U564 ( .A(KEYINPUT17), .B(KEYINPUT96), .Z(n458) );
  XNOR2_X1 U565 ( .A(n480), .B(n458), .ZN(n459) );
  NAND2_X1 U566 ( .A1(G224), .A2(n748), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n461), .B(n460), .ZN(n463) );
  XNOR2_X1 U568 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n520), .B(n464), .ZN(n465) );
  NAND2_X1 U570 ( .A1(n697), .A2(n627), .ZN(n467) );
  XOR2_X1 U571 ( .A(KEYINPUT74), .B(n466), .Z(n468) );
  XNOR2_X2 U572 ( .A(n467), .B(n434), .ZN(n571) );
  XNOR2_X2 U573 ( .A(n469), .B(KEYINPUT93), .ZN(n603) );
  XNOR2_X1 U574 ( .A(KEYINPUT19), .B(KEYINPUT77), .ZN(n470) );
  XNOR2_X1 U575 ( .A(n471), .B(KEYINPUT14), .ZN(n473) );
  NAND2_X1 U576 ( .A1(n473), .A2(G952), .ZN(n472) );
  XOR2_X1 U577 ( .A(KEYINPUT97), .B(n472), .Z(n677) );
  NOR2_X1 U578 ( .A1(G953), .A2(n677), .ZN(n562) );
  NAND2_X1 U579 ( .A1(n473), .A2(G902), .ZN(n474) );
  XOR2_X1 U580 ( .A(KEYINPUT99), .B(n474), .Z(n559) );
  XOR2_X1 U581 ( .A(G898), .B(KEYINPUT98), .Z(n732) );
  NAND2_X1 U582 ( .A1(G953), .A2(n732), .ZN(n740) );
  NOR2_X1 U583 ( .A1(n559), .A2(n740), .ZN(n475) );
  NOR2_X1 U584 ( .A1(n562), .A2(n475), .ZN(n476) );
  XOR2_X1 U585 ( .A(KEYINPUT100), .B(n476), .Z(n477) );
  NAND2_X1 U586 ( .A1(n477), .A2(n586), .ZN(n478) );
  XOR2_X1 U587 ( .A(KEYINPUT109), .B(G122), .Z(n482) );
  XNOR2_X1 U588 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U589 ( .A(n516), .B(n483), .Z(n486) );
  NAND2_X1 U590 ( .A1(G217), .A2(n484), .ZN(n485) );
  XNOR2_X1 U591 ( .A(n486), .B(n485), .ZN(n488) );
  XOR2_X1 U592 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n487) );
  XNOR2_X1 U593 ( .A(n488), .B(n487), .ZN(n723) );
  NOR2_X1 U594 ( .A1(n723), .A2(G902), .ZN(n489) );
  XNOR2_X1 U595 ( .A(n489), .B(G478), .ZN(n543) );
  INV_X1 U596 ( .A(n543), .ZN(n508) );
  XNOR2_X1 U597 ( .A(G104), .B(KEYINPUT106), .ZN(n490) );
  XNOR2_X1 U598 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U599 ( .A(n744), .B(n492), .ZN(n497) );
  XNOR2_X1 U600 ( .A(KEYINPUT11), .B(G122), .ZN(n493) );
  XNOR2_X1 U601 ( .A(n493), .B(KEYINPUT12), .ZN(n495) );
  XNOR2_X1 U602 ( .A(KEYINPUT105), .B(KEYINPUT107), .ZN(n494) );
  XNOR2_X1 U603 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U604 ( .A(n497), .B(n496), .ZN(n503) );
  XNOR2_X1 U605 ( .A(n500), .B(KEYINPUT76), .ZN(n510) );
  NAND2_X1 U606 ( .A1(n510), .A2(G214), .ZN(n501) );
  XNOR2_X1 U607 ( .A(n515), .B(n501), .ZN(n502) );
  XNOR2_X1 U608 ( .A(n503), .B(n502), .ZN(n694) );
  OR2_X1 U609 ( .A1(n694), .A2(G902), .ZN(n507) );
  XNOR2_X1 U610 ( .A(G475), .B(KEYINPUT13), .ZN(n505) );
  INV_X1 U611 ( .A(KEYINPUT108), .ZN(n504) );
  XNOR2_X1 U612 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U613 ( .A(n507), .B(n506), .ZN(n542) );
  NOR2_X1 U614 ( .A1(n508), .A2(n542), .ZN(n570) );
  NAND2_X1 U615 ( .A1(G210), .A2(n510), .ZN(n511) );
  XNOR2_X1 U616 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U617 ( .A(n514), .B(n513), .ZN(n517) );
  XNOR2_X1 U618 ( .A(n522), .B(n517), .ZN(n636) );
  NOR2_X1 U619 ( .A1(G902), .A2(n636), .ZN(n519) );
  XNOR2_X1 U620 ( .A(G472), .B(KEYINPUT71), .ZN(n518) );
  XNOR2_X2 U621 ( .A(n519), .B(n518), .ZN(n656) );
  XNOR2_X1 U622 ( .A(n656), .B(KEYINPUT6), .ZN(n600) );
  NAND2_X1 U623 ( .A1(G227), .A2(n748), .ZN(n521) );
  INV_X1 U624 ( .A(KEYINPUT1), .ZN(n523) );
  INV_X1 U625 ( .A(n650), .ZN(n608) );
  INV_X1 U626 ( .A(n563), .ZN(n647) );
  XNOR2_X1 U627 ( .A(n526), .B(KEYINPUT73), .ZN(n547) );
  NOR2_X1 U628 ( .A1(n547), .A2(n600), .ZN(n529) );
  XNOR2_X1 U629 ( .A(n529), .B(n528), .ZN(n678) );
  INV_X1 U630 ( .A(n542), .ZN(n531) );
  OR2_X1 U631 ( .A1(n543), .A2(n531), .ZN(n533) );
  INV_X1 U632 ( .A(KEYINPUT112), .ZN(n532) );
  XNOR2_X1 U633 ( .A(n533), .B(n532), .ZN(n598) );
  NAND2_X1 U634 ( .A1(n565), .A2(n608), .ZN(n534) );
  XNOR2_X1 U635 ( .A(KEYINPUT111), .B(n534), .ZN(n535) );
  AND2_X1 U636 ( .A1(n535), .A2(n600), .ZN(n536) );
  NAND2_X1 U637 ( .A1(n565), .A2(n524), .ZN(n538) );
  NOR2_X1 U638 ( .A1(n656), .A2(n538), .ZN(n539) );
  NAND2_X1 U639 ( .A1(n540), .A2(n539), .ZN(n704) );
  AND2_X1 U640 ( .A1(n543), .A2(n542), .ZN(n690) );
  INV_X1 U641 ( .A(n690), .ZN(n710) );
  OR2_X1 U642 ( .A1(n543), .A2(n542), .ZN(n713) );
  NAND2_X1 U643 ( .A1(n710), .A2(n713), .ZN(n667) );
  NOR2_X1 U644 ( .A1(n656), .A2(n575), .ZN(n545) );
  XOR2_X1 U645 ( .A(KEYINPUT103), .B(n546), .Z(n700) );
  XOR2_X1 U646 ( .A(KEYINPUT31), .B(KEYINPUT104), .Z(n550) );
  INV_X1 U647 ( .A(n656), .ZN(n548) );
  NOR2_X1 U648 ( .A1(n548), .A2(n547), .ZN(n658) );
  XNOR2_X1 U649 ( .A(n550), .B(n549), .ZN(n714) );
  XNOR2_X1 U650 ( .A(n552), .B(KEYINPUT110), .ZN(n553) );
  INV_X1 U651 ( .A(KEYINPUT45), .ZN(n557) );
  OR2_X1 U652 ( .A1(n748), .A2(n559), .ZN(n560) );
  NOR2_X1 U653 ( .A1(G900), .A2(n560), .ZN(n561) );
  NOR2_X1 U654 ( .A1(n562), .A2(n561), .ZN(n577) );
  NOR2_X1 U655 ( .A1(n563), .A2(n577), .ZN(n564) );
  AND2_X1 U656 ( .A1(n565), .A2(n564), .ZN(n599) );
  XNOR2_X1 U657 ( .A(KEYINPUT28), .B(KEYINPUT115), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n567), .B(n566), .ZN(n569) );
  NAND2_X1 U659 ( .A1(n569), .A2(n568), .ZN(n588) );
  INV_X1 U660 ( .A(n570), .ZN(n665) );
  XOR2_X1 U661 ( .A(n571), .B(KEYINPUT38), .Z(n663) );
  NAND2_X1 U662 ( .A1(n362), .A2(n662), .ZN(n668) );
  NOR2_X1 U663 ( .A1(n665), .A2(n668), .ZN(n572) );
  XNOR2_X1 U664 ( .A(n572), .B(KEYINPUT41), .ZN(n679) );
  NOR2_X1 U665 ( .A1(n588), .A2(n679), .ZN(n573) );
  XNOR2_X1 U666 ( .A(n573), .B(KEYINPUT42), .ZN(n757) );
  NAND2_X1 U667 ( .A1(n656), .A2(n662), .ZN(n578) );
  XOR2_X1 U668 ( .A(KEYINPUT30), .B(n578), .Z(n579) );
  NAND2_X1 U669 ( .A1(n580), .A2(n579), .ZN(n596) );
  INV_X1 U670 ( .A(n362), .ZN(n581) );
  INV_X1 U671 ( .A(KEYINPUT39), .ZN(n582) );
  INV_X1 U672 ( .A(KEYINPUT40), .ZN(n584) );
  XNOR2_X1 U673 ( .A(n585), .B(KEYINPUT46), .ZN(n613) );
  XNOR2_X1 U674 ( .A(n706), .B(KEYINPUT47), .ZN(n594) );
  AND2_X1 U675 ( .A1(KEYINPUT82), .A2(KEYINPUT47), .ZN(n589) );
  OR2_X1 U676 ( .A1(n667), .A2(n589), .ZN(n590) );
  INV_X1 U677 ( .A(KEYINPUT47), .ZN(n592) );
  INV_X1 U678 ( .A(KEYINPUT82), .ZN(n591) );
  NAND2_X1 U679 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U680 ( .A1(n706), .A2(n594), .ZN(n595) );
  INV_X1 U681 ( .A(n571), .ZN(n622) );
  NOR2_X1 U682 ( .A1(n596), .A2(n622), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n599), .A2(n690), .ZN(n601) );
  OR2_X1 U684 ( .A1(n601), .A2(n600), .ZN(n618) );
  INV_X1 U685 ( .A(KEYINPUT116), .ZN(n602) );
  XNOR2_X1 U686 ( .A(n618), .B(n602), .ZN(n604) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n607) );
  XNOR2_X1 U688 ( .A(KEYINPUT117), .B(KEYINPUT36), .ZN(n605) );
  XNOR2_X1 U689 ( .A(n605), .B(KEYINPUT92), .ZN(n606) );
  XNOR2_X1 U690 ( .A(n607), .B(n606), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n689) );
  XNOR2_X1 U692 ( .A(n689), .B(KEYINPUT89), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n617) );
  XNOR2_X1 U694 ( .A(KEYINPUT88), .B(KEYINPUT48), .ZN(n615) );
  INV_X1 U695 ( .A(KEYINPUT68), .ZN(n614) );
  XNOR2_X1 U696 ( .A(n615), .B(n614), .ZN(n616) );
  INV_X1 U697 ( .A(n618), .ZN(n620) );
  AND2_X1 U698 ( .A1(n524), .A2(n662), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n621), .B(KEYINPUT43), .ZN(n623) );
  AND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n717) );
  INV_X1 U702 ( .A(n717), .ZN(n624) );
  INV_X1 U703 ( .A(n713), .ZN(n705) );
  XNOR2_X1 U704 ( .A(n747), .B(KEYINPUT75), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n630) );
  XNOR2_X1 U706 ( .A(n627), .B(KEYINPUT85), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n628), .A2(KEYINPUT2), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n635) );
  INV_X1 U709 ( .A(n733), .ZN(n641) );
  NAND2_X1 U710 ( .A1(KEYINPUT2), .A2(n716), .ZN(n631) );
  XNOR2_X1 U711 ( .A(KEYINPUT81), .B(n631), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n369), .A2(n632), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n633), .B(KEYINPUT87), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n641), .A2(n634), .ZN(n644) );
  AND2_X2 U715 ( .A1(n635), .A2(n644), .ZN(n718) );
  NAND2_X1 U716 ( .A1(n718), .A2(G472), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n637), .B(n374), .ZN(n639) );
  INV_X1 U718 ( .A(G952), .ZN(n638) );
  AND2_X1 U719 ( .A1(n638), .A2(G953), .ZN(n729) );
  NAND2_X1 U720 ( .A1(n639), .A2(n389), .ZN(n640) );
  XNOR2_X1 U721 ( .A(n640), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U722 ( .A1(n641), .A2(n378), .ZN(n643) );
  INV_X1 U723 ( .A(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n683) );
  NOR2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U727 ( .A(KEYINPUT49), .B(n648), .ZN(n654) );
  XOR2_X1 U728 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n652) );
  NAND2_X1 U729 ( .A1(n524), .A2(n649), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U734 ( .A(KEYINPUT51), .B(n659), .Z(n660) );
  NOR2_X1 U735 ( .A1(n679), .A2(n660), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(KEYINPUT120), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n362), .A2(n662), .ZN(n664) );
  XOR2_X1 U738 ( .A(KEYINPUT121), .B(n664), .Z(n666) );
  NOR2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n671) );
  INV_X1 U740 ( .A(n667), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U743 ( .A1(n377), .A2(n672), .ZN(n673) );
  NOR2_X1 U744 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U745 ( .A(n675), .B(KEYINPUT52), .ZN(n676) );
  NOR2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n679), .A2(n377), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n748), .A2(n684), .ZN(n686) );
  XNOR2_X1 U750 ( .A(KEYINPUT53), .B(KEYINPUT123), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n687), .B(KEYINPUT37), .ZN(n688) );
  XNOR2_X1 U752 ( .A(n689), .B(n688), .ZN(G27) );
  NAND2_X1 U753 ( .A1(n706), .A2(n690), .ZN(n691) );
  XNOR2_X1 U754 ( .A(n691), .B(G146), .ZN(G48) );
  NOR2_X1 U755 ( .A1(n700), .A2(n710), .ZN(n692) );
  XOR2_X1 U756 ( .A(n692), .B(G104), .Z(G6) );
  NAND2_X1 U757 ( .A1(n718), .A2(G475), .ZN(n695) );
  XOR2_X1 U758 ( .A(KEYINPUT64), .B(KEYINPUT59), .Z(n693) );
  NAND2_X1 U759 ( .A1(n718), .A2(G210), .ZN(n698) );
  XNOR2_X1 U760 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n696) );
  XOR2_X1 U761 ( .A(n699), .B(G101), .Z(G3) );
  NOR2_X1 U762 ( .A1(n700), .A2(n713), .ZN(n702) );
  XNOR2_X1 U763 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n701) );
  XNOR2_X1 U764 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U765 ( .A(G107), .B(n703), .ZN(G9) );
  XNOR2_X1 U766 ( .A(G110), .B(n704), .ZN(G12) );
  XOR2_X1 U767 ( .A(G128), .B(KEYINPUT29), .Z(n708) );
  NAND2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U769 ( .A(n708), .B(n707), .ZN(G30) );
  XOR2_X1 U770 ( .A(G143), .B(n709), .Z(G45) );
  NOR2_X1 U771 ( .A1(n714), .A2(n710), .ZN(n711) );
  XOR2_X1 U772 ( .A(KEYINPUT118), .B(n711), .Z(n712) );
  XNOR2_X1 U773 ( .A(n359), .B(n712), .ZN(G15) );
  NOR2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U775 ( .A(G116), .B(n715), .Z(G18) );
  XNOR2_X1 U776 ( .A(G134), .B(n716), .ZN(G36) );
  XOR2_X1 U777 ( .A(G140), .B(n717), .Z(G42) );
  NAND2_X1 U778 ( .A1(n725), .A2(G469), .ZN(n722) );
  XOR2_X1 U779 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n719) );
  XNOR2_X1 U780 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U781 ( .A1(n725), .A2(G478), .ZN(n724) );
  NAND2_X1 U782 ( .A1(n725), .A2(G217), .ZN(n728) );
  NAND2_X1 U783 ( .A1(G953), .A2(G224), .ZN(n730) );
  XOR2_X1 U784 ( .A(KEYINPUT61), .B(n730), .Z(n731) );
  NOR2_X1 U785 ( .A1(n732), .A2(n731), .ZN(n735) );
  NOR2_X1 U786 ( .A1(G953), .A2(n365), .ZN(n734) );
  NOR2_X1 U787 ( .A1(n735), .A2(n734), .ZN(n743) );
  XNOR2_X1 U788 ( .A(n736), .B(KEYINPUT125), .ZN(n738) );
  XNOR2_X1 U789 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U790 ( .A(n739), .B(G101), .ZN(n741) );
  NAND2_X1 U791 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(G69) );
  XNOR2_X1 U793 ( .A(n744), .B(KEYINPUT4), .ZN(n745) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(n750) );
  XNOR2_X1 U795 ( .A(n747), .B(n750), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(n754) );
  XNOR2_X1 U797 ( .A(G227), .B(n750), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U799 ( .A1(G953), .A2(n752), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n754), .A2(n753), .ZN(G72) );
  XOR2_X1 U801 ( .A(n755), .B(G122), .Z(G24) );
  XOR2_X1 U802 ( .A(G137), .B(KEYINPUT126), .Z(n756) );
  XNOR2_X1 U803 ( .A(n757), .B(n756), .ZN(G39) );
  XOR2_X1 U804 ( .A(n758), .B(G119), .Z(G21) );
  XOR2_X1 U805 ( .A(n759), .B(G131), .Z(G33) );
endmodule

