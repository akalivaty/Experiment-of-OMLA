//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n570, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT69), .Z(new_n455));
  OR2_X1    g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(KEYINPUT71), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(G567), .B2(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(KEYINPUT71), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  XNOR2_X1  g039(.A(KEYINPUT72), .B(G2105), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  AND2_X1   g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(KEYINPUT73), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT73), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT72), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT72), .A2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n475), .A2(G137), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT75), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n471), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT74), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(G101), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(G101), .A3(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT74), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n479), .A2(new_n480), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n469), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n480), .B1(new_n479), .B2(new_n487), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(G160));
  AND2_X1   g066(.A1(new_n472), .A2(new_n474), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G136), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT76), .Z(new_n495));
  NOR2_X1   g070(.A1(new_n492), .A2(new_n478), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G124), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT77), .ZN(new_n498));
  OAI221_X1 g073(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n478), .C2(G112), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT78), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n500), .B(new_n501), .ZN(G162));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  MUX2_X1   g078(.A(G102), .B(G114), .S(G2105), .Z(new_n504));
  AOI22_X1  g079(.A1(new_n475), .A2(new_n503), .B1(new_n504), .B2(G2104), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n465), .B1(new_n472), .B2(new_n474), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G138), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT79), .ZN(new_n509));
  INV_X1    g084(.A(G138), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n510), .A2(KEYINPUT4), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(new_n484), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT72), .A2(G2105), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n509), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n478), .A2(new_n466), .A3(KEYINPUT79), .A4(new_n511), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n505), .B1(new_n508), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g099(.A(KEYINPUT80), .B(new_n505), .C1(new_n508), .C2(new_n521), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(G164));
  XNOR2_X1  g102(.A(KEYINPUT5), .B(G543), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G50), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n530), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G166));
  AND2_X1   g113(.A1(new_n529), .A2(G89), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n528), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(KEYINPUT6), .A2(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(KEYINPUT6), .A2(G651), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n548));
  AOI22_X1  g123(.A1(G51), .A2(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n541), .A2(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  INV_X1    g126(.A(new_n530), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n552), .A2(G90), .B1(G52), .B2(new_n545), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n536), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  XNOR2_X1  g134(.A(KEYINPUT82), .B(G81), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n545), .A2(G43), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n536), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  XOR2_X1   g144(.A(KEYINPUT83), .B(KEYINPUT8), .Z(new_n570));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G188));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n532), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n545), .A2(new_n576), .A3(G53), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n528), .A2(G65), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n575), .A2(new_n577), .B1(new_n580), .B2(G651), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n530), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT84), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n583), .A2(G91), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G166), .ZN(G303));
  AND2_X1   g162(.A1(new_n583), .A2(new_n584), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G87), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n528), .A2(G74), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G49), .B2(new_n545), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n528), .A2(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G48), .B2(new_n545), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n583), .A2(G86), .A3(new_n584), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT85), .ZN(G305));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n530), .A2(new_n600), .B1(new_n532), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n536), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT86), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(new_n588), .A2(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n588), .A2(KEYINPUT10), .A3(G92), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n545), .A2(G54), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n528), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n536), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  MUX2_X1   g194(.A(G301), .B(new_n618), .S(new_n619), .Z(G284));
  MUX2_X1   g195(.A(G301), .B(new_n618), .S(new_n619), .Z(G321));
  NOR2_X1   g196(.A1(G286), .A2(new_n619), .ZN(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n619), .ZN(G280));
  XNOR2_X1  g199(.A(G280), .B(KEYINPUT88), .ZN(G297));
  AOI21_X1  g200(.A(new_n616), .B1(new_n611), .B2(new_n612), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  NOR3_X1   g203(.A1(new_n563), .A2(G868), .A3(new_n565), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n618), .A2(G559), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G323));
  XNOR2_X1  g206(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n632));
  XNOR2_X1  g207(.A(G323), .B(new_n632), .ZN(G282));
  NAND2_X1  g208(.A1(new_n466), .A2(new_n481), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(KEYINPUT90), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(KEYINPUT90), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n635), .A2(KEYINPUT13), .ZN(new_n640));
  OR3_X1    g215(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n639), .B1(new_n638), .B2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n493), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n496), .A2(G123), .ZN(new_n644));
  OAI221_X1 g219(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n478), .C2(G111), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n641), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT91), .ZN(G156));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT14), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT92), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n651), .B2(new_n652), .ZN(new_n656));
  XOR2_X1   g231(.A(G2451), .B(G2454), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n656), .B(new_n658), .Z(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n663), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT93), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n669), .B2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n670), .B2(new_n671), .ZN(new_n675));
  INV_X1    g250(.A(new_n671), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n676), .A2(new_n672), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n673), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2096), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2100), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n685), .A2(new_n686), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n684), .A2(new_n689), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n684), .A2(new_n689), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n692));
  AOI211_X1 g267(.A(new_n688), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(new_n691), .B2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(G1981), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT95), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT96), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n698), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  NAND3_X1  g279(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT25), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n493), .A2(G139), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n706), .B(new_n707), .C1(new_n478), .C2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G33), .B(new_n709), .S(G29), .Z(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G2072), .Z(new_n711));
  INV_X1    g286(.A(G2084), .ZN(new_n712));
  NAND2_X1  g287(.A1(G160), .A2(G29), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  AND2_X1   g289(.A1(KEYINPUT24), .A2(G34), .ZN(new_n715));
  NOR2_X1   g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n493), .A2(G141), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n496), .A2(G129), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT26), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n723), .A2(new_n724), .B1(G105), .B2(new_n481), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n719), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G32), .B(new_n726), .S(G29), .Z(new_n727));
  XOR2_X1   g302(.A(KEYINPUT27), .B(G1996), .Z(new_n728));
  OAI221_X1 g303(.A(new_n711), .B1(new_n712), .B2(new_n718), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n714), .A2(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n714), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2078), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n734), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1961), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G19), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n566), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1341), .ZN(new_n740));
  INV_X1    g315(.A(G1966), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT102), .B1(G16), .B2(G21), .ZN(new_n742));
  NOR2_X1   g317(.A1(G286), .A2(new_n734), .ZN(new_n743));
  MUX2_X1   g318(.A(new_n742), .B(KEYINPUT102), .S(new_n743), .Z(new_n744));
  AOI21_X1  g319(.A(new_n740), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n741), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n714), .A2(G26), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  OAI221_X1 g323(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n478), .C2(G116), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT100), .Z(new_n750));
  AOI22_X1  g325(.A1(G128), .A2(new_n496), .B1(new_n493), .B2(G140), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n748), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2067), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT31), .B(G11), .Z(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT30), .B(G28), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n755), .B1(new_n714), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n646), .B2(new_n714), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n727), .B2(new_n728), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n745), .A2(new_n746), .A3(new_n754), .A4(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G4), .A2(G16), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n626), .B2(G16), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G1348), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n718), .A2(new_n712), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n734), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT23), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1956), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n762), .B2(G1348), .ZN(new_n770));
  OR4_X1    g345(.A1(new_n737), .A2(new_n760), .A3(new_n765), .A4(new_n770), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n730), .A2(new_n733), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G29), .A2(G35), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G162), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT29), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G2090), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(G2090), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT103), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n772), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  MUX2_X1   g354(.A(G6), .B(G305), .S(G16), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT98), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT32), .B(G1981), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  MUX2_X1   g359(.A(G23), .B(G288), .S(G16), .Z(new_n785));
  XOR2_X1   g360(.A(KEYINPUT33), .B(G1976), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G22), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G166), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT99), .B(G1971), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n783), .A2(new_n784), .A3(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n795));
  MUX2_X1   g370(.A(G24), .B(G290), .S(G16), .Z(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(G1986), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(G1986), .ZN(new_n798));
  NOR2_X1   g373(.A1(G95), .A2(G2105), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT97), .Z(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G107), .C2(new_n478), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n496), .A2(G119), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n493), .A2(G131), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G25), .B(new_n804), .S(G29), .Z(new_n805));
  XOR2_X1   g380(.A(KEYINPUT35), .B(G1991), .Z(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n805), .B(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n797), .A2(new_n798), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n794), .A2(new_n795), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(KEYINPUT36), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n794), .A2(new_n812), .A3(new_n795), .A4(new_n809), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n779), .B1(new_n811), .B2(new_n813), .ZN(G311));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n813), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n815), .A2(new_n776), .A3(new_n772), .A4(new_n778), .ZN(G150));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  INV_X1    g392(.A(G55), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n530), .A2(new_n817), .B1(new_n532), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n536), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n566), .A2(KEYINPUT104), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT104), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n563), .B2(new_n565), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n823), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n824), .A2(new_n823), .A3(new_n826), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n618), .A2(new_n627), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n834));
  AOI21_X1  g409(.A(G860), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n823), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT37), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(G145));
  INV_X1    g414(.A(KEYINPUT106), .ZN(new_n840));
  XNOR2_X1  g415(.A(G162), .B(G160), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(new_n646), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n804), .B(new_n635), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n493), .A2(G142), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n496), .A2(G130), .ZN(new_n845));
  OAI221_X1 g420(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n478), .C2(G118), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n843), .B(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n752), .B(new_n522), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n709), .A2(KEYINPUT105), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n726), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n840), .B1(new_n842), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n841), .B(new_n646), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n853), .A3(KEYINPUT106), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT107), .B(G37), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n842), .B2(new_n854), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(KEYINPUT40), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT40), .B1(new_n858), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(G395));
  XNOR2_X1  g440(.A(G305), .B(G166), .ZN(new_n866));
  XNOR2_X1  g441(.A(G290), .B(G288), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT42), .Z(new_n869));
  INV_X1    g444(.A(KEYINPUT108), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n630), .B(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(new_n830), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n830), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT109), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n618), .A2(new_n874), .A3(new_n623), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT109), .B1(new_n626), .B2(G299), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n626), .A2(G299), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n872), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(KEYINPUT41), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n875), .A2(new_n876), .A3(new_n882), .A4(new_n877), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n872), .A2(new_n873), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n869), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT110), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n869), .B1(new_n884), .B2(new_n880), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(G868), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(G868), .B2(new_n822), .ZN(G295));
  OAI21_X1  g466(.A(new_n890), .B1(G868), .B2(new_n822), .ZN(G331));
  NAND2_X1  g467(.A1(new_n881), .A2(new_n883), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n555), .A2(G168), .A3(new_n557), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G168), .B1(new_n555), .B2(new_n557), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n828), .B(new_n829), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  INV_X1    g473(.A(new_n829), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n898), .B(new_n894), .C1(new_n899), .C2(new_n827), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n879), .A2(new_n897), .A3(new_n900), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n868), .A3(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n866), .B(new_n867), .Z(new_n905));
  AOI22_X1  g480(.A1(new_n881), .A2(new_n883), .B1(new_n897), .B2(new_n900), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n901), .A2(new_n878), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  AND4_X1   g484(.A1(KEYINPUT43), .A2(new_n904), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n904), .A2(new_n908), .A3(new_n859), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(KEYINPUT43), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT111), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(new_n918), .A3(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n904), .A2(new_n908), .A3(new_n911), .A4(new_n909), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n921), .A2(KEYINPUT44), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT112), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n912), .A2(new_n918), .A3(KEYINPUT43), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n918), .B1(new_n912), .B2(KEYINPUT43), .ZN(new_n925));
  OAI211_X1 g500(.A(KEYINPUT112), .B(new_n922), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n915), .B1(new_n923), .B2(new_n927), .ZN(G397));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n522), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n490), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(G40), .A3(new_n488), .A4(new_n469), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n752), .A2(G2067), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n752), .B(G2067), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT113), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n726), .B(G1996), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n804), .A2(new_n807), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n804), .B(new_n806), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n936), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n936), .A2(G1986), .A3(G290), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT48), .ZN(new_n947));
  OAI22_X1  g522(.A1(new_n936), .A2(new_n943), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n935), .B1(new_n939), .B2(new_n726), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT126), .Z(new_n950));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n951));
  OAI22_X1  g526(.A1(new_n936), .A2(G1996), .B1(KEYINPUT125), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(KEYINPUT125), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n952), .B(new_n953), .Z(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OR3_X1    g530(.A1(new_n950), .A2(KEYINPUT47), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT47), .B1(new_n950), .B2(new_n955), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n948), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n941), .A2(new_n944), .ZN(new_n959));
  XNOR2_X1  g534(.A(G290), .B(G1986), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n935), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1981), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n596), .A2(new_n597), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT115), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n596), .A2(new_n597), .A3(new_n965), .A4(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n552), .A2(G86), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n962), .B1(new_n596), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT49), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT49), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n972), .B(new_n969), .C1(new_n964), .C2(new_n966), .ZN(new_n973));
  INV_X1    g548(.A(G40), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n489), .A2(new_n974), .A3(new_n490), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n475), .A2(G138), .A3(new_n478), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT4), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n519), .A3(new_n520), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n978), .B2(new_n505), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(G8), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n971), .A2(new_n973), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n589), .A2(G1976), .A3(new_n591), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n980), .A2(G8), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT52), .ZN(new_n985));
  INV_X1    g560(.A(G1976), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT52), .B1(G288), .B2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(G8), .A3(new_n980), .A4(new_n983), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  INV_X1    g566(.A(new_n525), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT80), .B1(new_n978), .B2(new_n505), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT50), .B(new_n929), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n930), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n934), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G2090), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n934), .B1(new_n979), .B2(KEYINPUT45), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n524), .B2(new_n525), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1002));
  INV_X1    g577(.A(G1971), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n991), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  OAI211_X1 g581(.A(G303), .B(G8), .C1(new_n1006), .C2(KEYINPUT55), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(KEYINPUT55), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n990), .A2(new_n1005), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n981), .ZN(new_n1011));
  INV_X1    g586(.A(new_n967), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n967), .A2(new_n970), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n972), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n967), .A2(KEYINPUT49), .A3(new_n970), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G288), .A2(G1976), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1011), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g595(.A(KEYINPUT116), .B(new_n1012), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1010), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT63), .ZN(new_n1023));
  AOI211_X1 g598(.A(G2090), .B(new_n934), .C1(new_n994), .C2(new_n996), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n929), .B1(new_n992), .B2(new_n993), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n931), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1971), .B1(new_n1026), .B2(new_n1000), .ZN(new_n1027));
  OAI211_X1 g602(.A(G8), .B(new_n1009), .C1(new_n1024), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(new_n998), .A3(new_n975), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n991), .B1(new_n1031), .B2(new_n1004), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1028), .B(new_n990), .C1(new_n1032), .C2(new_n1009), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n994), .A2(new_n996), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(new_n712), .A3(new_n975), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT45), .B(new_n929), .C1(new_n992), .C2(new_n993), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n934), .B1(new_n930), .B2(new_n931), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n741), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1040), .A2(G8), .A3(G168), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1023), .B1(new_n1033), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1028), .A2(new_n990), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1041), .A2(new_n1023), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1022), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G299), .A2(KEYINPUT117), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n1052));
  NAND3_X1  g627(.A1(G299), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1056), .B(new_n1050), .C1(new_n581), .C2(new_n585), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT118), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1956), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n930), .A2(new_n995), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n1025), .B2(new_n995), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1060), .B1(new_n1062), .B2(new_n934), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT56), .B(G2072), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1000), .B(new_n1064), .C1(new_n1001), .C2(KEYINPUT45), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1059), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1059), .A3(new_n1065), .ZN(new_n1067));
  INV_X1    g642(.A(G1348), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1070), .B2(new_n934), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n980), .A2(G2067), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n618), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1066), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n618), .B(new_n1072), .C1(new_n997), .C2(G1348), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT60), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1956), .B1(new_n1030), .B2(new_n975), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1065), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(new_n1067), .A3(KEYINPUT61), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT61), .B1(new_n1082), .B2(new_n1067), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n618), .A2(KEYINPUT60), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1072), .B(new_n1086), .C1(new_n997), .C2(G1348), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n1088));
  INV_X1    g663(.A(G1996), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(new_n1000), .C1(new_n1001), .C2(KEYINPUT45), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT58), .B(G1341), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT119), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n980), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n566), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1088), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  AOI211_X1 g673(.A(KEYINPUT59), .B(new_n1096), .C1(new_n1090), .C2(new_n1093), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1087), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1085), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1075), .B1(new_n1084), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1031), .A2(new_n1004), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1009), .B1(new_n1103), .B2(G8), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1043), .A2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1106));
  NAND3_X1  g681(.A1(new_n522), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(G2078), .ZN(new_n1109));
  AND4_X1   g684(.A1(new_n932), .A2(new_n975), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G2078), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(new_n1000), .C1(new_n1001), .C2(KEYINPUT45), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1110), .B1(new_n1112), .B2(new_n1108), .ZN(new_n1113));
  INV_X1    g688(.A(G1961), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1070), .B2(new_n934), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1113), .A2(G301), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1109), .ZN(new_n1117));
  AOI211_X1 g692(.A(new_n1117), .B(new_n934), .C1(new_n930), .C2(new_n931), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1112), .A2(new_n1108), .B1(new_n1036), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(G301), .B1(new_n1119), .B2(new_n1115), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1106), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G171), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1119), .A2(G301), .A3(new_n1115), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(KEYINPUT54), .A3(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(G168), .A2(new_n991), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT51), .B1(new_n1126), .B2(KEYINPUT121), .ZN(new_n1127));
  OAI211_X1 g702(.A(G8), .B(new_n1127), .C1(new_n1040), .C2(G286), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1126), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1127), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n997), .A2(new_n712), .B1(new_n1038), .B2(new_n741), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1129), .B(new_n1130), .C1(new_n1131), .C2(new_n991), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1040), .A2(G8), .A3(G286), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1128), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1105), .A2(new_n1121), .A3(new_n1125), .A4(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1048), .B1(new_n1102), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1128), .A2(new_n1132), .A3(new_n1133), .A4(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n1105), .A3(new_n1120), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT123), .B1(new_n1134), .B2(KEYINPUT62), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1138), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT124), .B(new_n961), .C1(new_n1136), .C2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1140), .A2(new_n1105), .A3(new_n1120), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1134), .A2(KEYINPUT62), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(new_n1149), .A3(new_n1137), .ZN(new_n1150));
  AND4_X1   g725(.A1(new_n1134), .A2(new_n1105), .A3(new_n1121), .A4(new_n1125), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1080), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1153), .B2(new_n1066), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1087), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1107), .A2(new_n975), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1025), .B2(new_n931), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1157), .A2(new_n1089), .B1(new_n980), .B2(new_n1092), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT59), .B1(new_n1158), .B2(new_n1096), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1094), .A2(new_n1088), .A3(new_n1097), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1155), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1154), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1074), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1151), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1150), .A2(new_n1165), .A3(new_n1048), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT124), .B1(new_n1166), .B2(new_n961), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n958), .B1(new_n1145), .B2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g743(.A1(G227), .A2(new_n463), .ZN(new_n1170));
  OAI211_X1 g744(.A(new_n703), .B(new_n1170), .C1(new_n664), .C2(new_n666), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1171), .B1(new_n858), .B2(new_n861), .ZN(new_n1172));
  AND2_X1   g746(.A1(new_n1172), .A2(new_n913), .ZN(G308));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n913), .ZN(G225));
endmodule


