//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1166;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n459), .A2(KEYINPUT68), .B1(G567), .B2(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT69), .B(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G137), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  AND2_X1   g050(.A1(new_n464), .A2(KEYINPUT70), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(KEYINPUT70), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n467), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  INV_X1    g055(.A(new_n465), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n481), .B1(new_n476), .B2(new_n477), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n465), .C2(G112), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n480), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n467), .A2(KEYINPUT69), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n492), .B(new_n494), .C1(new_n470), .C2(new_n471), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n464), .A2(new_n465), .A3(new_n498), .A4(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n491), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT71), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(new_n506), .B1(new_n502), .B2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n508), .A2(new_n509), .B1(G75), .B2(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n507), .A2(KEYINPUT72), .A3(G62), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n501), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(G88), .B1(G50), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n519), .B1(new_n512), .B2(new_n513), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n518), .A2(G51), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(G89), .B2(new_n517), .ZN(G168));
  AOI22_X1  g103(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n501), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n515), .A2(G543), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n516), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(new_n518), .A2(G43), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n507), .A2(G81), .A3(new_n515), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT74), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT74), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n501), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G860), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT77), .Z(G188));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n507), .B2(G65), .ZN(new_n555));
  INV_X1    g130(.A(G91), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n555), .A2(new_n501), .B1(new_n516), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n515), .A2(new_n561), .A3(G53), .A4(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n558), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n560), .A2(new_n558), .A3(new_n562), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n557), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  OAI21_X1  g145(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n518), .A2(G49), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n516), .ZN(G288));
  AOI22_X1  g149(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n501), .ZN(new_n576));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  INV_X1    g152(.A(G48), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n516), .A2(new_n577), .B1(new_n578), .B2(new_n533), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AND2_X1   g156(.A1(new_n507), .A2(G60), .ZN(new_n582));
  AND2_X1   g157(.A1(G72), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT80), .ZN(new_n586));
  XNOR2_X1  g161(.A(KEYINPUT81), .B(G85), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n517), .A2(new_n587), .B1(G47), .B2(new_n518), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  XNOR2_X1  g165(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT83), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n592), .A2(new_n516), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n516), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n594), .A2(new_n595), .B1(G54), .B2(new_n518), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n501), .B1(new_n597), .B2(KEYINPUT84), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(KEYINPUT84), .B2(new_n597), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n590), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n590), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n566), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(G868), .B2(new_n566), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n600), .B1(new_n606), .B2(G860), .ZN(G148));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n543), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n596), .A2(new_n599), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n608), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g188(.A1(G123), .A2(new_n483), .B1(new_n479), .B2(G135), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT85), .ZN(new_n615));
  NOR3_X1   g190(.A1(new_n465), .A2(new_n615), .A3(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n465), .B2(G111), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n617), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n614), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT86), .B(G2096), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(G156));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2430), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT87), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT88), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n631), .B2(new_n629), .ZN(new_n635));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n635), .B(new_n636), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(new_n638), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n640), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(G14), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n644), .B1(new_n640), .B2(new_n642), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n627), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n640), .A2(new_n642), .ZN(new_n649));
  INV_X1    g224(.A(new_n644), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g226(.A1(new_n651), .A2(KEYINPUT89), .A3(G14), .A4(new_n645), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2100), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G1986), .ZN(new_n669));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  AND2_X1   g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT91), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n678), .A2(new_n674), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n681), .A2(new_n671), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n677), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT92), .ZN(new_n684));
  INV_X1    g259(.A(G1981), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(KEYINPUT92), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n669), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n691), .A2(G1986), .A3(new_n687), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT93), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  AND3_X1   g270(.A1(new_n690), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n690), .B2(new_n692), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n668), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n690), .A2(new_n692), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(new_n694), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n690), .A2(new_n692), .A3(new_n695), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(new_n667), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT97), .ZN(new_n706));
  MUX2_X1   g281(.A(G23), .B(G288), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT33), .Z(new_n708));
  INV_X1    g283(.A(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT95), .B(G16), .Z(new_n711));
  NOR2_X1   g286(.A1(G166), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G22), .B2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G1971), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G6), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n580), .B2(new_n716), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT96), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT32), .B(G1981), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n721), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n710), .A2(new_n715), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n713), .A2(new_n714), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n706), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n722), .A2(new_n723), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n708), .B(G1976), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n725), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n729), .A2(KEYINPUT97), .A3(new_n730), .A4(new_n715), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n726), .A2(new_n731), .A3(KEYINPUT34), .ZN(new_n732));
  INV_X1    g307(.A(new_n711), .ZN(new_n733));
  MUX2_X1   g308(.A(G24), .B(G290), .S(new_n733), .Z(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(G1986), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(KEYINPUT94), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(KEYINPUT94), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n479), .A2(G131), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n483), .A2(G119), .ZN(new_n742));
  OAI221_X1 g317(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n465), .C2(G107), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(new_n739), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT35), .B(G1991), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n735), .A2(KEYINPUT98), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G1986), .B2(new_n734), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n732), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(KEYINPUT34), .B1(new_n726), .B2(new_n731), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n705), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n726), .A2(new_n731), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT34), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n756), .A2(KEYINPUT36), .A3(new_n732), .A4(new_n750), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n733), .A2(G19), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n541), .B(KEYINPUT75), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n733), .ZN(new_n760));
  INV_X1    g335(.A(G1341), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n736), .A2(G33), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n464), .A2(G127), .ZN(new_n764));
  NAND2_X1  g339(.A1(G115), .A2(G2104), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT100), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n465), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n767), .B2(new_n766), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n479), .A2(G139), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT25), .Z(new_n772));
  NAND3_X1  g347(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n763), .B1(new_n773), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G2072), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT101), .Z(new_n777));
  NOR2_X1   g352(.A1(new_n739), .A2(G27), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G164), .B2(new_n739), .ZN(new_n779));
  INV_X1    g354(.A(G2078), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n716), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n716), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(G1961), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n774), .A2(new_n775), .B1(G1961), .B2(new_n783), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n777), .A2(new_n781), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n739), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G35), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT103), .Z(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n486), .B2(new_n739), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT29), .Z(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G2090), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n711), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT23), .Z(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G299), .B2(G16), .ZN(new_n795));
  INV_X1    g370(.A(G1956), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n786), .A2(new_n792), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n791), .A2(G2090), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT104), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT102), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND3_X1  g379(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT26), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n803), .A2(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G141), .ZN(new_n810));
  INV_X1    g385(.A(G129), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n809), .B1(new_n478), .B2(new_n810), .C1(new_n811), .C2(new_n482), .ZN(new_n812));
  MUX2_X1   g387(.A(G32), .B(new_n812), .S(G29), .Z(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT27), .B(G1996), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n716), .A2(G21), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G168), .B2(new_n716), .ZN(new_n817));
  INV_X1    g392(.A(G1966), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G28), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT30), .ZN(new_n821));
  AOI21_X1  g396(.A(G29), .B1(new_n820), .B2(KEYINPUT30), .ZN(new_n822));
  OR2_X1    g397(.A1(KEYINPUT31), .A2(G11), .ZN(new_n823));
  NAND2_X1  g398(.A1(KEYINPUT31), .A2(G11), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n619), .B2(new_n787), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT24), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(G34), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(G34), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n787), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G160), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n736), .ZN(new_n832));
  INV_X1    g407(.A(G2084), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n826), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n815), .A2(new_n819), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n787), .A2(G26), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT28), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n483), .A2(G128), .ZN(new_n839));
  OAI221_X1 g414(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n465), .C2(G116), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n479), .A2(G140), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n838), .B1(new_n843), .B2(G29), .ZN(new_n844));
  INV_X1    g419(.A(G2067), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(G4), .A2(G16), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT99), .Z(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n610), .B2(new_n716), .ZN(new_n849));
  INV_X1    g424(.A(G1348), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n836), .A2(new_n846), .A3(new_n851), .ZN(new_n852));
  AND4_X1   g427(.A1(new_n762), .A2(new_n798), .A3(new_n800), .A4(new_n852), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n753), .A2(new_n757), .A3(new_n853), .ZN(G311));
  NAND3_X1  g429(.A1(new_n753), .A2(new_n757), .A3(new_n853), .ZN(G150));
  AOI22_X1  g430(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n501), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  INV_X1    g433(.A(G55), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n516), .A2(new_n858), .B1(new_n859), .B2(new_n533), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n543), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n541), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n600), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g445(.A(G860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n861), .A2(new_n544), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(G145));
  XNOR2_X1  g450(.A(new_n619), .B(G160), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n497), .A2(new_n499), .ZN(new_n879));
  INV_X1    g454(.A(new_n491), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n843), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n843), .A2(new_n881), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n745), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n886), .A2(new_n744), .A3(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n773), .B(new_n812), .ZN(new_n889));
  OAI221_X1 g464(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n465), .C2(G118), .ZN(new_n890));
  INV_X1    g465(.A(G142), .ZN(new_n891));
  INV_X1    g466(.A(G130), .ZN(new_n892));
  OAI221_X1 g467(.A(new_n890), .B1(new_n478), .B2(new_n891), .C1(new_n892), .C2(new_n482), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n623), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n889), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n888), .A2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n878), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n877), .A3(new_n896), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g479(.A1(new_n759), .A2(new_n861), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n611), .B1(new_n905), .B2(new_n864), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n600), .A2(new_n566), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n610), .A2(G299), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n611), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n863), .A2(new_n910), .A3(new_n865), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n906), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n906), .A2(new_n911), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n906), .A2(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n906), .A2(new_n909), .A3(new_n911), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G166), .B(G290), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n580), .B(G288), .Z(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n917), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(new_n917), .B2(new_n923), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n862), .A2(new_n608), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(G295));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n931), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  INV_X1    g511(.A(new_n926), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n938));
  AOI21_X1  g513(.A(G168), .B1(new_n938), .B2(G301), .ZN(new_n939));
  NAND2_X1  g514(.A1(G171), .A2(KEYINPUT106), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n866), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(G168), .A2(KEYINPUT106), .A3(G171), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n940), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n863), .A2(new_n865), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n914), .A3(new_n915), .ZN(new_n947));
  INV_X1    g522(.A(new_n909), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n942), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n937), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n919), .B1(new_n945), .B2(new_n942), .ZN(new_n951));
  INV_X1    g526(.A(new_n949), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n926), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n953), .A3(new_n902), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n936), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(G397));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(G164), .B2(G1384), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G40), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n469), .A2(new_n965), .A3(new_n474), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT46), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n843), .A2(G2067), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n841), .A2(new_n845), .A3(new_n842), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n974), .B2(new_n812), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT127), .Z(new_n977));
  OR2_X1    g552(.A1(new_n977), .A2(KEYINPUT47), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(KEYINPUT47), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n812), .B(G1996), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n747), .A3(new_n745), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n967), .B1(new_n982), .B2(new_n973), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n744), .B(new_n747), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G290), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n968), .A3(new_n669), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n985), .A2(new_n968), .B1(KEYINPUT48), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n988), .A2(KEYINPUT48), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n978), .A2(new_n979), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(G288), .A2(new_n709), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(KEYINPUT107), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n881), .A2(new_n966), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(G8), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n998));
  AND2_X1   g573(.A1(G288), .A2(new_n709), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(G8), .A3(new_n996), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n996), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n994), .C1(KEYINPUT52), .C2(new_n999), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(KEYINPUT108), .B(G1981), .Z(new_n1007));
  NAND2_X1  g582(.A1(new_n580), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n685), .B2(new_n580), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1008), .B(KEYINPUT49), .C1(new_n685), .C2(new_n580), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n1004), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1006), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(G166), .B2(new_n1003), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT55), .B(G8), .C1(new_n514), .C2(new_n520), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n966), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n881), .A2(new_n995), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n962), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n881), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n881), .A2(new_n1024), .A3(new_n995), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1025), .A2(new_n966), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2090), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1023), .A2(new_n714), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(new_n1003), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1018), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1016), .B(new_n1017), .C1(new_n1029), .C2(new_n1003), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1014), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT63), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1022), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1022), .A2(new_n1035), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1021), .A3(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1038), .A2(new_n818), .B1(new_n1027), .B2(new_n833), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1039), .A2(new_n1003), .A3(G286), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1033), .A2(KEYINPUT112), .A3(new_n1034), .A4(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1004), .B(KEYINPUT109), .ZN(new_n1042));
  NOR2_X1   g617(.A1(G288), .A2(G1976), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1013), .A2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(new_n1008), .B(KEYINPUT110), .Z(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1018), .A2(new_n1030), .A3(new_n1006), .A4(new_n1013), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1014), .A2(new_n1040), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT112), .B(KEYINPUT63), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1039), .A2(G168), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1003), .B1(new_n1039), .B2(G168), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1054), .A2(new_n1052), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT62), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n1038), .A2(new_n1058), .A3(G2078), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1021), .A2(new_n780), .A3(new_n1022), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1025), .A2(new_n966), .A3(new_n1026), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT123), .B(G1961), .Z(new_n1062));
  AOI22_X1  g637(.A1(new_n1060), .A2(new_n1058), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(G301), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1057), .A2(new_n1033), .A3(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1055), .A2(new_n1056), .A3(KEYINPUT62), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1041), .B(new_n1051), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1027), .B2(G1956), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1061), .A2(KEYINPUT113), .A3(new_n796), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1021), .A2(new_n1071), .A3(new_n1022), .A4(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1022), .A2(new_n963), .A3(new_n966), .A4(new_n1072), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1069), .A2(new_n1070), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n560), .A2(new_n562), .ZN(new_n1077));
  OR2_X1    g652(.A1(new_n557), .A2(new_n1077), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n566), .B2(KEYINPUT57), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n560), .A2(new_n558), .A3(new_n562), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(new_n563), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n1085));
  NOR4_X1   g660(.A1(new_n1084), .A2(KEYINPUT115), .A3(new_n1085), .A4(new_n557), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1080), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1076), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1061), .A2(new_n850), .B1(new_n1002), .B2(new_n845), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n610), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n1076), .B2(new_n1087), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1076), .A2(new_n1092), .A3(new_n1087), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1091), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n600), .B1(new_n1090), .B2(KEYINPUT60), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT122), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1090), .A2(KEYINPUT60), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1098), .B(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1022), .A2(new_n963), .A3(new_n969), .A4(new_n966), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(new_n761), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n996), .A2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1101), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1102), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT120), .B(new_n759), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n759), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1111), .A3(KEYINPUT59), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT113), .B1(new_n1061), .B2(new_n796), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1070), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1087), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1087), .B(new_n1117), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(KEYINPUT117), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1088), .B1(new_n1125), .B2(new_n1094), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1115), .B(new_n1124), .C1(new_n1126), .C2(KEYINPUT61), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1100), .B1(new_n1127), .B2(KEYINPUT121), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1089), .B1(new_n1095), .B2(new_n1093), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1116), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1113), .A2(new_n1114), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1096), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n466), .A2(KEYINPUT124), .A3(new_n468), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT124), .B1(new_n466), .B2(new_n468), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n780), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1137), .A2(new_n474), .A3(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1022), .A2(new_n963), .A3(new_n1136), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1063), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(G171), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1135), .B1(new_n1064), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1033), .B(new_n1143), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1135), .B1(new_n1145), .B2(G301), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1141), .A2(G171), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(KEYINPUT125), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1147), .A2(KEYINPUT125), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1146), .B(KEYINPUT126), .C1(new_n1149), .C2(new_n1148), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1144), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1067), .B1(new_n1134), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n985), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G290), .B(new_n669), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n967), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n992), .B1(new_n1155), .B2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g734(.A1(new_n956), .A2(new_n957), .ZN(new_n1161));
  NOR2_X1   g735(.A1(new_n462), .A2(G227), .ZN(new_n1162));
  AND2_X1   g736(.A1(new_n903), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g737(.A1(new_n1163), .A2(new_n653), .A3(new_n702), .A4(new_n698), .ZN(new_n1164));
  NOR2_X1   g738(.A1(new_n1161), .A2(new_n1164), .ZN(G308));
  NAND2_X1  g739(.A1(new_n959), .A2(new_n955), .ZN(new_n1166));
  NAND4_X1  g740(.A1(new_n1166), .A2(new_n703), .A3(new_n653), .A4(new_n1163), .ZN(G225));
endmodule


