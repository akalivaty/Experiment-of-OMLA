//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(G952), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G902), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AOI211_X1 g008(.A(new_n193), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT21), .B(G898), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G214), .B1(G237), .B2(G902), .ZN(new_n199));
  OAI21_X1  g013(.A(G210), .B1(G237), .B2(G902), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G104), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G107), .ZN(new_n204));
  OAI21_X1  g018(.A(G101), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n206));
  AOI21_X1  g020(.A(G101), .B1(new_n203), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n201), .A3(G104), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G116), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G113), .ZN(new_n217));
  INV_X1    g031(.A(G113), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT2), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n213), .B(new_n215), .C1(new_n217), .C2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT5), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(G113), .C1(KEYINPUT5), .C2(new_n213), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n211), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n213), .A2(new_n215), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT2), .B(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n220), .A2(new_n226), .A3(KEYINPUT64), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n203), .A2(G107), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n206), .A2(new_n209), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(G101), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n223), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G122), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(KEYINPUT77), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n240), .B(new_n223), .C1(new_n234), .C2(new_n236), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT6), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n245), .A2(new_n229), .A3(new_n227), .A4(new_n233), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n240), .B1(new_n246), .B2(new_n223), .ZN(new_n247));
  OAI211_X1 g061(.A(KEYINPUT78), .B(new_n242), .C1(new_n244), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n237), .A2(new_n241), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT6), .A4(new_n243), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT1), .B1(new_n253), .B2(G146), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(G146), .ZN(new_n255));
  INV_X1    g069(.A(G146), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G143), .ZN(new_n257));
  OAI211_X1 g071(.A(G128), .B(new_n254), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G125), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(G146), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n260), .B(new_n261), .C1(KEYINPUT1), .C2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT0), .A4(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n255), .A2(new_n257), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G128), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n264), .B1(new_n268), .B2(new_n259), .ZN(new_n269));
  INV_X1    g083(.A(G224), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n271), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n252), .A2(new_n275), .ZN(new_n276));
  OR2_X1    g090(.A1(new_n271), .A2(KEYINPUT7), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n240), .B(KEYINPUT8), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n222), .A2(new_n220), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n205), .A2(new_n210), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n223), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  OR3_X1    g098(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n271), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n278), .A2(new_n243), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n193), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n200), .B1(new_n276), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n274), .B1(new_n248), .B2(new_n251), .ZN(new_n290));
  INV_X1    g104(.A(new_n200), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n290), .A2(new_n291), .A3(new_n287), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n198), .B(new_n199), .C1(new_n289), .C2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(G113), .B(G122), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(new_n203), .ZN(new_n295));
  XNOR2_X1  g109(.A(G125), .B(G140), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(new_n256), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n190), .A2(new_n194), .A3(G214), .ZN(new_n298));
  NAND2_X1  g112(.A1(KEYINPUT79), .A2(G143), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(KEYINPUT79), .A2(G143), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OR2_X1    g116(.A1(KEYINPUT79), .A2(G143), .ZN(new_n303));
  NOR2_X1   g117(.A1(G237), .A2(G953), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(G214), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT18), .ZN(new_n307));
  INV_X1    g121(.A(G131), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n303), .A2(new_n299), .B1(new_n304), .B2(G214), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n298), .A2(new_n301), .ZN(new_n311));
  OAI21_X1  g125(.A(G131), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI221_X1 g126(.A(new_n297), .B1(new_n306), .B2(new_n309), .C1(new_n312), .C2(new_n307), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n302), .A2(new_n308), .A3(new_n305), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT17), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n296), .A2(KEYINPUT16), .ZN(new_n319));
  OR3_X1    g133(.A1(new_n259), .A2(KEYINPUT16), .A3(G140), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n319), .A2(G146), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(G146), .B1(new_n319), .B2(new_n320), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT81), .A4(new_n315), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n312), .A2(KEYINPUT80), .A3(new_n315), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n308), .B1(new_n302), .B2(new_n305), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(KEYINPUT17), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n325), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n295), .B(new_n313), .C1(new_n324), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n312), .A2(new_n314), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n296), .B(KEYINPUT19), .Z(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(G146), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n319), .A2(G146), .A3(new_n320), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n320), .A4(G146), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n313), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n295), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n331), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n344));
  NOR2_X1   g158(.A1(G475), .A2(G902), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n331), .A2(new_n342), .A3(KEYINPUT82), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT82), .B1(new_n331), .B2(new_n342), .ZN(new_n348));
  INV_X1    g162(.A(new_n345), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n346), .B1(new_n350), .B2(new_n344), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n313), .B1(new_n324), .B2(new_n330), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n341), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n331), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n193), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G475), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G122), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT83), .B1(new_n358), .B2(G116), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n214), .A3(G122), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT84), .B1(new_n362), .B2(KEYINPUT14), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(G116), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT84), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT14), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n359), .A2(new_n361), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(KEYINPUT14), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n364), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G107), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n362), .A2(new_n201), .A3(new_n364), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n253), .A2(G128), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n262), .A2(G143), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G134), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n373), .A3(G134), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n362), .A2(new_n201), .A3(new_n364), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n201), .B1(new_n362), .B2(new_n364), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n373), .A2(new_n384), .A3(G134), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n376), .A2(new_n377), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n372), .A2(new_n373), .A3(new_n384), .A4(G134), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT9), .B(G234), .ZN(new_n390));
  INV_X1    g204(.A(G217), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n390), .A2(new_n391), .A3(G953), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n380), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n392), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n378), .B1(new_n369), .B2(G107), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n383), .A2(new_n388), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(new_n193), .ZN(new_n400));
  INV_X1    g214(.A(G478), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n401), .A2(KEYINPUT15), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n400), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n293), .A2(new_n357), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G221), .ZN(new_n406));
  INV_X1    g220(.A(new_n390), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n406), .B1(new_n407), .B2(new_n193), .ZN(new_n408));
  INV_X1    g222(.A(new_n268), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n245), .A2(new_n409), .A3(new_n233), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n258), .A2(new_n205), .A3(new_n210), .A4(new_n263), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT11), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n375), .B2(G137), .ZN(new_n416));
  INV_X1    g230(.A(G137), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT11), .A3(G134), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n375), .A2(G137), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G131), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n416), .A2(new_n418), .A3(new_n308), .A4(new_n419), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT65), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(KEYINPUT65), .A3(new_n422), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n414), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT10), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n211), .A2(new_n431), .A3(new_n263), .A4(new_n258), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n231), .A2(new_n232), .A3(G101), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(new_n268), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n430), .A2(new_n432), .B1(new_n434), .B2(new_n245), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT75), .B1(new_n435), .B2(new_n427), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT75), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n414), .A2(new_n437), .A3(new_n428), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n429), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n194), .A2(G227), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT76), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n435), .A2(new_n427), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n435), .A2(KEYINPUT75), .A3(new_n427), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n437), .B1(new_n414), .B2(new_n428), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT76), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n442), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n429), .A2(new_n442), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n258), .A2(new_n263), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n281), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n411), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT12), .B1(new_n428), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n454), .A2(KEYINPUT12), .A3(new_n423), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n451), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n444), .A2(new_n450), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G469), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n193), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n436), .A2(new_n438), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n445), .B1(new_n455), .B2(new_n456), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n461), .A2(new_n451), .B1(new_n462), .B2(new_n442), .ZN(new_n463));
  OAI21_X1  g277(.A(G469), .B1(new_n463), .B2(G902), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n408), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n405), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n425), .A2(new_n409), .A3(new_n426), .ZN(new_n467));
  INV_X1    g281(.A(new_n419), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n375), .A2(G137), .ZN(new_n469));
  OAI21_X1  g283(.A(G131), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n422), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(new_n452), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n227), .A2(new_n229), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n467), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n474), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n268), .B1(new_n422), .B2(new_n421), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n472), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT28), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT28), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT67), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n475), .A2(KEYINPUT67), .A3(new_n481), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n480), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n304), .A2(G210), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT27), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(G101), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n467), .A2(KEYINPUT30), .A3(new_n473), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n477), .B2(new_n472), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n476), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n490), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n475), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT29), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n485), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT67), .B1(new_n475), .B2(new_n481), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n467), .A2(new_n473), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n476), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n475), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT28), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n490), .A2(KEYINPUT29), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n193), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(G472), .B1(new_n498), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(G472), .A2(G902), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT68), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n481), .B1(new_n475), .B2(new_n478), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n499), .A2(new_n513), .A3(new_n500), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n512), .B1(new_n514), .B2(new_n490), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n486), .A2(KEYINPUT68), .A3(new_n496), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT31), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n475), .A2(new_n490), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n518), .B1(new_n519), .B2(new_n495), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n495), .A3(new_n518), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI211_X1 g337(.A(KEYINPUT66), .B(new_n518), .C1(new_n519), .C2(new_n495), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI211_X1 g339(.A(KEYINPUT32), .B(new_n511), .C1(new_n517), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT32), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n521), .ZN(new_n528));
  INV_X1    g342(.A(new_n520), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n524), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n486), .A2(KEYINPUT68), .A3(new_n496), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT68), .B1(new_n486), .B2(new_n496), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n527), .B1(new_n534), .B2(new_n510), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n509), .B1(new_n526), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(KEYINPUT69), .B(new_n509), .C1(new_n526), .C2(new_n535), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT24), .B(G110), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n212), .A2(G128), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT70), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n212), .A2(KEYINPUT70), .A3(G128), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n543), .B(new_n544), .C1(new_n212), .C2(G128), .ZN(new_n545));
  OAI22_X1  g359(.A1(new_n321), .A2(new_n322), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(new_n212), .B2(G128), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n541), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n551), .A2(G110), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT72), .B1(new_n546), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n322), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n335), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT72), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(G110), .A3(new_n552), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n545), .A2(new_n540), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n556), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n545), .A2(new_n540), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n550), .A2(G110), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n562), .A2(new_n563), .B1(new_n256), .B2(new_n296), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n337), .A3(new_n338), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT22), .B(G137), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n406), .A2(new_n189), .A3(G953), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n567), .B(new_n568), .Z(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n561), .A2(new_n565), .A3(new_n569), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n193), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT25), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n391), .B1(G234), .B2(new_n193), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n572), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n576), .A2(G902), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n575), .A2(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n538), .A2(new_n539), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT74), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT74), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n538), .A2(new_n583), .A3(new_n539), .A4(new_n580), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n466), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT86), .B(G101), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G3));
  INV_X1    g401(.A(new_n199), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n276), .A2(new_n200), .A3(new_n288), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n291), .B1(new_n290), .B2(new_n287), .ZN(new_n590));
  AOI211_X1 g404(.A(new_n197), .B(new_n588), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n398), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n401), .A2(G902), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n392), .B(KEYINPUT87), .Z(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n395), .B2(new_n396), .ZN(new_n596));
  OAI211_X1 g410(.A(KEYINPUT33), .B(new_n596), .C1(new_n393), .C2(KEYINPUT88), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n393), .A2(KEYINPUT88), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n593), .B(new_n594), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n398), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n401), .B1(new_n600), .B2(G902), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT89), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT89), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n599), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n591), .A2(new_n357), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT90), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n511), .B1(new_n517), .B2(new_n525), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n534), .A2(new_n193), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(G472), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n580), .A3(new_n465), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT91), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT34), .B(G104), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  NAND2_X1  g431(.A1(new_n350), .A2(new_n344), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT82), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n343), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n331), .A2(new_n342), .A3(KEYINPUT82), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n345), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT20), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n356), .A3(new_n404), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n293), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n613), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT92), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT35), .B(G107), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  AND2_X1   g444(.A1(new_n573), .A2(new_n574), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n573), .A2(new_n574), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n576), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n570), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT93), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n566), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n579), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n611), .A2(new_n405), .A3(new_n465), .A4(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  INV_X1    g455(.A(new_n465), .ZN(new_n642));
  INV_X1    g456(.A(new_n638), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n192), .B1(new_n195), .B2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n625), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n538), .A2(new_n539), .A3(new_n644), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  NOR2_X1   g465(.A1(new_n532), .A2(new_n533), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n530), .A2(new_n531), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n510), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT32), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n609), .A2(new_n527), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n495), .A2(new_n475), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n490), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n193), .B1(new_n504), .B2(new_n490), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT94), .Z(new_n664));
  XOR2_X1   g478(.A(new_n648), .B(KEYINPUT39), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n465), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n643), .A2(new_n199), .A3(new_n357), .A4(new_n404), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n289), .A2(new_n292), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT38), .ZN(new_n671));
  OR3_X1    g485(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n664), .A2(new_n667), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n253), .ZN(G45));
  INV_X1    g488(.A(new_n648), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n357), .A2(new_n606), .A3(new_n645), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT95), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n677), .A2(new_n538), .A3(new_n539), .A4(new_n644), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  AOI21_X1  g493(.A(KEYINPUT69), .B1(new_n657), .B2(new_n509), .ZN(new_n680));
  INV_X1    g494(.A(new_n539), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n458), .A2(new_n193), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G469), .ZN(new_n684));
  INV_X1    g498(.A(new_n408), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n460), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT96), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT96), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n684), .A2(new_n688), .A3(new_n685), .A4(new_n460), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n682), .A2(new_n580), .A3(new_n608), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n682), .A2(new_n580), .A3(new_n626), .A4(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  AOI22_X1  g509(.A1(new_n623), .A2(new_n346), .B1(G475), .B2(new_n355), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n198), .A3(new_n403), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n458), .A2(new_n459), .A3(new_n193), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n459), .B1(new_n458), .B2(new_n193), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT97), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n701), .A3(new_n685), .A4(new_n645), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n684), .A2(new_n685), .A3(new_n460), .A4(new_n645), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT97), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n697), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n682), .A2(new_n638), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  NOR3_X1   g521(.A1(new_n293), .A2(new_n696), .A3(new_n403), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n687), .A2(new_n689), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n610), .A2(G472), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n510), .B(KEYINPUT98), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n529), .A2(new_n522), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n490), .B1(new_n501), .B2(new_n505), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n710), .A2(new_n580), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT99), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n710), .A2(KEYINPUT99), .A3(new_n580), .A4(new_n714), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n709), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n358), .ZN(G24));
  NAND2_X1  g534(.A1(new_n702), .A2(new_n704), .ZN(new_n721));
  AOI21_X1  g535(.A(G902), .B1(new_n517), .B2(new_n525), .ZN(new_n722));
  INV_X1    g536(.A(G472), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n638), .B(new_n714), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n357), .A2(new_n606), .A3(new_n675), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n721), .A2(new_n726), .A3(KEYINPUT100), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT100), .B1(new_n721), .B2(new_n726), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n259), .ZN(G27));
  AND2_X1   g544(.A1(new_n536), .A2(new_n580), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n289), .A2(new_n292), .A3(new_n588), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n465), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n725), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n731), .A2(KEYINPUT42), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n538), .A2(new_n539), .A3(new_n734), .A4(new_n580), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT101), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n735), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NOR3_X1   g556(.A1(new_n733), .A2(new_n625), .A3(new_n648), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n538), .A2(new_n743), .A3(new_n539), .A4(new_n580), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  AND2_X1   g559(.A1(new_n603), .A2(new_n605), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n357), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT102), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n747), .B(KEYINPUT43), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT102), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n611), .A2(new_n643), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n755), .A2(KEYINPUT104), .A3(new_n756), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n755), .A2(new_n756), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n463), .A2(KEYINPUT45), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n463), .A2(KEYINPUT45), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(G469), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(G469), .A2(G902), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n460), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n766), .A2(new_n767), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n685), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n665), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n732), .B(KEYINPUT103), .Z(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  INV_X1    g591(.A(new_n732), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n725), .A2(new_n580), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n771), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(KEYINPUT47), .B(new_n685), .C1(new_n769), .C2(new_n770), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n680), .B2(new_n681), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NOR2_X1   g599(.A1(new_n408), .A2(new_n588), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n580), .A2(new_n671), .A3(new_n747), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n700), .B(KEYINPUT49), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n664), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n591), .A2(KEYINPUT105), .A3(new_n696), .A4(new_n404), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT105), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n351), .A2(new_n404), .A3(new_n356), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n793), .B2(new_n293), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n791), .A2(new_n794), .A3(new_n607), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n639), .B1(new_n795), .B2(new_n612), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n719), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(new_n706), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n582), .A2(new_n584), .ZN(new_n799));
  INV_X1    g613(.A(new_n466), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n798), .A2(new_n801), .A3(new_n691), .A4(new_n694), .ZN(new_n802));
  INV_X1    g616(.A(new_n724), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n734), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n744), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n624), .A2(new_n356), .A3(new_n403), .A4(new_n675), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n733), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n538), .A2(new_n539), .A3(new_n638), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT106), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n805), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n741), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n802), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n650), .B1(new_n727), .B2(new_n728), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT107), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT107), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n817), .B(new_n650), .C1(new_n727), .C2(new_n728), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n646), .A2(new_n696), .A3(new_n403), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n642), .A2(new_n638), .A3(new_n648), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n663), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n678), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(new_n818), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n823), .B1(new_n815), .B2(new_n822), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(KEYINPUT108), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT108), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n814), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OR3_X1    g645(.A1(new_n815), .A2(new_n823), .A3(new_n822), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n826), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n814), .A2(KEYINPUT53), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT109), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n790), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n814), .B(KEYINPUT53), .C1(new_n827), .C2(new_n828), .ZN(new_n840));
  INV_X1    g654(.A(new_n833), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n691), .A2(new_n694), .A3(new_n706), .A4(new_n797), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n585), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n741), .A3(new_n812), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n830), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n840), .A2(new_n845), .A3(new_n790), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n191), .B(new_n749), .C1(new_n717), .C2(new_n718), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n700), .A2(new_n408), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n781), .A2(new_n782), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n774), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n686), .A2(new_n778), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n852), .A2(new_n580), .A3(new_n192), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n664), .A2(new_n696), .A3(new_n746), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n749), .A2(new_n191), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n803), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n671), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n858), .A2(new_n199), .A3(new_n686), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n848), .A2(new_n859), .ZN(new_n860));
  OR3_X1    g674(.A1(new_n860), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(KEYINPUT110), .B2(KEYINPUT50), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n857), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n851), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(KEYINPUT111), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n851), .A2(new_n866), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n863), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n848), .A2(new_n721), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT112), .Z(new_n872));
  NAND3_X1  g686(.A1(new_n855), .A2(new_n731), .A3(new_n852), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT48), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n746), .A2(new_n696), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n664), .A2(new_n875), .A3(new_n853), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n188), .A2(new_n872), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n867), .A2(new_n870), .A3(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n839), .A2(new_n847), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(G952), .A2(G953), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT113), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n789), .B1(new_n879), .B2(new_n881), .ZN(G75));
  NAND2_X1  g696(.A1(new_n187), .A2(G953), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT116), .Z(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT117), .Z(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n840), .A2(new_n845), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(G902), .ZN(new_n888));
  INV_X1    g702(.A(G210), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n252), .B(new_n275), .ZN(new_n891));
  XNOR2_X1  g705(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n885), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n893), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT115), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n897), .A3(new_n893), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n896), .B2(new_n898), .ZN(G51));
  INV_X1    g713(.A(new_n884), .ZN(new_n900));
  INV_X1    g714(.A(new_n764), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n843), .A2(KEYINPUT53), .A3(new_n741), .A4(new_n812), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n825), .A2(new_n826), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT108), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n825), .A2(KEYINPUT108), .A3(new_n826), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT53), .B1(new_n814), .B2(new_n833), .ZN(new_n908));
  OAI211_X1 g722(.A(G902), .B(new_n901), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT120), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n887), .A2(new_n911), .A3(G902), .A4(new_n901), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n458), .B(KEYINPUT118), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n907), .B2(new_n908), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n846), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n765), .B(KEYINPUT57), .Z(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n913), .B1(new_n918), .B2(KEYINPUT119), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  INV_X1    g734(.A(new_n917), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n915), .B2(new_n846), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n922), .B2(new_n914), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n900), .B1(new_n919), .B2(new_n923), .ZN(G54));
  NAND2_X1  g738(.A1(new_n620), .A2(new_n621), .ZN(new_n925));
  NAND2_X1  g739(.A1(KEYINPUT58), .A2(G475), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n888), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n884), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n888), .A2(new_n925), .A3(new_n926), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G60));
  OAI21_X1  g744(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT121), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT59), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n916), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n885), .ZN(new_n937));
  INV_X1    g751(.A(new_n934), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n839), .B2(new_n847), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n939), .B2(new_n932), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT123), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n887), .A2(new_n636), .A3(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n887), .A2(new_n944), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n885), .B(new_n945), .C1(new_n946), .C2(new_n578), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G66));
  OAI21_X1  g763(.A(G953), .B1(new_n196), .B2(new_n270), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n843), .B2(G953), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n248), .B(new_n251), .C1(G898), .C2(new_n194), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G69));
  NAND3_X1  g767(.A1(new_n773), .A2(new_n731), .A3(new_n819), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n784), .A2(new_n744), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n776), .A2(new_n955), .A3(new_n741), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n816), .A2(new_n678), .A3(new_n818), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n194), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n647), .A2(G953), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n958), .B2(new_n960), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(G227), .A2(G900), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n492), .A2(new_n494), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n333), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n963), .A2(G953), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n961), .B2(new_n962), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n964), .A2(G953), .ZN(new_n969));
  INV_X1    g783(.A(new_n875), .ZN(new_n970));
  AOI211_X1 g784(.A(new_n778), .B(new_n666), .C1(new_n970), .C2(new_n793), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n799), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT124), .Z(new_n973));
  AND3_X1   g787(.A1(new_n973), .A2(new_n776), .A3(new_n784), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n957), .A2(new_n673), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(KEYINPUT62), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n966), .A2(G953), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n968), .B(new_n969), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n967), .A2(new_n981), .ZN(G72));
  NAND3_X1  g796(.A1(new_n838), .A2(new_n831), .A3(new_n836), .ZN(new_n983));
  XNOR2_X1  g797(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n723), .A2(new_n193), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n983), .A2(new_n497), .A3(new_n659), .A4(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n978), .B2(new_n802), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n660), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n956), .A2(new_n957), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n986), .B1(new_n990), .B2(new_n802), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n497), .B(KEYINPUT127), .Z(new_n992));
  AOI21_X1  g806(.A(new_n900), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n987), .A2(new_n989), .A3(new_n993), .ZN(G57));
endmodule


