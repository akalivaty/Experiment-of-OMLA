//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n458), .B1(new_n449), .B2(new_n455), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT67), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n468), .A2(new_n465), .A3(G101), .A4(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n464), .A2(G137), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n463), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n463), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n465), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n463), .B2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n480), .B1(new_n485), .B2(G136), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT69), .Z(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n461), .B2(new_n462), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n462), .C2(new_n461), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  XOR2_X1   g075(.A(KEYINPUT5), .B(G543), .Z(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G88), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n506), .A2(KEYINPUT70), .A3(new_n509), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT71), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR3_X1    g092(.A1(new_n515), .A2(KEYINPUT71), .A3(new_n516), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n512), .A2(new_n513), .B1(new_n517), .B2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n520));
  XOR2_X1   g095(.A(new_n520), .B(KEYINPUT72), .Z(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT74), .B(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n505), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n526), .A2(new_n527), .B1(new_n508), .B2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n521), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G168));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  INV_X1    g106(.A(G77), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n501), .A2(new_n531), .B1(new_n532), .B2(new_n507), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT75), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n535), .B1(new_n532), .B2(new_n507), .C1(new_n501), .C2(new_n531), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n534), .A2(G651), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n505), .A2(G90), .B1(new_n508), .B2(G52), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n502), .A2(new_n503), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n514), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n544), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n516), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n546), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n508), .A2(new_n560), .A3(G53), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OR3_X1    g137(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT77), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n547), .A2(KEYINPUT77), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(new_n564), .A3(G91), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n516), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT78), .A4(new_n567), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n529), .A2(KEYINPUT79), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n521), .A2(new_n528), .A3(new_n575), .A4(new_n523), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n574), .A2(new_n576), .ZN(G286));
  NAND2_X1  g152(.A1(new_n512), .A2(new_n513), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n518), .A2(new_n517), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G303));
  NAND3_X1  g155(.A1(new_n563), .A2(new_n564), .A3(G87), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n514), .A2(G74), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(new_n508), .B2(G49), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G288));
  NAND3_X1  g159(.A1(new_n563), .A2(new_n564), .A3(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n501), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n508), .B2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n514), .A2(G60), .ZN(new_n591));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n516), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n505), .A2(G85), .B1(new_n508), .B2(G47), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n563), .A2(new_n564), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n603));
  INV_X1    g178(.A(G54), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n546), .B2(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n501), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n603), .A2(new_n605), .B1(G651), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n599), .B1(new_n610), .B2(G868), .ZN(G321));
  XOR2_X1   g186(.A(G321), .B(KEYINPUT82), .Z(G284));
  MUX2_X1   g187(.A(G299), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g188(.A(G280), .B(KEYINPUT83), .Z(G297));
  NAND2_X1  g189(.A1(new_n602), .A2(new_n609), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(G559), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G860), .B2(new_n610), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT84), .Z(G148));
  INV_X1    g193(.A(new_n552), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n616), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g198(.A(G2104), .ZN(new_n624));
  NOR3_X1   g199(.A1(new_n463), .A2(new_n624), .A3(G2105), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT86), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n476), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n465), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n632), .B1(new_n633), .B2(new_n634), .C1(new_n484), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n629), .A2(G2100), .ZN(new_n639));
  NAND4_X1  g214(.A1(new_n631), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT87), .Z(G401));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  INV_X1    g237(.A(new_n659), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n663), .B2(new_n657), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n657), .B(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n664), .B1(new_n666), .B2(new_n663), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n663), .A3(new_n660), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n673), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n673), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G24), .ZN(new_n690));
  INV_X1    g265(.A(G290), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  INV_X1    g267(.A(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G25), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g273(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n699));
  OAI221_X1 g274(.A(G2104), .B1(G107), .B2(new_n465), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT90), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n485), .A2(G131), .ZN(new_n702));
  AOI211_X1 g277(.A(new_n701), .B(new_n702), .C1(G119), .C2(new_n476), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n696), .B1(new_n703), .B2(new_n695), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT91), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n704), .B(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G6), .B(G305), .S(G16), .Z(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT32), .B(G1981), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G1971), .ZN(new_n712));
  NAND2_X1  g287(.A1(G166), .A2(G16), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G16), .B2(G22), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G23), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT92), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G288), .B2(new_n689), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT33), .B(G1976), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT93), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n715), .B(new_n721), .C1(new_n712), .C2(new_n714), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n694), .B(new_n708), .C1(new_n722), .C2(KEYINPUT34), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(KEYINPUT34), .B2(new_n722), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT36), .Z(new_n725));
  NAND2_X1  g300(.A1(G160), .A2(G29), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT99), .B(KEYINPUT24), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(new_n695), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G2084), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT100), .Z(new_n732));
  NOR2_X1   g307(.A1(G168), .A2(new_n689), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n689), .B2(G21), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT31), .B(G11), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n738), .A2(G28), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n695), .B1(new_n738), .B2(G28), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n737), .B1(new_n739), .B2(new_n740), .C1(new_n636), .C2(new_n695), .ZN(new_n741));
  INV_X1    g316(.A(new_n730), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n695), .A2(G27), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G164), .B2(new_n695), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2078), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n734), .B2(new_n735), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n732), .A2(new_n736), .A3(new_n744), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n689), .A2(G19), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n552), .B2(new_n689), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT94), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1341), .ZN(new_n753));
  NOR2_X1   g328(.A1(G4), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n610), .B2(G16), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(G1348), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n749), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n695), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n476), .A2(G128), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n465), .A2(G116), .ZN(new_n761));
  OAI21_X1  g336(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n762));
  INV_X1    g337(.A(G140), .ZN(new_n763));
  OAI221_X1 g338(.A(new_n760), .B1(new_n761), .B2(new_n762), .C1(new_n484), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT96), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT95), .B(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n695), .A2(G32), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n485), .A2(G141), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT26), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n771), .B(new_n773), .C1(G129), .C2(new_n476), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT101), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n769), .B1(new_n776), .B2(new_n695), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT27), .B(G1996), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n757), .A2(new_n768), .A3(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n695), .A2(G33), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT25), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n485), .A2(G139), .ZN(new_n784));
  NAND2_X1  g359(.A1(G115), .A2(G2104), .ZN(new_n785));
  INV_X1    g360(.A(G127), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n463), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT97), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n465), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n788), .B2(new_n787), .ZN(new_n790));
  AOI211_X1 g365(.A(new_n783), .B(new_n784), .C1(KEYINPUT98), .C2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(KEYINPUT98), .B2(new_n790), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n781), .B1(new_n792), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2072), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  NOR2_X1   g371(.A1(G171), .A2(new_n689), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G5), .B2(new_n689), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n796), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n793), .B2(new_n794), .ZN(new_n801));
  NOR2_X1   g376(.A1(G29), .A2(G35), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G162), .B2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT29), .B(G2090), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n689), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT23), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n572), .B2(new_n689), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT102), .B(G1956), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n755), .A2(G1348), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n803), .A2(new_n804), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n805), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n780), .A2(new_n799), .A3(new_n801), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n725), .A2(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  XOR2_X1   g391(.A(KEYINPUT104), .B(G93), .Z(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT103), .B(G55), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n547), .A2(new_n817), .B1(new_n546), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n516), .ZN(new_n821));
  OAI21_X1  g396(.A(G860), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n610), .A2(G559), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT105), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n819), .A2(new_n821), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n552), .B(new_n828), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n831));
  AOI21_X1  g406(.A(G860), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT106), .ZN(new_n833));
  INV_X1    g408(.A(new_n829), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n827), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n833), .B1(new_n832), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n823), .B1(new_n837), .B2(new_n838), .ZN(G145));
  XOR2_X1   g414(.A(KEYINPUT108), .B(G37), .Z(new_n840));
  NOR2_X1   g415(.A1(new_n792), .A2(new_n776), .ZN(new_n841));
  INV_X1    g416(.A(new_n775), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n841), .B1(new_n792), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  INV_X1    g419(.A(G118), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n844), .B1(new_n845), .B2(G2105), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n485), .A2(G142), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT107), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  AOI211_X1 g424(.A(new_n846), .B(new_n849), .C1(G130), .C2(new_n476), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n764), .B(G164), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n703), .B(new_n627), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n851), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n853), .B1(new_n852), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n843), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(G162), .B(new_n636), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(G160), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n850), .B(new_n851), .ZN(new_n861));
  INV_X1    g436(.A(new_n853), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n843), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n855), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n858), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n860), .B1(new_n858), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n840), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g444(.A1(new_n615), .A2(new_n572), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT109), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n602), .A2(new_n570), .A3(new_n571), .A4(new_n609), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(G299), .A2(new_n610), .A3(KEYINPUT109), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(KEYINPUT41), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n870), .A2(new_n876), .A3(new_n872), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n616), .B(new_n834), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n616), .B(new_n829), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(new_n874), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT42), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n886), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(G166), .B(new_n691), .ZN(new_n889));
  XOR2_X1   g464(.A(G305), .B(G288), .Z(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(KEYINPUT110), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n885), .A2(new_n893), .A3(new_n887), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n620), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n828), .A2(G868), .ZN(new_n898));
  OR3_X1    g473(.A1(new_n897), .A2(KEYINPUT111), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT111), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(G295));
  OR2_X1    g476(.A1(new_n897), .A2(new_n898), .ZN(G331));
  NAND2_X1  g477(.A1(G301), .A2(G168), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT112), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n540), .A2(new_n541), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n906), .A2(new_n574), .A3(new_n539), .A4(new_n576), .ZN(new_n907));
  NAND3_X1  g482(.A1(G301), .A2(KEYINPUT112), .A3(G168), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n905), .A2(new_n834), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n907), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT112), .B1(G301), .B2(G168), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n829), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n909), .A2(new_n912), .B1(new_n875), .B2(new_n877), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n912), .A2(new_n882), .A3(new_n909), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n892), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n913), .A2(new_n914), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n917), .B2(new_n891), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n918), .B2(KEYINPUT113), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT113), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n913), .A2(new_n914), .A3(new_n892), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(G37), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT43), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n876), .B1(new_n912), .B2(new_n909), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n870), .A2(new_n872), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n882), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n926), .B(new_n891), .C1(new_n927), .C2(new_n924), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(new_n915), .A3(new_n840), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n923), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n919), .B2(new_n922), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n932), .B1(new_n935), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g511(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G164), .B2(G1384), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n470), .A2(new_n474), .A3(G40), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  INV_X1    g517(.A(new_n499), .ZN(new_n943));
  XNOR2_X1  g518(.A(KEYINPUT3), .B(G2104), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n498), .B1(new_n944), .B2(new_n495), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g521(.A(KEYINPUT45), .B(new_n942), .C1(new_n946), .C2(new_n493), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(G2078), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n470), .A2(new_n474), .A3(G40), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT115), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT50), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n956), .B(new_n942), .C1(new_n946), .C2(new_n493), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n942), .B1(new_n946), .B2(new_n493), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n953), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n952), .B1(new_n961), .B2(G1961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT123), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n939), .A2(new_n964), .A3(new_n947), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n959), .A2(KEYINPUT114), .A3(new_n938), .ZN(new_n966));
  AOI211_X1 g541(.A(G2078), .B(new_n953), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n967), .B2(KEYINPUT53), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n966), .ZN(new_n969));
  INV_X1    g544(.A(G2078), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n970), .A3(new_n940), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(KEYINPUT123), .A3(new_n950), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n962), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n973), .A2(KEYINPUT124), .A3(G301), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT124), .ZN(new_n975));
  INV_X1    g550(.A(new_n962), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n953), .B1(new_n965), .B2(new_n966), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n963), .B(KEYINPUT53), .C1(new_n977), .C2(new_n970), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT123), .B1(new_n971), .B2(new_n950), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(new_n980), .B2(G171), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n974), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n976), .B(G301), .C1(new_n978), .C2(new_n979), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT125), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n973), .A2(KEYINPUT125), .A3(G301), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n937), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT126), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT54), .B1(new_n973), .B2(G301), .ZN(new_n990));
  INV_X1    g565(.A(new_n983), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n980), .A2(G171), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(KEYINPUT126), .A3(KEYINPUT54), .A4(new_n983), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n954), .A2(new_n940), .A3(new_n957), .ZN(new_n996));
  INV_X1    g571(.A(G1956), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(KEYINPUT117), .A3(new_n997), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n568), .B(KEYINPUT57), .Z(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT56), .B(G2072), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n977), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n961), .A2(G1348), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n959), .A2(new_n953), .ZN(new_n1009));
  INV_X1    g584(.A(G2067), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n615), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1006), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT118), .B(new_n1006), .C1(new_n1007), .C2(new_n1012), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT61), .ZN(new_n1017));
  AND4_X1   g592(.A1(new_n1003), .A2(new_n1005), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1007), .B2(new_n1018), .ZN(new_n1019));
  OAI221_X1 g594(.A(new_n1011), .B1(new_n961), .B2(G1348), .C1(new_n610), .C2(KEYINPUT60), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n610), .A2(KEYINPUT60), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1008), .A2(KEYINPUT60), .A3(new_n610), .A4(new_n1011), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1003), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1005), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1006), .A2(new_n1028), .A3(KEYINPUT61), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1019), .A2(new_n1024), .A3(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n552), .A2(KEYINPUT120), .ZN(new_n1031));
  AOI211_X1 g606(.A(G1996), .B(new_n953), .C1(new_n965), .C2(new_n966), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT58), .B(G1341), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1032), .A2(KEYINPUT119), .B1(new_n1009), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1996), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n977), .A2(KEYINPUT119), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1031), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT59), .B(new_n1031), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1015), .B(new_n1016), .C1(new_n1030), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n588), .A2(G651), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n508), .A2(G48), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n505), .A2(G86), .ZN(new_n1046));
  OAI21_X1  g621(.A(G1981), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n585), .A2(new_n1048), .A3(new_n589), .ZN(new_n1049));
  OR2_X1    g624(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G8), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G164), .A2(G1384), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n940), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1050), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G288), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G1976), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1059), .A2(new_n1054), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n1059), .B2(new_n1054), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1057), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(G166), .B2(new_n1052), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n977), .A2(G1971), .ZN(new_n1070));
  AOI211_X1 g645(.A(G2090), .B(new_n953), .C1(new_n958), .C2(new_n960), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1069), .B(G8), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1065), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1069), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n996), .A2(G2090), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n969), .A2(new_n940), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(new_n712), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1077), .B2(new_n1052), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n940), .A2(new_n743), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n958), .B2(new_n960), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n953), .B1(new_n959), .B2(new_n938), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1966), .B1(new_n1083), .B2(new_n947), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1082), .A2(new_n1084), .A3(new_n529), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1080), .B1(new_n1085), .B2(new_n1052), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n958), .A2(new_n960), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1081), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n735), .B1(new_n941), .B2(new_n948), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(G168), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n529), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1086), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1094), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1079), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n988), .A2(new_n995), .A3(new_n1042), .A4(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1099), .A2(new_n1052), .A3(G286), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1078), .A2(new_n1072), .A3(new_n1065), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G286), .A2(new_n1052), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(KEYINPUT63), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(G8), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1074), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1073), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1072), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1049), .B1(new_n1057), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1111), .A2(new_n1065), .B1(new_n1054), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1086), .A2(new_n1093), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1086), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT62), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT124), .B1(new_n973), .B2(G301), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n980), .A2(new_n975), .A3(G171), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1079), .B1(new_n1124), .B2(KEYINPUT62), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1115), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1098), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n939), .A2(new_n953), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n776), .A2(new_n1035), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n764), .B(new_n1010), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1130), .B(new_n1131), .C1(new_n1035), .C2(new_n842), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n703), .B(new_n707), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(G290), .B(new_n693), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1129), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1127), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n691), .A2(new_n1128), .A3(new_n693), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT48), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1134), .B2(new_n1129), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n703), .A2(new_n707), .ZN(new_n1142));
  OAI22_X1  g717(.A1(new_n1132), .A2(new_n1142), .B1(G2067), .B2(new_n764), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1128), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1129), .B1(new_n1131), .B2(new_n842), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT46), .B1(new_n1129), .B2(G1996), .ZN(new_n1147));
  OR3_X1    g722(.A1(new_n1129), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT47), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1138), .A2(KEYINPUT127), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1136), .B1(new_n1098), .B2(new_n1126), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1151), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1152), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g732(.A(G319), .ZN(new_n1159));
  NOR4_X1   g733(.A1(G229), .A2(new_n1159), .A3(new_n655), .A4(G227), .ZN(new_n1160));
  OAI211_X1 g734(.A(new_n868), .B(new_n1160), .C1(new_n933), .C2(new_n934), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


