//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980;
  AND2_X1   g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT29), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT65), .A2(KEYINPUT27), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT65), .A2(KEYINPUT27), .ZN(new_n214));
  OAI21_X1  g013(.A(G183gat), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g016(.A(KEYINPUT66), .B(G183gat), .C1(new_n213), .C2(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  AOI21_X1  g018(.A(G190gat), .B1(new_n219), .B2(KEYINPUT27), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT28), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT28), .A3(new_n220), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n212), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NOR3_X1   g028(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n209), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  AND2_X1   g031(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n211), .A2(new_n232), .B1(new_n233), .B2(G190gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n227), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n211), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n209), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n205), .A3(new_n206), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n241), .B2(new_n228), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n242), .A3(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n203), .B1(new_n226), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n212), .ZN(new_n247));
  INV_X1    g046(.A(new_n220), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n248), .B1(new_n215), .B2(new_n216), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT28), .B1(new_n249), .B2(new_n218), .ZN(new_n250));
  INV_X1    g049(.A(new_n225), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n238), .A2(new_n242), .A3(KEYINPUT25), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT25), .B1(new_n238), .B2(new_n242), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT64), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n235), .A2(new_n256), .A3(new_n243), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n252), .A2(new_n202), .A3(new_n255), .A4(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT72), .ZN(new_n259));
  INV_X1    g058(.A(G211gat), .ZN(new_n260));
  INV_X1    g059(.A(G218gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G211gat), .A2(G218gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT22), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n262), .A2(new_n259), .A3(new_n263), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n265), .A2(new_n267), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n267), .ZN(new_n271));
  INV_X1    g070(.A(new_n269), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n272), .B2(new_n264), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n246), .A2(new_n258), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT73), .ZN(new_n278));
  XNOR2_X1  g077(.A(G64gat), .B(G92gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n226), .A2(new_n245), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n251), .B1(new_n221), .B2(new_n222), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n255), .B(new_n257), .C1(new_n283), .C2(new_n212), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n282), .A2(new_n202), .B1(new_n284), .B2(new_n203), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n276), .B(new_n281), .C1(new_n285), .C2(new_n275), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT74), .ZN(new_n287));
  INV_X1    g086(.A(new_n203), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n235), .A2(new_n256), .A3(new_n243), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n256), .B1(new_n235), .B2(new_n243), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n288), .B1(new_n291), .B2(new_n252), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n252), .A2(new_n202), .A3(new_n244), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n274), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n276), .A4(new_n281), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n281), .B1(new_n295), .B2(new_n276), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n287), .A2(new_n297), .B1(KEYINPUT30), .B2(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n246), .A2(new_n275), .A3(new_n258), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n255), .A2(new_n257), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n203), .B1(new_n301), .B2(new_n226), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n275), .B1(new_n302), .B2(new_n293), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n280), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT75), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT30), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n307), .B(new_n280), .C1(new_n300), .C2(new_n303), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n299), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G1gat), .B(G29gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT0), .ZN(new_n313));
  XNOR2_X1  g112(.A(G57gat), .B(G85gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G162gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT78), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G162gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n316), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT79), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT79), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT78), .B(G162gat), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n324), .B(KEYINPUT2), .C1(new_n325), .C2(new_n316), .ZN(new_n326));
  NOR2_X1   g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327));
  AND2_X1   g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n316), .A2(new_n317), .ZN(new_n330));
  AOI211_X1 g129(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n323), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n329), .ZN(new_n333));
  NOR2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT76), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OR3_X1    g134(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT76), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n328), .B2(new_n327), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(KEYINPUT2), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n328), .A2(new_n327), .A3(new_n337), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n335), .B(new_n336), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT3), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n332), .A2(new_n345), .A3(new_n342), .ZN(new_n346));
  INV_X1    g145(.A(G134gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G127gat), .ZN(new_n348));
  INV_X1    g147(.A(G127gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G134gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n351), .A2(KEYINPUT1), .ZN(new_n352));
  INV_X1    g151(.A(G113gat), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT67), .B1(new_n353), .B2(G120gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT67), .ZN(new_n355));
  INV_X1    g154(.A(G120gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(G113gat), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n354), .B(new_n357), .C1(G113gat), .C2(new_n356), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n353), .A2(G120gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n356), .A2(G113gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n352), .A2(new_n358), .B1(new_n362), .B2(new_n351), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n344), .A2(new_n346), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n332), .A2(new_n342), .A3(new_n363), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n332), .A2(new_n342), .A3(KEYINPUT4), .A4(new_n363), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n365), .A2(new_n366), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n343), .A2(new_n364), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n367), .ZN(new_n374));
  INV_X1    g173(.A(new_n366), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n344), .A2(new_n346), .A3(new_n364), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n369), .A2(new_n370), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n379), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n378), .B1(new_n381), .B2(new_n372), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n371), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n315), .B(new_n377), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT6), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n379), .A2(new_n380), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n387), .A2(new_n378), .A3(new_n372), .A4(new_n366), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT80), .B1(new_n371), .B2(KEYINPUT5), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n388), .A2(new_n389), .B1(new_n371), .B2(new_n376), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(new_n315), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n377), .B1(new_n382), .B2(new_n383), .ZN(new_n393));
  INV_X1    g192(.A(new_n315), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT6), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n311), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n275), .B1(new_n346), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n270), .A2(new_n273), .A3(new_n398), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n400), .A2(new_n345), .B1(new_n342), .B2(new_n332), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT82), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G228gat), .ZN(new_n403));
  INV_X1    g202(.A(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n346), .A2(new_n398), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n274), .ZN(new_n408));
  INV_X1    g207(.A(new_n401), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n402), .B(new_n405), .C1(new_n410), .C2(KEYINPUT82), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n400), .A2(new_n345), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n407), .A2(new_n274), .B1(new_n413), .B2(new_n343), .ZN(new_n414));
  OAI221_X1 g213(.A(new_n412), .B1(new_n403), .B2(new_n404), .C1(new_n414), .C2(new_n406), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G22gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(G22gat), .A3(new_n415), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT31), .B(G50gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  AOI21_X1  g222(.A(G22gat), .B1(new_n411), .B2(new_n415), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n418), .A2(new_n425), .A3(new_n419), .A4(new_n423), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT34), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n284), .A2(new_n363), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n252), .A2(new_n364), .A3(new_n255), .A4(new_n257), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G227gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(new_n404), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n429), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  AOI211_X1 g235(.A(KEYINPUT34), .B(new_n434), .C1(new_n430), .C2(new_n431), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT71), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n434), .A3(new_n431), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT32), .ZN(new_n440));
  XOR2_X1   g239(.A(G15gat), .B(G43gat), .Z(new_n441));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n440), .B1(new_n446), .B2(KEYINPUT33), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n440), .A2(KEYINPUT33), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n439), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n451), .B2(new_n446), .ZN(new_n452));
  AOI211_X1 g251(.A(KEYINPUT70), .B(new_n445), .C1(new_n439), .C2(new_n450), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n438), .B(new_n448), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n448), .B1(new_n452), .B2(new_n453), .ZN(new_n455));
  INV_X1    g254(.A(new_n438), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n427), .A2(new_n428), .A3(new_n454), .A4(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT35), .B1(new_n397), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n427), .A2(new_n428), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n310), .A2(KEYINPUT84), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n299), .A2(new_n309), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT6), .B1(new_n390), .B2(new_n315), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n393), .A2(new_n394), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n395), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n436), .A2(new_n437), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n469), .B(new_n448), .C1(new_n452), .C2(new_n453), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n460), .A2(new_n464), .A3(new_n468), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n369), .A2(new_n370), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n366), .B1(new_n477), .B2(new_n365), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT39), .B1(new_n374), .B2(new_n375), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(new_n375), .C1(new_n379), .C2(new_n380), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n480), .A2(KEYINPUT40), .A3(new_n315), .A4(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n482), .B(new_n315), .C1(new_n478), .C2(new_n479), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT40), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(new_n391), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n461), .A2(new_n463), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n300), .A2(new_n303), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n281), .B1(new_n490), .B2(KEYINPUT37), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT38), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n302), .A2(new_n293), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT37), .B1(new_n493), .B2(new_n274), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n275), .B1(new_n246), .B2(new_n258), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT85), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n281), .A2(KEYINPUT37), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n286), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n495), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n500), .B(KEYINPUT37), .C1(new_n493), .C2(new_n274), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT85), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n499), .A2(new_n501), .A3(new_n502), .A4(new_n492), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n490), .A2(KEYINPUT37), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n492), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n305), .A2(new_n308), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n467), .A2(new_n504), .A3(new_n508), .A4(new_n395), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n460), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n427), .A2(new_n428), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n397), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n471), .A2(new_n513), .A3(new_n473), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n513), .B1(new_n457), .B2(new_n454), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n510), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n476), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(KEYINPUT92), .Z(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n523));
  INV_X1    g322(.A(G8gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(KEYINPUT16), .A3(new_n526), .ZN(new_n528));
  AOI211_X1 g327(.A(new_n523), .B(new_n524), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n523), .A2(new_n524), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n527), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n522), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(new_n528), .A3(new_n531), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT91), .A3(G8gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(KEYINPUT93), .A3(new_n532), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT87), .B1(G29gat), .B2(G36gat), .ZN(new_n539));
  INV_X1    g338(.A(G29gat), .ZN(new_n540));
  INV_X1    g339(.A(G36gat), .ZN(new_n541));
  OAI22_X1  g340(.A1(new_n539), .A2(KEYINPUT14), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n539), .A2(KEYINPUT14), .ZN(new_n543));
  OR3_X1    g342(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT88), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n546), .B2(KEYINPUT15), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n547), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n546), .A2(new_n549), .A3(KEYINPUT15), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n545), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n551), .A2(new_n545), .A3(KEYINPUT89), .A4(new_n552), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(KEYINPUT17), .A3(new_n556), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n529), .B2(new_n533), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n555), .B2(new_n556), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n521), .B(new_n558), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT18), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n563), .A2(KEYINPUT94), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(new_n563), .B2(KEYINPUT94), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n520), .B(KEYINPUT13), .Z(new_n567));
  OR2_X1    g366(.A1(new_n538), .A2(new_n557), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n567), .B1(new_n568), .B2(new_n558), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n565), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G113gat), .B(G141gat), .Z(new_n571));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT12), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n563), .A2(KEYINPUT94), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n569), .B1(new_n578), .B2(KEYINPUT18), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT94), .A3(new_n564), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n576), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n518), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n561), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n557), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT102), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G99gat), .B(G106gat), .Z(new_n598));
  OAI21_X1  g397(.A(new_n590), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n600), .A2(KEYINPUT102), .A3(new_n592), .A4(new_n596), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n559), .A3(new_n604), .ZN(new_n605));
  AND3_X1   g404(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n604), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n557), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n587), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT101), .Z(new_n612));
  XNOR2_X1  g411(.A(G134gat), .B(G162gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  NAND3_X1  g413(.A1(new_n605), .A2(new_n587), .A3(new_n608), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT103), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n609), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n605), .A2(KEYINPUT103), .A3(new_n587), .A4(new_n608), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n614), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI211_X1 g421(.A(KEYINPUT104), .B(new_n614), .C1(new_n618), .C2(new_n619), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n616), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(KEYINPUT105), .B(new_n616), .C1(new_n622), .C2(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n629));
  INV_X1    g428(.A(G57gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(G64gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(G64gat), .ZN(new_n632));
  INV_X1    g431(.A(G64gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(KEYINPUT96), .A3(G57gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT97), .ZN(new_n636));
  XOR2_X1   g435(.A(G71gat), .B(G78gat), .Z(new_n637));
  AOI21_X1  g436(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n633), .A2(G57gat), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT95), .B1(new_n632), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n638), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n632), .A2(new_n641), .A3(KEYINPUT95), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n637), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n538), .B1(KEYINPUT21), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT100), .ZN(new_n650));
  XNOR2_X1  g449(.A(G127gat), .B(G155gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT20), .ZN(new_n652));
  NAND2_X1  g451(.A1(G231gat), .A2(G233gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT98), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n650), .B(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n648), .A2(KEYINPUT21), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT99), .B(KEYINPUT19), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(G183gat), .B(G211gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n656), .A2(new_n661), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n628), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n598), .B(KEYINPUT106), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n597), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n602), .A2(new_n640), .A3(new_n646), .A4(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n671), .B(new_n672), .C1(new_n607), .C2(new_n648), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n607), .A2(new_n648), .A3(KEYINPUT10), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n668), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n671), .B1(new_n607), .B2(new_n648), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n668), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G120gat), .B(G148gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  OR2_X1    g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n585), .A2(new_n666), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n468), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  INV_X1    g486(.A(new_n464), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT107), .B(KEYINPUT16), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G8gat), .ZN(new_n692));
  OR3_X1    g491(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(G8gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n690), .B1(new_n689), .B2(new_n692), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT108), .ZN(G1325gat));
  INV_X1    g496(.A(G15gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n471), .A2(new_n473), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT109), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n451), .A2(new_n446), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT70), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n451), .A2(new_n449), .A3(new_n446), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n438), .B1(new_n707), .B2(new_n448), .ZN(new_n708));
  INV_X1    g507(.A(new_n454), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT36), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n471), .A2(new_n513), .A3(new_n473), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n703), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n702), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n684), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n701), .B1(new_n715), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g515(.A1(new_n684), .A2(new_n511), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT43), .B(G22gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  AND2_X1   g518(.A1(new_n626), .A2(new_n627), .ZN(new_n720));
  INV_X1    g519(.A(new_n584), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n665), .A2(new_n683), .A3(new_n721), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n518), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n540), .A3(new_n685), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT45), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n720), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n310), .B1(new_n467), .B2(new_n395), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT110), .B1(new_n460), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT110), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n397), .A2(new_n730), .A3(new_n511), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(new_n713), .A3(new_n510), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n727), .B1(new_n733), .B2(new_n476), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n726), .B1(new_n518), .B2(new_n720), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n722), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT111), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n738), .B(new_n722), .C1(new_n734), .C2(new_n735), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n737), .A2(new_n685), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n725), .B1(new_n740), .B2(new_n540), .ZN(G1328gat));
  NAND3_X1  g540(.A1(new_n723), .A2(new_n541), .A3(new_n688), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT46), .Z(new_n743));
  AND3_X1   g542(.A1(new_n737), .A2(new_n688), .A3(new_n739), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n541), .ZN(G1329gat));
  OAI21_X1  g544(.A(G43gat), .B1(new_n736), .B2(new_n713), .ZN(new_n746));
  INV_X1    g545(.A(G43gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n723), .A2(new_n747), .A3(new_n700), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(KEYINPUT47), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n748), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n737), .A2(new_n714), .A3(new_n739), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(G43gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n752), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g552(.A(G50gat), .B1(new_n736), .B2(new_n460), .ZN(new_n754));
  INV_X1    g553(.A(G50gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n723), .A2(new_n755), .A3(new_n511), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(KEYINPUT48), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n737), .A2(new_n511), .A3(new_n739), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G50gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n756), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n759), .B2(G50gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n765), .A2(KEYINPUT112), .A3(KEYINPUT48), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n757), .B1(new_n763), .B2(new_n766), .ZN(G1331gat));
  NAND2_X1  g566(.A1(new_n733), .A2(new_n476), .ZN(new_n768));
  INV_X1    g567(.A(new_n683), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n666), .A2(new_n769), .A3(new_n584), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n685), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n688), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT49), .B(G64gat), .Z(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(G1333gat));
  NAND2_X1  g576(.A1(new_n771), .A2(new_n714), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n699), .A2(G71gat), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n778), .A2(G71gat), .B1(new_n771), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g580(.A1(new_n771), .A2(new_n511), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n720), .A3(new_n664), .A4(new_n721), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n786), .A2(new_n594), .A3(new_n685), .A4(new_n683), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n734), .A2(new_n735), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n665), .A2(new_n769), .A3(new_n584), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n791), .B2(new_n468), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G85gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n791), .A2(new_n788), .A3(new_n468), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n787), .B1(new_n793), .B2(new_n794), .ZN(G1336gat));
  NAND3_X1  g594(.A1(new_n789), .A2(new_n688), .A3(new_n790), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT114), .B1(new_n796), .B2(G92gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(KEYINPUT52), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n464), .A2(G92gat), .A3(new_n769), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n786), .A2(new_n799), .B1(new_n796), .B2(G92gat), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n798), .B(new_n800), .ZN(G1337gat));
  NOR3_X1   g600(.A1(new_n769), .A2(new_n699), .A3(G99gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G99gat), .B1(new_n791), .B2(new_n713), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1338gat));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n511), .A3(new_n790), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G106gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n460), .A2(G106gat), .A3(new_n769), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n786), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT115), .B1(new_n786), .B2(new_n808), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT53), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n806), .A2(KEYINPUT116), .ZN(new_n815));
  OAI21_X1  g614(.A(G106gat), .B1(new_n806), .B2(KEYINPUT116), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n814), .B(new_n809), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n813), .A2(new_n817), .ZN(G1339gat));
  NOR2_X1   g617(.A1(new_n688), .A2(new_n468), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n673), .A2(new_n674), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n667), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n673), .A2(new_n668), .A3(new_n674), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n680), .B1(new_n675), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n682), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT55), .B1(new_n824), .B2(new_n826), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n558), .B1(new_n560), .B2(new_n562), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n520), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n568), .A2(new_n558), .A3(new_n567), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n575), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(new_n570), .B2(new_n576), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n626), .A2(new_n627), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n584), .A2(new_n830), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n683), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n626), .A2(new_n627), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n664), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n628), .A2(new_n665), .A3(new_n769), .A4(new_n721), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n820), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n511), .A2(new_n699), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n353), .A3(new_n721), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n468), .B1(new_n841), .B2(new_n842), .ZN(new_n847));
  INV_X1    g646(.A(new_n458), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n688), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n584), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n846), .B1(new_n851), .B2(new_n353), .ZN(G1340gat));
  NOR3_X1   g651(.A1(new_n845), .A2(new_n356), .A3(new_n769), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n683), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n356), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n349), .A3(new_n665), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n845), .B2(new_n664), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1342gat));
  NAND2_X1  g657(.A1(new_n720), .A2(new_n464), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT117), .Z(new_n860));
  NOR3_X1   g659(.A1(new_n849), .A2(new_n860), .A3(G134gat), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n845), .B2(new_n628), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(KEYINPUT56), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G1343gat));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n460), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT119), .B1(new_n828), .B2(new_n829), .ZN(new_n869));
  INV_X1    g668(.A(new_n829), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n682), .A4(new_n827), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n584), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n839), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n628), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n837), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n626), .A2(new_n627), .B1(new_n873), .B2(new_n839), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT120), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n665), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n842), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n868), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n460), .B1(new_n841), .B2(new_n842), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT118), .B1(new_n883), .B2(KEYINPUT57), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n838), .A2(new_n839), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n628), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n626), .A2(new_n627), .A3(new_n836), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n665), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n511), .B1(new_n888), .B2(new_n881), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n867), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n882), .A2(new_n884), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n714), .A2(new_n820), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n584), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G141gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n714), .A2(new_n460), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n843), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n721), .A2(G141gat), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT121), .Z(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT58), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n895), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1344gat));
  INV_X1    g704(.A(G148gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n897), .A2(new_n906), .A3(new_n683), .ZN(new_n907));
  XOR2_X1   g706(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n908));
  OAI21_X1  g707(.A(new_n868), .B1(new_n888), .B2(new_n881), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n664), .B1(new_n837), .B2(new_n878), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n460), .B1(new_n910), .B2(new_n842), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n911), .B2(KEYINPUT57), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n683), .A3(new_n893), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n906), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n908), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n906), .A2(KEYINPUT59), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n892), .A2(new_n893), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n683), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n907), .B1(new_n917), .B2(new_n920), .ZN(G1345gat));
  NAND3_X1  g720(.A1(new_n892), .A2(new_n665), .A3(new_n893), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G155gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n897), .A2(new_n316), .A3(new_n665), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n923), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(G1346gat));
  INV_X1    g728(.A(new_n860), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n930), .A2(new_n325), .A3(new_n847), .A4(new_n896), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n919), .A2(new_n720), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n325), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n685), .A2(new_n464), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n935), .B1(new_n841), .B2(new_n842), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n844), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n205), .A3(new_n721), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n936), .A2(new_n848), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT125), .Z(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n584), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n938), .B1(new_n941), .B2(new_n205), .ZN(G1348gat));
  NAND3_X1  g741(.A1(new_n940), .A2(new_n206), .A3(new_n683), .ZN(new_n943));
  OAI21_X1  g742(.A(G176gat), .B1(new_n937), .B2(new_n769), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1349gat));
  NAND2_X1  g744(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n939), .A2(new_n665), .A3(new_n946), .A4(new_n224), .ZN(new_n947));
  OAI21_X1  g746(.A(G183gat), .B1(new_n937), .B2(new_n664), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g749(.A(G190gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n940), .A2(new_n951), .A3(new_n720), .ZN(new_n952));
  XNOR2_X1  g751(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n720), .A3(new_n844), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(G190gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(G190gat), .A3(new_n953), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n952), .B1(new_n955), .B2(new_n957), .ZN(G1351gat));
  NOR2_X1   g757(.A1(new_n714), .A2(new_n935), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n912), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(G197gat), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n721), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n883), .A2(new_n584), .A3(new_n959), .ZN(new_n963));
  AOI22_X1  g762(.A1(new_n960), .A2(new_n962), .B1(new_n961), .B2(new_n963), .ZN(G1352gat));
  NAND2_X1  g763(.A1(new_n883), .A2(new_n959), .ZN(new_n965));
  INV_X1    g764(.A(G204gat), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(KEYINPUT127), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n965), .A2(new_n769), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(KEYINPUT127), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n969), .B(new_n970), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n912), .A2(new_n683), .A3(new_n959), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n972), .B2(new_n966), .ZN(G1353gat));
  NAND2_X1  g772(.A1(new_n960), .A2(new_n665), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n665), .A2(new_n260), .ZN(new_n977));
  OAI22_X1  g776(.A1(new_n975), .A2(new_n976), .B1(new_n965), .B2(new_n977), .ZN(G1354gat));
  AND2_X1   g777(.A1(new_n960), .A2(new_n720), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n720), .A2(new_n261), .ZN(new_n980));
  OAI22_X1  g779(.A1(new_n979), .A2(new_n261), .B1(new_n965), .B2(new_n980), .ZN(G1355gat));
endmodule


