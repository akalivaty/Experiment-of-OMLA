//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G214), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G131), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT17), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(new_n195), .A3(new_n191), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(KEYINPUT17), .A3(G131), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT76), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT76), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(G125), .A2(G140), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n205), .B2(G140), .ZN(new_n210));
  OAI211_X1 g024(.A(G146), .B(new_n208), .C1(new_n210), .C2(new_n206), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n209), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT76), .B(G125), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(new_n207), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT16), .ZN(new_n217));
  AOI21_X1  g031(.A(G146), .B1(new_n217), .B2(new_n208), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n203), .A2(G125), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n201), .A2(KEYINPUT76), .ZN(new_n222));
  OAI21_X1  g036(.A(G140), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n206), .B1(new_n223), .B2(new_n214), .ZN(new_n224));
  INV_X1    g038(.A(new_n208), .ZN(new_n225));
  OAI211_X1 g039(.A(KEYINPUT77), .B(new_n220), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n200), .B1(new_n219), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G113), .B(G122), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT87), .B(G104), .ZN(new_n230));
  XOR2_X1   g044(.A(new_n229), .B(new_n230), .Z(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT18), .A2(G131), .ZN(new_n233));
  OR2_X1    g047(.A1(new_n192), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G125), .B(G140), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n220), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n216), .B2(new_n220), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n192), .A2(new_n233), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n228), .A2(new_n232), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n220), .B1(new_n224), .B2(new_n225), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n212), .A3(new_n211), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n199), .B1(new_n242), .B2(new_n226), .ZN(new_n243));
  INV_X1    g057(.A(new_n239), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n231), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G902), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G475), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G475), .A2(G902), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n243), .A2(new_n231), .A3(new_n244), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n210), .A2(KEYINPUT19), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(KEYINPUT86), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT19), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n235), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT86), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(KEYINPUT19), .B2(new_n210), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n220), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n193), .A2(new_n196), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n211), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n232), .B1(new_n263), .B2(new_n239), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n252), .A2(new_n264), .A3(KEYINPUT88), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n253), .A2(KEYINPUT86), .A3(new_n256), .ZN(new_n267));
  OR3_X1    g081(.A1(new_n216), .A2(KEYINPUT86), .A3(new_n255), .ZN(new_n268));
  AOI21_X1  g082(.A(G146), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n239), .B1(new_n269), .B2(new_n261), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n231), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n266), .B1(new_n240), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n251), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT20), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT20), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n275), .B(new_n251), .C1(new_n252), .C2(new_n264), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n250), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT9), .B(G234), .ZN(new_n278));
  OAI21_X1  g092(.A(G221), .B1(new_n278), .B2(G902), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G137), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G134), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT11), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT11), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT66), .ZN(new_n286));
  OAI211_X1 g100(.A(KEYINPUT67), .B(new_n282), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G134), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(G137), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n283), .A2(KEYINPUT11), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n281), .A2(KEYINPUT11), .A3(G134), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n287), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n288), .A2(G137), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G131), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n300));
  AOI21_X1  g114(.A(G131), .B1(new_n288), .B2(G137), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n300), .B1(new_n296), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(G104), .B(G107), .ZN(new_n305));
  INV_X1    g119(.A(G101), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT79), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G107), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G104), .ZN(new_n309));
  INV_X1    g123(.A(G104), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G107), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(G101), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n310), .B2(G107), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n308), .A3(G104), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n315), .A2(new_n317), .A3(new_n306), .A4(new_n311), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n307), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G128), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(KEYINPUT1), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n220), .A2(G143), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n189), .A2(G146), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n220), .B2(G143), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n189), .A2(KEYINPUT65), .A3(G146), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n326), .A2(new_n327), .B1(G143), .B2(new_n220), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n320), .B1(new_n322), .B2(KEYINPUT1), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n319), .B(new_n324), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n322), .B2(new_n323), .ZN(new_n331));
  INV_X1    g145(.A(new_n324), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n330), .B1(new_n333), .B2(new_n319), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n304), .A2(new_n334), .A3(KEYINPUT12), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT82), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n304), .A2(new_n334), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT12), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n304), .A2(new_n334), .A3(KEYINPUT82), .A4(KEYINPUT12), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n333), .B2(new_n319), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT10), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n347), .B2(new_n319), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT0), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n320), .A3(KEYINPUT64), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT64), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n351), .B1(KEYINPUT0), .B2(G128), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(KEYINPUT0), .A2(G128), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n322), .A2(new_n323), .ZN(new_n356));
  OAI22_X1  g170(.A1(new_n355), .A2(new_n328), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n315), .A2(new_n317), .A3(new_n311), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G101), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(KEYINPUT4), .A3(new_n318), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n362), .A3(G101), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n319), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n365), .A2(KEYINPUT80), .A3(KEYINPUT10), .A4(new_n346), .ZN(new_n366));
  AND4_X1   g180(.A1(new_n344), .A2(new_n348), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n195), .B1(new_n296), .B2(new_n297), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n290), .A2(new_n291), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n295), .B1(new_n282), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n371), .A2(new_n294), .A3(new_n289), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n301), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT68), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n368), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n299), .B(new_n377), .C1(new_n302), .C2(new_n303), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n367), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n342), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G140), .ZN(new_n383));
  INV_X1    g197(.A(G227), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G953), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n383), .B(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n364), .A2(new_n348), .A3(new_n366), .A4(new_n344), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n304), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n304), .A2(KEYINPUT81), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n379), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n390), .B2(new_n367), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n382), .A2(new_n386), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G469), .B1(new_n392), .B2(G902), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n342), .A2(new_n391), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n387), .B1(new_n389), .B2(new_n379), .ZN(new_n395));
  INV_X1    g209(.A(new_n388), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n386), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G469), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT74), .B(G902), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n280), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n400), .ZN(new_n403));
  INV_X1    g217(.A(G217), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n278), .A2(new_n404), .A3(G953), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G122), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G116), .ZN(new_n408));
  INV_X1    g222(.A(G116), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G122), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(new_n308), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n189), .A2(G128), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT13), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n320), .A2(G143), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT89), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT89), .B1(new_n320), .B2(G143), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G134), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n416), .B(new_n417), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n288), .A4(new_n413), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n288), .B(new_n413), .C1(new_n418), .C2(new_n419), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT90), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n412), .A2(new_n421), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n410), .A2(KEYINPUT14), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT14), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n409), .A3(G122), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n428), .A2(new_n430), .A3(KEYINPUT91), .A4(new_n408), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n431), .B(G107), .C1(KEYINPUT91), .C2(new_n430), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n411), .A2(new_n308), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n288), .B1(new_n422), .B2(new_n413), .ZN(new_n434));
  INV_X1    g248(.A(new_n425), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n432), .B(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n427), .A2(new_n436), .A3(KEYINPUT92), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT92), .B1(new_n427), .B2(new_n436), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n406), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n439), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n405), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n403), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n443), .B(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G953), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n449), .A2(G952), .ZN(new_n450));
  INV_X1    g264(.A(G234), .ZN(new_n451));
  INV_X1    g265(.A(G237), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n449), .B(new_n400), .C1(G234), .C2(G237), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(G898), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G210), .B1(G237), .B2(G902), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n357), .A2(new_n205), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n324), .B(new_n215), .C1(new_n328), .C2(new_n329), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT84), .ZN(new_n463));
  INV_X1    g277(.A(G224), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT84), .B1(new_n357), .B2(new_n205), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n463), .A2(KEYINPUT7), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G119), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G116), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n409), .A2(G119), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT2), .B(G113), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT5), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G113), .B1(new_n471), .B2(KEYINPUT5), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n365), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n473), .A2(new_n474), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n361), .A2(new_n482), .A3(new_n363), .ZN(new_n483));
  XNOR2_X1  g297(.A(G110), .B(G122), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n460), .B2(new_n461), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT7), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n466), .A2(new_n490), .ZN(new_n491));
  OAI22_X1  g305(.A1(new_n487), .A2(new_n467), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n319), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n480), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n484), .B(KEYINPUT8), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n469), .A2(new_n485), .A3(new_n492), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n247), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n485), .A2(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n480), .A2(new_n483), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT83), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n484), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(KEYINPUT6), .A3(new_n503), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n465), .B1(new_n487), .B2(new_n467), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n459), .B1(new_n499), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n485), .A2(KEYINPUT6), .B1(new_n501), .B2(new_n503), .ZN(new_n512));
  INV_X1    g326(.A(new_n506), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(new_n247), .A3(new_n458), .A4(new_n498), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n448), .B(new_n457), .C1(new_n510), .C2(new_n515), .ZN(new_n516));
  AND4_X1   g330(.A1(new_n277), .A2(new_n402), .A3(new_n446), .A4(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n376), .A2(new_n519), .A3(new_n357), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT69), .B1(new_n304), .B2(new_n358), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n282), .A2(new_n297), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G131), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n346), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n302), .B2(new_n303), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(KEYINPUT70), .B(new_n525), .C1(new_n302), .C2(new_n303), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n518), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n304), .A2(new_n358), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT30), .A3(new_n526), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n482), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n482), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n526), .B(new_n537), .C1(new_n376), .C2(new_n357), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT26), .B(G101), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT72), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n187), .A2(G210), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(G210), .A3(new_n187), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n536), .A2(new_n538), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n400), .B1(new_n550), .B2(KEYINPUT29), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n538), .A2(KEYINPUT28), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n532), .A2(new_n553), .A3(new_n526), .A4(new_n537), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n537), .B1(new_n532), .B2(new_n526), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT29), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT29), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n519), .B1(new_n376), .B2(new_n357), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n304), .A2(KEYINPUT69), .A3(new_n358), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n530), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n555), .B(new_n560), .C1(new_n563), .C2(new_n537), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n559), .A2(new_n548), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G472), .B1(new_n551), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n561), .A2(new_n562), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n374), .A2(new_n375), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT70), .B1(new_n570), .B2(new_n525), .ZN(new_n571));
  INV_X1    g385(.A(new_n529), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT30), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT73), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n538), .A2(new_n575), .A3(new_n548), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n538), .B2(new_n548), .ZN(new_n577));
  OAI22_X1  g391(.A1(new_n574), .A2(new_n534), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n555), .B1(new_n563), .B2(new_n537), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n578), .A2(KEYINPUT31), .B1(new_n579), .B2(new_n549), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  OAI221_X1 g395(.A(new_n581), .B1(new_n576), .B2(new_n577), .C1(new_n574), .C2(new_n534), .ZN(new_n582));
  AOI211_X1 g396(.A(KEYINPUT32), .B(new_n568), .C1(new_n580), .C2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT32), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n569), .A2(new_n573), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n534), .B1(new_n585), .B2(new_n518), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n576), .A2(new_n577), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT31), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n579), .A2(new_n549), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n582), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n584), .B1(new_n590), .B2(new_n567), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n566), .B1(new_n583), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n404), .B1(new_n400), .B2(G234), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n211), .A2(new_n236), .ZN(new_n595));
  XNOR2_X1  g409(.A(G119), .B(G128), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT75), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT24), .B(G110), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT23), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n470), .B2(G128), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n320), .A2(KEYINPUT23), .A3(G119), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n601), .B(new_n602), .C1(G119), .C2(new_n320), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n603), .A2(G110), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n599), .A2(KEYINPUT78), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT78), .B1(new_n599), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n595), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n597), .ZN(new_n608));
  INV_X1    g422(.A(new_n598), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n608), .A2(new_n609), .B1(G110), .B2(new_n603), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n242), .A2(new_n610), .A3(new_n226), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT22), .B(G137), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n449), .A2(G221), .A3(G234), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n612), .B(new_n613), .Z(new_n614));
  AND3_X1   g428(.A1(new_n607), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n607), .B2(new_n611), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(KEYINPUT25), .A3(new_n400), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n607), .A2(new_n611), .ZN(new_n619));
  INV_X1    g433(.A(new_n614), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n607), .A2(new_n611), .A3(new_n614), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n400), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT25), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n594), .B1(new_n618), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n617), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n593), .A2(G902), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n517), .A2(new_n592), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  INV_X1    g447(.A(G472), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n590), .B2(new_n400), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n567), .B2(new_n590), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n631), .A3(new_n402), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT93), .ZN(new_n638));
  INV_X1    g452(.A(new_n251), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT88), .B1(new_n252), .B2(new_n264), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n240), .A2(new_n266), .A3(new_n271), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n276), .B1(new_n642), .B2(new_n275), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n249), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n427), .A2(new_n436), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n405), .A2(KEYINPUT95), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n440), .A2(new_n442), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(G478), .A3(new_n400), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n400), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(KEYINPUT96), .A3(new_n444), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n443), .B2(G478), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n644), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n510), .A2(KEYINPUT94), .A3(new_n515), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT94), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n661), .B(new_n459), .C1(new_n499), .C2(new_n509), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n447), .A3(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n659), .A2(new_n457), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n638), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT34), .B(G104), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G6));
  INV_X1    g481(.A(KEYINPUT97), .ZN(new_n668));
  INV_X1    g482(.A(new_n445), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n443), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n640), .A2(new_n641), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n275), .B1(new_n671), .B2(new_n251), .ZN(new_n672));
  AOI211_X1 g486(.A(KEYINPUT20), .B(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n670), .B(new_n249), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n668), .B1(new_n674), .B2(new_n457), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n642), .A2(new_n275), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n250), .B1(new_n274), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n457), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n677), .A2(KEYINPUT97), .A3(new_n670), .A4(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n663), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n675), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n638), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT98), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT35), .B(G107), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G9));
  NAND2_X1  g499(.A1(new_n618), .A2(new_n625), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n593), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n620), .A2(KEYINPUT36), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n619), .B(new_n688), .Z(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n629), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n687), .A2(KEYINPUT99), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT99), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n626), .B2(new_n690), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n517), .A2(new_n636), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT37), .B(G110), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G12));
  AND3_X1   g512(.A1(new_n695), .A2(new_n402), .A3(new_n680), .ZN(new_n699));
  INV_X1    g513(.A(G900), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n454), .B1(new_n455), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n674), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n699), .A2(new_n592), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  INV_X1    g518(.A(new_n695), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n510), .A2(new_n515), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT38), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n447), .A3(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n708), .A2(new_n277), .A3(new_n446), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n701), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n402), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT40), .Z(new_n712));
  INV_X1    g526(.A(new_n577), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n538), .A2(new_n575), .A3(new_n548), .ZN(new_n714));
  AOI22_X1  g528(.A1(new_n531), .A2(new_n535), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n548), .B1(new_n557), .B2(new_n538), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n247), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G472), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n583), .B2(new_n591), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n709), .A2(new_n712), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  INV_X1    g535(.A(new_n701), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n644), .A2(new_n658), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n699), .A2(new_n592), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  NAND2_X1  g540(.A1(new_n381), .A2(new_n388), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n386), .A2(new_n727), .B1(new_n342), .B2(new_n391), .ZN(new_n728));
  OAI21_X1  g542(.A(G469), .B1(new_n728), .B2(new_n403), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(KEYINPUT100), .A3(new_n401), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT100), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n731), .B(G469), .C1(new_n728), .C2(new_n403), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n280), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n592), .A2(new_n733), .A3(new_n631), .A4(new_n664), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT101), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND4_X1  g551(.A1(new_n681), .A2(new_n592), .A3(new_n631), .A4(new_n733), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  AOI211_X1 g553(.A(new_n280), .B(new_n663), .C1(new_n732), .C2(new_n730), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n644), .A2(new_n670), .A3(new_n457), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n592), .A2(new_n740), .A3(new_n695), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  AOI211_X1 g557(.A(KEYINPUT104), .B(new_n446), .C1(new_n643), .C2(new_n249), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n644), .B2(new_n670), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n740), .A2(new_n747), .A3(new_n678), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n556), .B1(new_n552), .B2(new_n554), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT102), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n549), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI211_X1 g565(.A(KEYINPUT102), .B(new_n556), .C1(new_n552), .C2(new_n554), .ZN(new_n752));
  OAI22_X1  g566(.A1(new_n715), .A2(new_n581), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT103), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n582), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n558), .A2(KEYINPUT102), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n749), .A2(new_n750), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n549), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT103), .B1(new_n758), .B2(new_n588), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n567), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n635), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n631), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT105), .B1(new_n748), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n631), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n753), .A2(new_n754), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n758), .A2(KEYINPUT103), .A3(new_n588), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n582), .A3(new_n766), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n764), .B(new_n635), .C1(new_n767), .C2(new_n567), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n730), .A2(new_n732), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n279), .A3(new_n678), .A4(new_n680), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT104), .B1(new_n277), .B2(new_n446), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n644), .A2(new_n745), .A3(new_n670), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n768), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n763), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G122), .ZN(G24));
  AOI21_X1  g592(.A(new_n635), .B1(new_n767), .B2(new_n567), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n695), .A3(new_n724), .A4(new_n740), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G125), .ZN(G27));
  INV_X1    g595(.A(new_n591), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n590), .A2(new_n584), .A3(new_n567), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT107), .B1(new_n583), .B2(new_n591), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n786), .A3(new_n566), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n706), .A2(new_n448), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n391), .A2(new_n388), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n342), .A2(new_n381), .ZN(new_n790));
  INV_X1    g604(.A(new_n386), .ZN(new_n791));
  OAI211_X1 g605(.A(G469), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(G469), .A2(G902), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n401), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n788), .B(new_n279), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n723), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n787), .A2(KEYINPUT42), .A3(new_n631), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n592), .A2(new_n631), .A3(new_n797), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT42), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n799), .A2(KEYINPUT106), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT106), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G131), .ZN(G33));
  INV_X1    g618(.A(new_n592), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n764), .ZN(new_n806));
  INV_X1    g620(.A(new_n796), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n702), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(KEYINPUT108), .B(G134), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(G36));
  INV_X1    g624(.A(new_n788), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n277), .A2(new_n658), .ZN(new_n812));
  AND2_X1   g626(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n813));
  NOR2_X1   g627(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n812), .A2(new_n814), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n705), .B(new_n636), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n811), .B1(new_n817), .B2(KEYINPUT44), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(KEYINPUT44), .B2(new_n817), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n392), .A2(KEYINPUT45), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(G469), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT46), .B1(new_n824), .B2(new_n793), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n795), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(KEYINPUT46), .A3(new_n793), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n279), .A3(new_n710), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n819), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G137), .ZN(G39));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n279), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT47), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n723), .A2(new_n631), .A3(new_n811), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n805), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G140), .ZN(G42));
  AOI21_X1  g651(.A(new_n453), .B1(new_n816), .B2(new_n815), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n707), .A2(new_n447), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n768), .A3(new_n733), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT115), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT50), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT116), .Z(new_n846));
  AND2_X1   g660(.A1(new_n733), .A2(new_n788), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n838), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT117), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n695), .A3(new_n779), .ZN(new_n850));
  INV_X1    g664(.A(new_n719), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n631), .A3(new_n454), .A4(new_n847), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n852), .A2(new_n644), .A3(new_n658), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n832), .B(KEYINPUT47), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n834), .A2(KEYINPUT114), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n769), .A2(new_n280), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n838), .A2(new_n768), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n811), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n854), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT51), .B1(new_n846), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n855), .A2(new_n859), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n862), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(KEYINPUT51), .A3(new_n850), .A4(new_n853), .ZN(new_n867));
  INV_X1    g681(.A(new_n740), .ZN(new_n868));
  OAI221_X1 g682(.A(new_n450), .B1(new_n852), .B2(new_n659), .C1(new_n868), .C2(new_n861), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n787), .A2(new_n631), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n849), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT48), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT48), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n849), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n869), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n867), .A2(new_n845), .B1(new_n875), .B2(KEYINPUT118), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n864), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n699), .B(new_n592), .C1(new_n702), .C2(new_n724), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n744), .A2(new_n746), .A3(new_n663), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n626), .A2(new_n690), .A3(new_n701), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n402), .A3(new_n719), .A4(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n780), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT52), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n880), .A2(new_n780), .A3(new_n883), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(KEYINPUT111), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n738), .A2(new_n734), .A3(new_n742), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n776), .B2(new_n763), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n670), .B(KEYINPUT110), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n277), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n659), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n402), .A2(new_n516), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n636), .A3(new_n631), .A4(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n895), .A2(new_n632), .A3(new_n696), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n890), .A2(new_n885), .A3(new_n887), .A4(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n779), .A2(new_n724), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n891), .A2(new_n701), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n592), .A2(new_n677), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n695), .B(new_n807), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n803), .A2(new_n808), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n879), .B(new_n888), .C1(new_n897), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n885), .A2(new_n887), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n738), .A2(new_n734), .A3(new_n742), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n777), .A3(new_n896), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n888), .A2(new_n879), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n803), .A2(new_n808), .A3(new_n901), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT113), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n885), .A2(KEYINPUT53), .A3(new_n887), .A4(new_n896), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n748), .A2(new_n762), .A3(KEYINPUT105), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n775), .B1(new_n768), .B2(new_n774), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT112), .B1(new_n918), .B2(new_n889), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT112), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n905), .A2(new_n777), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n915), .A2(new_n909), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n879), .B1(new_n897), .B2(new_n902), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n912), .A2(new_n913), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n925), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n903), .B2(new_n910), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT113), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n878), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(G952), .B2(G953), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n769), .B(KEYINPUT49), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n631), .A2(new_n279), .A3(new_n447), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n933), .A2(new_n707), .A3(new_n812), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n851), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n931), .A2(new_n935), .ZN(G75));
  NOR2_X1   g750(.A1(new_n449), .A2(G952), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n400), .B1(new_n922), .B2(new_n923), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT56), .B1(new_n938), .B2(new_n459), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n505), .A2(new_n506), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n511), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT55), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n937), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n919), .A2(new_n921), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n945), .A2(new_n902), .A3(new_n914), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT53), .B1(new_n907), .B2(new_n909), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n403), .B(new_n459), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT119), .B1(new_n950), .B2(new_n942), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT119), .ZN(new_n952));
  AOI211_X1 g766(.A(new_n952), .B(new_n943), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n944), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT120), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(KEYINPUT120), .B(new_n944), .C1(new_n951), .C2(new_n953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(G51));
  OAI21_X1  g772(.A(KEYINPUT54), .B1(new_n946), .B2(new_n947), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(KEYINPUT121), .A3(new_n925), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n922), .A2(new_n923), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT54), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n793), .B(KEYINPUT57), .Z(new_n964));
  NAND3_X1  g778(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n398), .ZN(new_n966));
  AOI211_X1 g780(.A(new_n400), .B(new_n824), .C1(new_n922), .C2(new_n923), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT122), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n937), .B1(new_n966), .B2(new_n968), .ZN(G54));
  NAND3_X1  g783(.A1(new_n938), .A2(KEYINPUT58), .A3(G475), .ZN(new_n970));
  INV_X1    g784(.A(new_n671), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n972), .A2(new_n973), .A3(new_n937), .ZN(G60));
  NAND2_X1  g788(.A1(G478), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT59), .Z(new_n976));
  AOI211_X1 g790(.A(new_n976), .B(new_n649), .C1(new_n648), .C2(new_n650), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n960), .A2(new_n963), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n937), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n976), .B1(new_n929), .B2(new_n926), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n651), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n980), .A2(new_n983), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT60), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n961), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n937), .B1(new_n987), .B2(new_n627), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n689), .B2(new_n987), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g804(.A(G953), .B1(new_n456), .B2(new_n464), .ZN(new_n991));
  INV_X1    g805(.A(new_n906), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(G953), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n505), .B(new_n506), .C1(G898), .C2(new_n449), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(G69));
  NAND2_X1  g809(.A1(new_n531), .A2(new_n533), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n267), .A2(new_n268), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(G900), .B2(G953), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n880), .A2(new_n780), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n836), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n870), .A2(new_n881), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n829), .B1(new_n819), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n803), .A2(new_n808), .ZN(new_n1004));
  OR3_X1    g818(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n999), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n711), .A2(new_n811), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n806), .A2(new_n893), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n830), .A2(new_n836), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n720), .A2(new_n1000), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT62), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n449), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n998), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1006), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(G953), .B1(new_n384), .B2(new_n700), .ZN(new_n1015));
  INV_X1    g829(.A(new_n998), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(new_n1016), .B2(KEYINPUT124), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1014), .B(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(new_n536), .A2(new_n538), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n1009), .A2(new_n906), .A3(new_n1011), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n548), .B(new_n1019), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(KEYINPUT127), .B1(new_n1019), .B2(new_n549), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1025), .A2(new_n715), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1019), .A2(KEYINPUT127), .A3(new_n549), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n911), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1022), .B1(new_n1005), .B2(new_n906), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n550), .B(KEYINPUT125), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n937), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT126), .ZN(new_n1034));
  OR2_X1    g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1030), .B1(new_n1035), .B2(new_n1036), .ZN(G57));
endmodule


