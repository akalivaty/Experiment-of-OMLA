//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  INV_X1    g0006(.A(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n202), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G116), .C2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G1), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT66), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n223), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n232), .A2(new_n221), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n226), .A2(new_n230), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G58), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(new_n213), .ZN(new_n255));
  OAI21_X1  g0055(.A(G20), .B1(new_n255), .B2(new_n201), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G159), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT82), .B1(new_n261), .B2(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n261), .A2(KEYINPUT82), .A3(G33), .ZN(new_n265));
  AOI21_X1  g0065(.A(G20), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  OAI21_X1  g0067(.A(G68), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n261), .A2(KEYINPUT82), .A3(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n263), .B2(new_n262), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n270), .A2(KEYINPUT7), .A3(G20), .ZN(new_n271));
  OAI211_X1 g0071(.A(KEYINPUT16), .B(new_n260), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n233), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT16), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n267), .B1(new_n276), .B2(G20), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n263), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n213), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n275), .B1(new_n282), .B2(new_n259), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n272), .A2(new_n274), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n220), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT72), .ZN(new_n286));
  INV_X1    g0086(.A(new_n285), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n274), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n220), .A2(G20), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(new_n289), .C1(new_n286), .C2(new_n274), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  MUX2_X1   g0092(.A(new_n285), .B(new_n290), .S(new_n292), .Z(new_n293));
  AND2_X1   g0093(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G200), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n212), .A2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G223), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n264), .A2(new_n265), .A3(new_n296), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT83), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G87), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  OAI211_X1 g0105(.A(G1), .B(G13), .C1(new_n278), .C2(new_n305), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G45), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT69), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G45), .ZN(new_n311));
  AOI21_X1  g0111(.A(G41), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT70), .B1(new_n312), .B2(G1), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n306), .A2(G274), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT70), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT69), .B(G45), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n220), .C1(new_n316), .C2(G41), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n220), .B1(G41), .B2(G45), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n306), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G232), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n295), .B1(new_n307), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n300), .A2(new_n302), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT83), .ZN(new_n326));
  INV_X1    g0126(.A(new_n306), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n318), .A2(new_n322), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n294), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT17), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT18), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n307), .A2(new_n337), .A3(new_n323), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n329), .B2(new_n331), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n336), .B1(new_n341), .B2(new_n294), .ZN(new_n342));
  OAI21_X1  g0142(.A(G169), .B1(new_n307), .B2(new_n323), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n329), .A2(G179), .A3(new_n331), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n284), .A2(new_n293), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(KEYINPUT18), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n335), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n321), .A2(G226), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n298), .A2(G222), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n276), .B(new_n351), .C1(new_n297), .C2(new_n298), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n280), .A2(new_n206), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n327), .A3(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n318), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT71), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n318), .A2(KEYINPUT71), .A3(new_n350), .A4(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G190), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n203), .A2(G20), .ZN(new_n361));
  INV_X1    g0161(.A(G150), .ZN(new_n362));
  INV_X1    g0162(.A(new_n257), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n278), .A2(G20), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n361), .B1(new_n362), .B2(new_n363), .C1(new_n365), .C2(new_n291), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n274), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n287), .A2(new_n202), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n367), .B(new_n368), .C1(new_n202), .C2(new_n290), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT9), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n357), .A2(G200), .A3(new_n358), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n369), .A2(new_n370), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n360), .A2(new_n371), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT10), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n369), .A2(new_n370), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(G190), .B2(new_n359), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n371), .A4(new_n372), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n280), .B1(G232), .B2(new_n298), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n214), .B2(new_n298), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n382), .B(new_n327), .C1(G107), .C2(new_n276), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(new_n318), .C1(new_n207), .C2(new_n320), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n384), .A2(G179), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n339), .ZN(new_n386));
  INV_X1    g0186(.A(new_n274), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n289), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(new_n206), .ZN(new_n389));
  XOR2_X1   g0189(.A(KEYINPUT15), .B(G87), .Z(new_n390));
  AOI22_X1  g0190(.A1(new_n292), .A2(new_n257), .B1(new_n390), .B2(new_n364), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n221), .B2(new_n206), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n392), .B2(new_n274), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n285), .A2(G77), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT75), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n385), .A2(new_n386), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n357), .A2(new_n339), .A3(new_n358), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT73), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n398), .A2(new_n399), .A3(new_n369), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n398), .B2(new_n369), .ZN(new_n401));
  AOI211_X1 g0201(.A(KEYINPUT74), .B(G179), .C1(new_n357), .C2(new_n358), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT74), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n359), .B2(new_n337), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n400), .A2(new_n401), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n384), .A2(G200), .ZN(new_n406));
  INV_X1    g0206(.A(new_n396), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(new_n407), .C1(new_n330), .C2(new_n384), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n380), .A2(new_n397), .A3(new_n405), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n212), .A2(new_n298), .ZN(new_n410));
  INV_X1    g0210(.A(G232), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G1698), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n263), .A2(new_n410), .A3(new_n279), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT76), .B1(new_n415), .B2(new_n327), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT76), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n417), .B(new_n306), .C1(new_n413), .C2(new_n414), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n321), .A2(G238), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n318), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT13), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G226), .A2(G1698), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n411), .B2(G1698), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(new_n276), .B1(G33), .B2(G97), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n417), .B1(new_n425), .B2(new_n306), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n415), .A2(KEYINPUT76), .A3(new_n327), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n318), .A4(new_n420), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n430), .A3(KEYINPUT77), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n419), .A2(new_n421), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT77), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n429), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(G200), .A3(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n364), .A2(G77), .B1(G20), .B2(new_n213), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT78), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n202), .B2(new_n363), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n274), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT11), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n287), .A2(KEYINPUT12), .A3(new_n213), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT12), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n285), .B2(G68), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n444), .C1(new_n388), .C2(new_n213), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT79), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n438), .A2(KEYINPUT11), .A3(new_n274), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n441), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n422), .A2(new_n430), .A3(G190), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n435), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT80), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT80), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n435), .A2(new_n448), .A3(new_n452), .A4(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n431), .A2(G169), .A3(new_n434), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT14), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n422), .A2(new_n430), .A3(G179), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT14), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n431), .A2(new_n459), .A3(new_n434), .A4(G169), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n448), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT81), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT81), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n455), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  AOI211_X1 g0267(.A(new_n349), .B(new_n409), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n263), .A2(new_n279), .A3(G250), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n298), .B1(new_n469), .B2(KEYINPUT4), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n298), .A2(KEYINPUT4), .A3(G244), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n280), .A2(new_n473), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n470), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n264), .A2(new_n265), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(new_n207), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n306), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n308), .A2(G1), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  AND2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n480), .B(G274), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n306), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n218), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n339), .B1(new_n479), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n287), .A2(new_n217), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n387), .B(new_n285), .C1(G1), .C2(new_n278), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G97), .ZN(new_n491));
  INV_X1    g0291(.A(G107), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n277), .B2(new_n281), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n363), .A2(new_n206), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n217), .A2(new_n492), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G97), .A2(G107), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n492), .A2(KEYINPUT6), .A3(G97), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n221), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n493), .A2(new_n494), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n488), .B(new_n491), .C1(new_n501), .C2(new_n387), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT84), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n486), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(KEYINPUT84), .B(new_n483), .C1(new_n485), .C2(new_n218), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n276), .A2(KEYINPUT4), .A3(G244), .A4(new_n298), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n476), .B1(new_n276), .B2(G250), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n471), .B(new_n507), .C1(new_n508), .C2(new_n298), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT4), .B1(new_n270), .B2(G244), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n327), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n506), .A2(new_n337), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n487), .A2(new_n502), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT85), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n487), .A2(new_n502), .A3(new_n512), .A4(KEYINPUT85), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n486), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n330), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n295), .B1(new_n506), .B2(new_n511), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n520), .A2(new_n521), .A3(new_n502), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n517), .A2(KEYINPUT86), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(G20), .B1(new_n278), .B2(G97), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n471), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT88), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT88), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n528), .A3(new_n471), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G20), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n527), .A2(new_n529), .A3(new_n274), .A4(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n387), .B1(KEYINPUT88), .B2(new_n526), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(KEYINPUT20), .A3(new_n531), .A4(new_n529), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n285), .A2(G116), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n490), .A2(G116), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G264), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n218), .A2(new_n298), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n264), .A2(new_n265), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G303), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n276), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n327), .ZN(new_n549));
  INV_X1    g0349(.A(new_n485), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G270), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n483), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G200), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n542), .B(new_n553), .C1(new_n330), .C2(new_n552), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n306), .B(G250), .C1(G1), .C2(new_n308), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n207), .A2(G1698), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n214), .A2(new_n298), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n264), .A2(new_n265), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n278), .B2(new_n530), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n556), .B1(new_n560), .B2(new_n327), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n480), .A2(G274), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(G190), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G200), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n270), .A2(new_n221), .A3(G68), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n569), .A2(new_n221), .A3(G33), .A4(G97), .ZN(new_n570));
  NOR3_X1   g0370(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n221), .B2(new_n414), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n570), .B1(new_n572), .B2(new_n569), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n274), .ZN(new_n575));
  INV_X1    g0375(.A(new_n390), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n287), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n490), .A2(G87), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n561), .A2(KEYINPUT87), .A3(G190), .A4(new_n562), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n565), .A2(new_n567), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n566), .A2(new_n339), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n575), .B(new_n577), .C1(new_n576), .C2(new_n489), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(G179), .C2(new_n566), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n287), .A2(new_n492), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n489), .A2(new_n492), .B1(KEYINPUT25), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n208), .A2(G20), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n263), .A3(new_n279), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT22), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT23), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n221), .B2(G107), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n492), .A2(KEYINPUT23), .A3(G20), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n588), .A2(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n264), .A2(KEYINPUT22), .A3(new_n265), .A4(new_n587), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n364), .A2(G116), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g0396(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n593), .A2(new_n594), .A3(new_n597), .A4(new_n595), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n586), .B1(new_n601), .B2(new_n274), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n218), .A2(G1698), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n209), .A2(new_n298), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n264), .A2(new_n265), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G294), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n327), .B1(G264), .B2(new_n550), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n483), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G200), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(G190), .A3(new_n483), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n585), .A2(KEYINPUT25), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n602), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n581), .A2(new_n584), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n524), .A2(new_n554), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n541), .A2(new_n552), .A3(G169), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n552), .A2(new_n337), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n541), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n541), .A2(new_n552), .A3(KEYINPUT21), .A4(G169), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n602), .A2(new_n612), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n609), .A2(new_n339), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n608), .A2(new_n337), .A3(new_n483), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n522), .B1(new_n515), .B2(new_n516), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n624), .B(new_n628), .C1(new_n629), .C2(KEYINPUT86), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n616), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n468), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g0432(.A(new_n632), .B(KEYINPUT90), .Z(G372));
  NAND2_X1  g0433(.A1(new_n581), .A2(new_n584), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n513), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n515), .A2(new_n516), .A3(new_n581), .A4(new_n584), .ZN(new_n636));
  XNOR2_X1  g0436(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI22_X1  g0438(.A1(new_n635), .A2(KEYINPUT26), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n628), .A2(new_n621), .A3(new_n619), .A4(new_n622), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n615), .A2(new_n640), .A3(new_n629), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n584), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n468), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT17), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n334), .B(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n397), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n450), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n463), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT92), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n345), .A2(KEYINPUT18), .A3(new_n346), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT18), .B1(new_n345), .B2(new_n346), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n342), .A2(KEYINPUT92), .A3(new_n347), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n380), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n405), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n643), .A2(new_n657), .ZN(G369));
  INV_X1    g0458(.A(G13), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G20), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n220), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n623), .A2(new_n541), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n666), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n554), .B1(new_n542), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n623), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n667), .B1(new_n670), .B2(KEYINPUT93), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(KEYINPUT93), .B2(new_n667), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n628), .A2(new_n666), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n625), .A2(new_n666), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n613), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n675), .B1(new_n628), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n624), .A2(new_n666), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n628), .B2(new_n666), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n680), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n227), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G1), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n571), .A2(new_n530), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n688), .A2(new_n689), .B1(new_n231), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n566), .A2(new_n519), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n608), .A3(new_n620), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n506), .A2(new_n511), .B1(new_n608), .B2(new_n483), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n337), .A3(new_n552), .A4(new_n566), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(new_n666), .ZN(new_n700));
  XNOR2_X1  g0500(.A(KEYINPUT94), .B(KEYINPUT31), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n517), .A2(new_n523), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT86), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n640), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n614), .B1(new_n629), .B2(KEYINPUT86), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n705), .A2(new_n554), .A3(new_n706), .A4(new_n668), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n702), .B(new_n707), .C1(KEYINPUT31), .C2(new_n700), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n642), .A2(new_n668), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT95), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n642), .A2(KEYINPUT95), .A3(new_n668), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT29), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n641), .A2(new_n584), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n635), .A2(KEYINPUT26), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n636), .A2(new_n638), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n666), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n710), .A2(new_n715), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n691), .B1(new_n723), .B2(G1), .ZN(G364));
  AOI21_X1  g0524(.A(new_n688), .B1(G45), .B2(new_n660), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n674), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G330), .B2(new_n672), .ZN(new_n727));
  INV_X1    g0527(.A(new_n725), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n221), .A2(new_n337), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n330), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n330), .A2(G179), .A3(G200), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(new_n221), .ZN(new_n733));
  AOI22_X1  g0533(.A1(G326), .A2(new_n731), .B1(new_n733), .B2(G294), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n730), .A2(G190), .ZN(new_n735));
  INV_X1    g0535(.A(G317), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT33), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(KEYINPUT33), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n221), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n330), .A3(G200), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT97), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n729), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT97), .B1(new_n221), .B2(new_n337), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G190), .A2(G200), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G311), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n280), .B1(new_n741), .B2(new_n743), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n742), .A2(new_n747), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n740), .B(new_n751), .C1(G329), .C2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(G322), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n745), .A2(G190), .A3(new_n295), .A4(new_n746), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n754), .B1(new_n547), .B2(new_n755), .C1(new_n756), .C2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT99), .Z(new_n763));
  INV_X1    g0563(.A(G159), .ZN(new_n764));
  OR3_X1    g0564(.A1(new_n752), .A2(KEYINPUT32), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n733), .A2(G97), .ZN(new_n766));
  INV_X1    g0566(.A(new_n755), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G87), .ZN(new_n768));
  OAI21_X1  g0568(.A(KEYINPUT32), .B1(new_n752), .B2(new_n764), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n765), .A2(new_n766), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n731), .ZN(new_n771));
  INV_X1    g0571(.A(new_n735), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n276), .B1(new_n771), .B2(new_n202), .C1(new_n213), .C2(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n770), .B(new_n773), .C1(G77), .C2(new_n748), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n774), .B1(new_n254), .B2(new_n761), .C1(new_n492), .C2(new_n743), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n763), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n233), .B1(G20), .B2(new_n339), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n728), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n777), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n249), .A2(new_n308), .B1(new_n232), .B2(new_n316), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n685), .A2(new_n270), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n227), .A2(new_n276), .ZN(new_n788));
  XOR2_X1   g0588(.A(G355), .B(KEYINPUT96), .Z(new_n789));
  OAI22_X1  g0589(.A1(new_n785), .A2(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n530), .B2(new_n685), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n778), .B1(new_n672), .B2(new_n782), .C1(new_n784), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n727), .A2(new_n792), .ZN(G396));
  AOI22_X1  g0593(.A1(new_n748), .A2(G159), .B1(G150), .B2(new_n735), .ZN(new_n794));
  INV_X1    g0594(.A(G137), .ZN(new_n795));
  INV_X1    g0595(.A(G143), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n794), .B1(new_n795), .B2(new_n771), .C1(new_n761), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT34), .ZN(new_n798));
  INV_X1    g0598(.A(new_n733), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n799), .A2(new_n254), .B1(new_n743), .B2(new_n213), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n477), .B(new_n800), .C1(G132), .C2(new_n753), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n798), .B(new_n801), .C1(new_n202), .C2(new_n755), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n743), .A2(new_n208), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n748), .A2(G116), .B1(G283), .B2(new_n735), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT100), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n766), .B(new_n280), .C1(new_n750), .C2(new_n752), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n771), .A2(new_n547), .B1(new_n492), .B2(new_n755), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n805), .B(new_n808), .C1(new_n761), .C2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n802), .B1(new_n803), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n777), .A2(new_n779), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n811), .A2(new_n777), .B1(new_n206), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n408), .B1(new_n407), .B2(new_n668), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n397), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n397), .A2(new_n666), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n779), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n813), .A2(new_n725), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n713), .A2(new_n714), .A3(new_n818), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n666), .B1(new_n716), .B2(new_n639), .ZN(new_n822));
  INV_X1    g0622(.A(new_n818), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n728), .B1(new_n825), .B2(new_n709), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT101), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n709), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n820), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT102), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(G384));
  NOR2_X1   g0634(.A1(new_n463), .A2(new_n666), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT38), .ZN(new_n836));
  INV_X1    g0636(.A(new_n664), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n346), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n654), .B2(new_n335), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n334), .A2(KEYINPUT92), .A3(new_n838), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT37), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n345), .A2(new_n346), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n334), .A2(new_n842), .A3(new_n838), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n334), .A2(new_n838), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n845), .A2(new_n649), .A3(KEYINPUT37), .A4(new_n842), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n836), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT39), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n272), .A2(new_n274), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT7), .B1(new_n270), .B2(G20), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n266), .A2(new_n267), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n852), .A3(G68), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT16), .B1(new_n853), .B2(new_n260), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n293), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n837), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n650), .A2(new_n651), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n645), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n294), .A2(new_n333), .B1(new_n345), .B2(new_n855), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n857), .B1(new_n861), .B2(KEYINPUT103), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT103), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n346), .B1(new_n332), .B2(new_n324), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n260), .B1(new_n268), .B2(new_n271), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n275), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n274), .A3(new_n272), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n293), .A2(new_n867), .B1(new_n343), .B2(new_n344), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n863), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n860), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  AND4_X1   g0670(.A1(new_n860), .A2(new_n334), .A3(new_n842), .A4(new_n838), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n859), .B(KEYINPUT38), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n848), .A2(new_n849), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n345), .A2(new_n855), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n334), .A2(new_n874), .A3(KEYINPUT103), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n869), .A2(new_n875), .A3(new_n856), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n871), .B1(new_n876), .B2(KEYINPUT37), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n856), .B1(new_n335), .B2(new_n348), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n836), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n849), .B1(new_n879), .B2(new_n872), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n873), .A2(KEYINPUT104), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT104), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n872), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n848), .A2(new_n849), .A3(new_n872), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n835), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n654), .A2(new_n837), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n816), .B1(new_n822), .B2(new_n823), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n462), .B(new_n666), .C1(new_n454), .C2(new_n461), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n462), .A2(new_n666), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n463), .A2(new_n450), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n883), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n887), .A2(new_n889), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n468), .B1(new_n715), .B2(new_n722), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n899), .A2(new_n657), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n898), .B(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  INV_X1    g0702(.A(new_n883), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n818), .B1(new_n891), .B2(new_n893), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n699), .A2(new_n666), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n707), .A2(new_n905), .A3(new_n701), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(KEYINPUT31), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n904), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n902), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n700), .B1(new_n631), .B2(new_n668), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n907), .B1(new_n911), .B2(new_n701), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n848), .A2(new_n872), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n913), .A4(new_n904), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n468), .A2(new_n912), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n915), .B(new_n916), .Z(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(G330), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n901), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n220), .B2(new_n660), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n498), .A2(new_n499), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT35), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n221), .B(new_n233), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(G116), .C1(new_n922), .C2(new_n921), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT36), .ZN(new_n925));
  OAI21_X1  g0725(.A(G77), .B1(new_n254), .B2(new_n213), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n926), .A2(new_n231), .B1(G50), .B2(new_n213), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(G1), .A3(new_n659), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n920), .A2(new_n925), .A3(new_n928), .ZN(G367));
  OAI22_X1  g0729(.A1(new_n772), .A2(new_n809), .B1(new_n217), .B2(new_n743), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(G311), .B2(new_n731), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n492), .B2(new_n799), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n767), .A2(KEYINPUT46), .A3(G116), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n749), .B2(new_n741), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT46), .B1(new_n767), .B2(G116), .ZN(new_n935));
  NOR4_X1   g0735(.A1(new_n932), .A2(new_n270), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n936), .B1(new_n547), .B2(new_n761), .C1(new_n736), .C2(new_n752), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n733), .A2(G68), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n254), .B2(new_n755), .C1(new_n771), .C2(new_n796), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n749), .A2(new_n202), .B1(new_n206), .B2(new_n743), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n276), .B1(new_n752), .B2(new_n795), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n942), .B1(new_n764), .B2(new_n772), .C1(new_n761), .C2(new_n362), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT110), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT47), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n728), .B1(new_n946), .B2(new_n777), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n783), .B1(new_n227), .B2(new_n576), .C1(new_n787), .C2(new_n244), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n579), .A2(new_n668), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n581), .A2(new_n584), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT105), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n584), .A2(new_n949), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n950), .A2(new_n951), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n947), .B(new_n948), .C1(new_n782), .C2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n220), .B1(new_n660), .B2(G45), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n513), .A2(new_n668), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n502), .A2(new_n666), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n959), .B1(new_n629), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n683), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT44), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n962), .B(new_n964), .Z(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n963), .B2(KEYINPUT44), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n683), .A2(new_n961), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n680), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n966), .A2(new_n679), .A3(new_n969), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n678), .B(new_n681), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n673), .B(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n723), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n723), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n686), .B(KEYINPUT41), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n958), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n682), .A2(new_n703), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT42), .Z(new_n982));
  INV_X1    g0782(.A(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT106), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n983), .A2(KEYINPUT106), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n955), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n961), .A2(new_n628), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n666), .B1(new_n987), .B2(new_n517), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n982), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n986), .B1(new_n982), .B2(new_n988), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n679), .A2(new_n961), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n992), .B1(KEYINPUT107), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT107), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n994), .B(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n956), .B1(new_n980), .B2(new_n996), .ZN(G387));
  OR2_X1    g0797(.A1(new_n723), .A2(new_n976), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(new_n686), .A3(new_n977), .ZN(new_n999));
  INV_X1    g0799(.A(new_n777), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n748), .A2(G303), .B1(G311), .B2(new_n735), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n756), .B2(new_n771), .C1(new_n761), .C2(new_n736), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT48), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n741), .B2(new_n799), .C1(new_n809), .C2(new_n755), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT49), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n753), .A2(G326), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n743), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n270), .B1(G116), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n270), .B1(new_n217), .B2(new_n743), .C1(new_n362), .C2(new_n752), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n799), .A2(new_n576), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n206), .B2(new_n755), .C1(new_n764), .C2(new_n771), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1012), .B(new_n1015), .C1(G68), .C2(new_n748), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n202), .B2(new_n761), .C1(new_n291), .C2(new_n772), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1000), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n678), .A2(new_n782), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n316), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n786), .B1(new_n241), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n227), .A2(new_n276), .A3(new_n689), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n213), .A2(new_n206), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n292), .A2(new_n202), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n689), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n308), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1023), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n685), .A2(new_n492), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n784), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OR3_X1    g0831(.A1(new_n1018), .A2(new_n1019), .A3(new_n1031), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n999), .B1(new_n728), .B2(new_n1032), .C1(new_n957), .C2(new_n975), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT112), .ZN(G393));
  AOI22_X1  g0834(.A1(new_n760), .A2(G311), .B1(G317), .B2(new_n731), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT52), .Z(new_n1036));
  OAI22_X1  g0836(.A1(new_n749), .A2(new_n809), .B1(new_n492), .B2(new_n743), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n799), .A2(new_n530), .B1(new_n755), .B2(new_n741), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n280), .B1(new_n752), .B2(new_n756), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1036), .B(new_n1040), .C1(new_n547), .C2(new_n772), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n760), .A2(G159), .B1(G150), .B2(new_n731), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT51), .Z(new_n1043));
  AOI21_X1  g0843(.A(new_n477), .B1(G143), .B2(new_n753), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n733), .A2(G77), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n213), .C2(new_n755), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n748), .A2(new_n292), .B1(G50), .B2(new_n735), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1046), .B1(KEYINPUT113), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(KEYINPUT113), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(new_n803), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1043), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1041), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n728), .B1(new_n1052), .B2(new_n777), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n783), .B1(new_n217), .B2(new_n227), .C1(new_n787), .C2(new_n252), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n961), .A2(new_n781), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n973), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1057), .B1(new_n1058), .B2(new_n958), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n973), .A2(new_n977), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n686), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n973), .A2(new_n977), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(G390));
  NAND3_X1  g0863(.A1(new_n468), .A2(G330), .A3(new_n912), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n899), .A2(new_n657), .A3(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n823), .A2(G330), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n708), .A2(new_n894), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT114), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n708), .A2(KEYINPUT114), .A3(new_n894), .A4(new_n1066), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n912), .A2(new_n1066), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n895), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n816), .B1(new_n720), .B2(new_n815), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n890), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n912), .A2(new_n894), .A3(new_n1066), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n894), .B1(new_n708), .B2(new_n1066), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1065), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT104), .B1(new_n873), .B2(new_n880), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n884), .A2(new_n882), .A3(new_n885), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n835), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n890), .B2(new_n895), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1085), .B(new_n913), .C1(new_n1074), .C2(new_n895), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1077), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1071), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1091), .A3(new_n1088), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1082), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1087), .A2(new_n1091), .A3(new_n1088), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1078), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1081), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n686), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n958), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1045), .B1(new_n771), .B2(new_n741), .C1(new_n492), .C2(new_n772), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n276), .B(new_n1100), .C1(G97), .C2(new_n748), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n760), .A2(G116), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n743), .A2(new_n213), .B1(new_n752), .B2(new_n809), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT115), .Z(new_n1104));
  NAND4_X1  g0904(.A1(new_n1101), .A2(new_n768), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n276), .B1(new_n799), .B2(new_n764), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n767), .A2(G150), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT53), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT54), .B(G143), .Z(new_n1109));
  AOI211_X1 g0909(.A(new_n1106), .B(new_n1108), .C1(new_n748), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n753), .A2(G125), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n760), .A2(G132), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n772), .A2(new_n795), .B1(new_n771), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G50), .B2(new_n1009), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .A4(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1000), .B1(new_n1105), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n291), .B2(new_n812), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n725), .B(new_n1118), .C1(new_n1119), .C2(new_n780), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1097), .A2(new_n1099), .A3(new_n1120), .ZN(G378));
  NAND3_X1  g0921(.A1(new_n910), .A2(new_n914), .A3(G330), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n369), .A2(new_n837), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT55), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n380), .A2(new_n405), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n380), .B2(new_n405), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n380), .A2(new_n405), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT55), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n380), .A2(new_n405), .A3(new_n1125), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n1123), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1128), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1122), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT119), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1128), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1134), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1136), .A2(KEYINPUT119), .A3(new_n1137), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1145), .A2(G330), .A3(new_n910), .A4(new_n914), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n898), .A2(new_n1139), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1119), .A2(new_n835), .B1(new_n883), .B2(new_n896), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n889), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1150), .A3(new_n958), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n731), .A2(G125), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n767), .A2(new_n1109), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n733), .A2(G150), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G137), .B2(new_n748), .ZN(new_n1156));
  INV_X1    g0956(.A(G132), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n772), .C1(new_n761), .C2(new_n1113), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT116), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(KEYINPUT116), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT59), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT59), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n1163), .A3(new_n1160), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G33), .B1(new_n753), .B2(G124), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G41), .B1(new_n1009), .B2(G159), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n305), .B1(new_n477), .B2(new_n278), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n202), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n735), .A2(G97), .B1(new_n1009), .B2(G58), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n477), .C1(new_n530), .C2(new_n771), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G107), .B2(new_n760), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n938), .B1(new_n206), .B2(new_n755), .C1(new_n741), .C2(new_n752), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n390), .B2(new_n748), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1172), .A2(new_n305), .A3(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT58), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1167), .A2(new_n1169), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n777), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT117), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n777), .A2(G50), .A3(new_n779), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1181), .B(new_n725), .C1(new_n1145), .C2(new_n780), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT120), .Z(new_n1183));
  NAND2_X1  g0983(.A1(new_n1151), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(KEYINPUT121), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT121), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1151), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1065), .B1(new_n1098), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1190), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n898), .B(new_n1148), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1065), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1096), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1197), .A3(KEYINPUT57), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1194), .A2(new_n686), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1189), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(G375));
  NAND3_X1  g1002(.A1(new_n1075), .A2(new_n1080), .A3(new_n1065), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(KEYINPUT122), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1203), .A2(KEYINPUT122), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n979), .B(new_n1082), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1014), .B1(new_n530), .B2(new_n772), .C1(new_n809), .C2(new_n771), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n280), .B1(new_n752), .B2(new_n547), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n749), .A2(new_n492), .B1(new_n206), .B2(new_n743), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n217), .B2(new_n755), .C1(new_n761), .C2(new_n741), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n270), .B1(new_n254), .B2(new_n743), .C1(new_n1113), .C2(new_n752), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n735), .A2(new_n1109), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n799), .B2(new_n202), .C1(new_n1157), .C2(new_n771), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(G150), .C2(new_n748), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n795), .B2(new_n761), .C1(new_n764), .C2(new_n755), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1000), .B1(new_n1212), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n213), .B2(new_n812), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n725), .B(new_n1219), .C1(new_n894), .C2(new_n780), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1191), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1220), .B1(new_n1221), .B2(new_n957), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1207), .A2(new_n1223), .ZN(G381));
  NOR2_X1   g1024(.A1(G375), .A2(G378), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1033), .A2(KEYINPUT112), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1033), .A2(KEYINPUT112), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n792), .A3(new_n727), .A4(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1228), .A2(G384), .A3(G390), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G387), .A2(G381), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1225), .A2(new_n1229), .A3(new_n1230), .ZN(G407));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1225), .B2(new_n665), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(G407), .ZN(G409));
  INV_X1    g1034(.A(KEYINPUT63), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1188), .A2(new_n1199), .A3(G378), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT123), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1188), .A2(new_n1199), .A3(KEYINPUT123), .A4(G378), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT124), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1147), .A2(new_n1150), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n957), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1182), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1241), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1195), .A2(new_n1197), .A3(new_n979), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n958), .B1(new_n1195), .B2(new_n1242), .ZN(new_n1249));
  OAI211_X1 g1049(.A(KEYINPUT125), .B(new_n1182), .C1(new_n1249), .C2(new_n1243), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(G378), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1240), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(G384), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT60), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1205), .A2(new_n1206), .B1(new_n1256), .B2(new_n1081), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1203), .A2(new_n1256), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1257), .A2(new_n686), .A3(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1255), .B1(new_n1260), .B2(new_n1222), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1257), .B(new_n686), .C1(new_n1256), .C2(new_n1203), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(G384), .A3(new_n1223), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1232), .A2(G343), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1254), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(G2897), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1261), .A2(new_n1263), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1269), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1238), .A2(new_n1239), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1273), .B2(new_n1266), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1235), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G390), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G387), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G390), .B(new_n956), .C1(new_n980), .C2(new_n996), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT126), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1228), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1228), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G387), .A2(new_n1276), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1279), .A2(new_n1284), .B1(KEYINPUT126), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1283), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  AOI211_X1 g1088(.A(new_n1264), .B(new_n1266), .C1(new_n1240), .C2(new_n1253), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(KEYINPUT63), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1275), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1269), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1264), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1261), .A2(new_n1263), .A3(new_n1269), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1254), .B2(new_n1267), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT63), .B1(new_n1297), .B2(new_n1289), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1283), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n1268), .B2(new_n1235), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT127), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT62), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1266), .B1(new_n1240), .B2(new_n1253), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1304), .B2(new_n1265), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1302), .A2(KEYINPUT61), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n1292), .A2(new_n1301), .B1(new_n1306), .B2(new_n1308), .ZN(G405));
  OAI21_X1  g1109(.A(new_n1240), .B1(G378), .B2(new_n1201), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(new_n1265), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(new_n1307), .ZN(G402));
endmodule


