//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT76), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n190), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G137), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G134), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n199), .A2(new_n200), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n200), .B1(new_n199), .B2(new_n206), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT0), .B(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT3), .B1(new_n220), .B2(G107), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n222));
  INV_X1    g036(.A(G107), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G104), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(G107), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(G101), .A3(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n226), .A2(G101), .ZN(new_n229));
  INV_X1    g043(.A(G101), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n221), .A2(new_n224), .A3(new_n230), .A4(new_n225), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT4), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n219), .B(new_n228), .C1(new_n229), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT1), .B1(new_n212), .B2(G146), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n212), .A2(G146), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n210), .A2(G143), .ZN(new_n236));
  OAI211_X1 g050(.A(G128), .B(new_n234), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G128), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n211), .B(new_n213), .C1(KEYINPUT1), .C2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n223), .A2(G104), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n220), .A2(G107), .ZN(new_n242));
  OAI21_X1  g056(.A(G101), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n231), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n244), .A3(KEYINPUT10), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n237), .A2(new_n231), .A3(new_n243), .A4(new_n239), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT10), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n233), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n209), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n233), .A2(new_n245), .A3(KEYINPUT79), .A4(new_n248), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n251), .A2(KEYINPUT80), .A3(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n233), .A2(new_n245), .A3(new_n209), .A4(new_n248), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT80), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n251), .B2(new_n252), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n194), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT78), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n246), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n240), .B2(new_n244), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n239), .A2(new_n237), .B1(new_n231), .B2(new_n243), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n259), .A3(new_n246), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n209), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT12), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n254), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n209), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n262), .B1(new_n259), .B2(new_n246), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n240), .A2(new_n244), .A3(KEYINPUT78), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(KEYINPUT12), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n193), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n258), .A2(G469), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G469), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n249), .A2(new_n250), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n267), .A3(new_n252), .ZN(new_n280));
  INV_X1    g094(.A(new_n256), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n251), .A2(KEYINPUT80), .A3(new_n252), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n193), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n264), .A2(new_n265), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n270), .A2(KEYINPUT12), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n254), .A4(new_n194), .ZN(new_n287));
  AOI211_X1 g101(.A(G469), .B(G902), .C1(new_n284), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n189), .B1(new_n278), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G214), .B1(G237), .B2(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(KEYINPUT2), .A2(G113), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NOR3_X1   g107(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G116), .B(G119), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n300));
  INV_X1    g114(.A(G113), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n292), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n291), .A3(new_n296), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n226), .A2(G101), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT4), .A3(new_n231), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n307), .A3(new_n228), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n296), .A2(KEYINPUT5), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT81), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT5), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(G116), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n309), .A2(new_n310), .A3(G113), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(G116), .ZN(new_n315));
  INV_X1    g129(.A(G116), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G119), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT5), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(G113), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT81), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n244), .A2(new_n314), .A3(new_n320), .A4(new_n304), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n308), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT82), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n308), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  XNOR2_X1  g139(.A(G110), .B(G122), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n323), .A2(new_n325), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n237), .A2(new_n330), .A3(new_n239), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n215), .B(G125), .C1(new_n216), .C2(new_n217), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n191), .A2(G224), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n334), .A2(KEYINPUT84), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(KEYINPUT84), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n333), .B(new_n337), .Z(new_n338));
  AND3_X1   g152(.A1(new_n308), .A2(new_n324), .A3(new_n321), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n324), .B1(new_n308), .B2(new_n321), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n339), .A2(new_n340), .A3(new_n326), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n308), .A2(new_n321), .A3(new_n326), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT6), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n329), .B(new_n338), .C1(new_n341), .C2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G210), .B1(G237), .B2(G902), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n336), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n333), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n326), .B(KEYINPUT8), .Z(new_n348));
  OAI21_X1  g162(.A(new_n304), .B1(new_n318), .B2(new_n319), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(new_n244), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n231), .A2(new_n243), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n314), .A2(new_n320), .A3(new_n304), .A4(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n347), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n333), .A2(new_n346), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n333), .A2(KEYINPUT85), .A3(new_n346), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n353), .A2(new_n342), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(new_n275), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n344), .A2(new_n345), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n345), .B1(new_n344), .B2(new_n359), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n290), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n203), .A2(new_n205), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT91), .B1(new_n238), .B2(G143), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT91), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n212), .A3(G128), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n238), .A2(G143), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n364), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT13), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n365), .A2(new_n367), .A3(KEYINPUT13), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n374), .B2(G134), .ZN(new_n375));
  OR2_X1    g189(.A1(KEYINPUT89), .A2(G122), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT89), .A2(G122), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n316), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n316), .A2(G122), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT90), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n377), .ZN(new_n382));
  NOR2_X1   g196(.A1(KEYINPUT89), .A2(G122), .ZN(new_n383));
  OAI21_X1  g197(.A(G116), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT90), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(new_n379), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n223), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n223), .B1(new_n381), .B2(new_n386), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n375), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n368), .A2(new_n369), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n203), .A2(new_n205), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n364), .A2(new_n368), .A3(new_n369), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n379), .A2(KEYINPUT14), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n379), .A2(KEYINPUT14), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n384), .A3(new_n396), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n393), .A2(new_n394), .B1(new_n397), .B2(G107), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n387), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT70), .B(G217), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n188), .A2(G953), .A3(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n390), .A2(KEYINPUT92), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n381), .A2(new_n386), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G107), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n387), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n405), .A2(new_n375), .B1(new_n398), .B2(new_n387), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n406), .B2(new_n401), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT92), .B1(new_n406), .B2(new_n401), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n275), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT93), .ZN(new_n410));
  INV_X1    g224(.A(G478), .ZN(new_n411));
  NOR2_X1   g225(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n390), .A2(new_n399), .A3(new_n401), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT92), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n390), .A2(new_n399), .ZN(new_n419));
  INV_X1    g233(.A(new_n401), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n421), .A3(new_n402), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT93), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n275), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n410), .A2(new_n415), .A3(new_n424), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n409), .A2(new_n415), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n330), .A2(KEYINPUT16), .A3(G140), .ZN(new_n428));
  XNOR2_X1  g242(.A(G125), .B(G140), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(KEYINPUT16), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G146), .ZN(new_n431));
  AOI211_X1 g245(.A(new_n210), .B(new_n428), .C1(KEYINPUT16), .C2(new_n429), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g247(.A1(KEYINPUT86), .A2(G143), .ZN(new_n434));
  NOR2_X1   g248(.A1(G237), .A2(G953), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(G214), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(KEYINPUT86), .A2(G143), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n434), .A2(new_n438), .B1(new_n435), .B2(G214), .ZN(new_n439));
  OAI211_X1 g253(.A(KEYINPUT17), .B(G131), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G131), .B1(new_n437), .B2(new_n439), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n434), .A2(new_n438), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n435), .A2(G214), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(new_n200), .A3(new_n436), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n433), .B(new_n440), .C1(new_n446), .C2(KEYINPUT17), .ZN(new_n447));
  XNOR2_X1  g261(.A(G113), .B(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(G104), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G140), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G125), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n330), .A2(G140), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(G146), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n210), .B1(new_n452), .B2(new_n453), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT87), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n456), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n429), .A2(new_n210), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT18), .B(G131), .C1(new_n437), .C2(new_n439), .ZN(new_n463));
  NAND2_X1  g277(.A1(KEYINPUT18), .A2(G131), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n444), .A2(new_n464), .A3(new_n436), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT88), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n462), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n465), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n444), .B2(new_n436), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n457), .A2(new_n461), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT88), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n447), .B(new_n450), .C1(new_n468), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n467), .B1(new_n462), .B2(new_n466), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(KEYINPUT88), .A3(new_n472), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n450), .B1(new_n478), .B2(new_n447), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n275), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G475), .ZN(new_n481));
  NAND2_X1  g295(.A1(G234), .A2(G237), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n482), .A2(G952), .A3(new_n191), .ZN(new_n483));
  XOR2_X1   g297(.A(KEYINPUT21), .B(G898), .Z(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT95), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n482), .A2(G902), .A3(G953), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n429), .B(KEYINPUT19), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n432), .B1(new_n490), .B2(new_n210), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n476), .A2(new_n477), .B1(new_n446), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n474), .B1(new_n492), .B2(new_n450), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  NOR2_X1   g308(.A1(G475), .A2(G902), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n481), .B(new_n489), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  NOR4_X1   g313(.A1(new_n289), .A2(new_n363), .A3(new_n427), .A4(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n219), .B1(new_n207), .B2(new_n208), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n303), .A2(new_n291), .A3(new_n296), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n296), .B1(new_n303), .B2(new_n291), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n199), .A2(new_n200), .A3(new_n206), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n200), .B1(G134), .B2(G137), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n392), .B2(G137), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n505), .A2(new_n239), .A3(new_n237), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n501), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT67), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n501), .A2(new_n508), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n514), .B2(new_n305), .ZN(new_n515));
  AOI211_X1 g329(.A(KEYINPUT67), .B(new_n504), .C1(new_n501), .C2(new_n508), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n512), .B1(new_n517), .B2(KEYINPUT28), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n435), .A2(G210), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT27), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT26), .B(G101), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(KEYINPUT66), .A2(KEYINPUT31), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AND4_X1   g338(.A1(new_n505), .A2(new_n239), .A3(new_n237), .A4(new_n507), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n196), .A2(new_n198), .ZN(new_n527));
  OAI21_X1  g341(.A(G131), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n218), .B1(new_n528), .B2(new_n505), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n525), .A2(new_n529), .A3(new_n305), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT30), .B1(new_n525), .B2(new_n529), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n501), .A2(new_n532), .A3(new_n508), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n530), .B1(new_n534), .B2(new_n305), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT66), .A2(KEYINPUT31), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n522), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n524), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n504), .B1(new_n531), .B2(new_n533), .ZN(new_n540));
  NOR4_X1   g354(.A1(new_n540), .A2(new_n530), .A3(new_n523), .A4(new_n537), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n518), .A2(new_n522), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(G472), .A2(G902), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(KEYINPUT32), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n305), .B1(new_n525), .B2(new_n529), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT67), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n514), .A2(new_n513), .A3(new_n305), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n530), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n511), .B1(new_n550), .B2(new_n510), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n522), .ZN(new_n552));
  INV_X1    g366(.A(new_n522), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n535), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT29), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n504), .B1(new_n501), .B2(new_n508), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT28), .B1(new_n530), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n557), .A2(KEYINPUT29), .A3(new_n511), .A4(new_n522), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n275), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT68), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n561), .A3(new_n275), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G472), .B1(new_n555), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n542), .A2(new_n543), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT32), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n542), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n543), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n546), .A2(new_n564), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT72), .B1(new_n312), .B2(G128), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT23), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT23), .ZN(new_n572));
  OAI211_X1 g386(.A(KEYINPUT72), .B(new_n572), .C1(new_n312), .C2(G128), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n312), .A2(G128), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G110), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(KEYINPUT71), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT71), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n312), .A3(G128), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n577), .A2(new_n579), .B1(G119), .B2(new_n238), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT24), .B(G110), .Z(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n576), .B(new_n582), .C1(new_n431), .C2(new_n432), .ZN(new_n583));
  OAI22_X1  g397(.A1(new_n575), .A2(G110), .B1(new_n580), .B2(new_n581), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n455), .B1(new_n430), .B2(G146), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT22), .B(G137), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n583), .A2(new_n586), .A3(new_n590), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n275), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n592), .A2(KEYINPUT25), .A3(new_n275), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n400), .B1(G234), .B2(new_n275), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n593), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n590), .B1(new_n583), .B2(new_n586), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n599), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n275), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT73), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n600), .A2(new_n607), .A3(KEYINPUT74), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT74), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n604), .B1(new_n596), .B2(new_n597), .ZN(new_n610));
  INV_X1    g424(.A(new_n607), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n569), .A2(KEYINPUT75), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT75), .B1(new_n569), .B2(new_n614), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n500), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  NAND3_X1  g432(.A1(new_n410), .A2(new_n411), .A3(new_n424), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT96), .B(KEYINPUT33), .Z(new_n620));
  NAND2_X1  g434(.A1(new_n422), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n421), .A2(KEYINPUT33), .A3(new_n416), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(G478), .A3(new_n275), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n481), .B1(new_n497), .B2(new_n498), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n489), .B(new_n290), .C1(new_n361), .C2(new_n362), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT97), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n627), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n493), .A2(new_n495), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n496), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n619), .A2(new_n623), .B1(new_n632), .B2(new_n481), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n629), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n628), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n542), .B2(new_n275), .ZN(new_n638));
  INV_X1    g452(.A(new_n543), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n534), .A2(new_n305), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n509), .A3(new_n538), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n523), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n535), .A2(new_n524), .A3(new_n538), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n551), .A2(new_n553), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n613), .A2(new_n638), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n289), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n636), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  AND2_X1   g466(.A1(new_n425), .A2(new_n426), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT98), .B1(new_n653), .B2(new_n499), .ZN(new_n654));
  INV_X1    g468(.A(new_n290), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n344), .A2(new_n359), .ZN(new_n656));
  INV_X1    g470(.A(new_n345), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n655), .B1(new_n658), .B2(new_n360), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n631), .A2(new_n496), .B1(G475), .B2(new_n480), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n427), .A2(new_n660), .A3(new_n489), .A4(new_n661), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n654), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n649), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n587), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n606), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n600), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n290), .C1(new_n361), .C2(new_n362), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n289), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n427), .A2(new_n499), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n638), .A2(new_n646), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(new_n483), .ZN(new_n678));
  INV_X1    g492(.A(new_n487), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n678), .B1(new_n679), .B2(G900), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n427), .A2(new_n661), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n569), .A2(new_n672), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  INV_X1    g497(.A(new_n535), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n522), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n530), .A2(new_n556), .ZN(new_n686));
  AOI21_X1  g500(.A(G902), .B1(new_n686), .B2(new_n553), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n637), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n565), .B2(new_n566), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n546), .A3(new_n568), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n361), .A2(new_n362), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT38), .ZN(new_n693));
  INV_X1    g507(.A(new_n670), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n427), .A2(new_n625), .A3(new_n290), .A4(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n680), .B(KEYINPUT39), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n648), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  AND3_X1   g516(.A1(new_n624), .A2(new_n625), .A3(new_n680), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n569), .A2(new_n672), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  AOI21_X1  g519(.A(G902), .B1(new_n284), .B2(new_n287), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n274), .ZN(new_n707));
  INV_X1    g521(.A(new_n189), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n707), .A2(new_n288), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n569), .A2(new_n614), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n636), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT41), .B(G113), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT99), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n711), .B(new_n713), .ZN(G15));
  NAND3_X1  g528(.A1(new_n569), .A2(new_n614), .A3(new_n709), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n654), .A2(new_n659), .A3(new_n662), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n316), .ZN(G18));
  NOR4_X1   g532(.A1(new_n363), .A2(new_n707), .A3(new_n288), .A4(new_n708), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n427), .A2(new_n499), .A3(new_n694), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n569), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  XNOR2_X1  g536(.A(new_n543), .B(KEYINPUT100), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n557), .A2(new_n511), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n553), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n723), .B1(new_n644), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n600), .A2(new_n607), .ZN(new_n727));
  NOR4_X1   g541(.A1(new_n638), .A2(new_n726), .A3(new_n727), .A4(new_n488), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n427), .A2(new_n659), .A3(new_n625), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n709), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NOR3_X1   g545(.A1(new_n638), .A2(new_n694), .A3(new_n726), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n719), .A2(new_n703), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  NOR2_X1   g548(.A1(new_n708), .A2(new_n655), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n658), .A2(new_n360), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n272), .A2(KEYINPUT101), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n272), .A2(KEYINPUT101), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(G469), .A3(new_n258), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n276), .B1(new_n706), .B2(new_n274), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n569), .A2(new_n614), .A3(new_n703), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n703), .A2(new_n741), .A3(KEYINPUT42), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n554), .B1(new_n518), .B2(new_n553), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n558), .A2(new_n561), .A3(new_n275), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n561), .B1(new_n558), .B2(new_n275), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n637), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g566(.A(new_n566), .B(new_n639), .C1(new_n644), .C2(new_n645), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT32), .B1(new_n542), .B2(new_n543), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT102), .B1(new_n755), .B2(new_n727), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n564), .A2(new_n567), .A3(new_n544), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT102), .ZN(new_n758));
  INV_X1    g572(.A(new_n727), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n745), .B1(new_n756), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n744), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n200), .ZN(G33));
  NAND4_X1  g577(.A1(new_n569), .A2(new_n614), .A3(new_n681), .A4(new_n741), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND3_X1  g579(.A1(new_n658), .A2(new_n290), .A3(new_n360), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  AOI211_X1 g581(.A(KEYINPUT43), .B(new_n625), .C1(new_n619), .C2(new_n623), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n625), .B(KEYINPUT104), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n624), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n768), .B1(new_n770), .B2(KEYINPUT43), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n771), .B(new_n670), .C1(new_n646), .C2(new_n638), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n767), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT105), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n737), .A2(KEYINPUT45), .A3(new_n258), .A4(new_n738), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT103), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n258), .A2(new_n272), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT45), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n778), .A2(G469), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n782), .B2(new_n277), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n288), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n277), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n708), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n772), .A2(new_n773), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n775), .A2(new_n697), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  AND2_X1   g603(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n569), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n613), .A3(new_n703), .A4(new_n767), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT106), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  NAND3_X1  g611(.A1(new_n693), .A2(new_n759), .A3(new_n735), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n770), .ZN(new_n799));
  OR3_X1    g613(.A1(new_n707), .A2(new_n288), .A3(KEYINPUT49), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT49), .B1(new_n707), .B2(new_n288), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n799), .A2(new_n691), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT107), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n710), .B1(new_n663), .B2(new_n636), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n721), .A2(new_n675), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n427), .A2(new_n661), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n626), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n647), .A3(new_n648), .A4(new_n629), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(new_n730), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n617), .A2(new_n805), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n632), .A2(new_n670), .A3(new_n481), .A4(new_n680), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n427), .A3(new_n766), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n569), .A3(new_n648), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n703), .A2(new_n741), .A3(new_n732), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n764), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n744), .B2(new_n761), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n804), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n628), .A2(new_n635), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n715), .B1(new_n819), .B2(new_n716), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n809), .A2(new_n721), .A3(new_n675), .A4(new_n730), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n764), .A2(new_n814), .A3(new_n815), .ZN(new_n823));
  INV_X1    g637(.A(new_n745), .ZN(new_n824));
  INV_X1    g638(.A(new_n760), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n758), .B1(new_n757), .B2(new_n759), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n742), .A2(new_n743), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n822), .A2(new_n829), .A3(KEYINPUT107), .A4(new_n617), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n818), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n740), .A2(new_n739), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n694), .A2(new_n189), .A3(new_n680), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n690), .A2(new_n729), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n682), .A3(new_n704), .A4(new_n733), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n682), .A2(new_n733), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT108), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n834), .A2(new_n704), .A3(KEYINPUT52), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT108), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n682), .A2(new_n733), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT109), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT109), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n839), .A2(new_n840), .A3(new_n845), .A4(new_n842), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n837), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n803), .B1(new_n831), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT110), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(KEYINPUT110), .B(new_n803), .C1(new_n831), .C2(new_n847), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n822), .A2(new_n829), .A3(new_n617), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n835), .B(KEYINPUT52), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT53), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT54), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n803), .B1(new_n852), .B2(new_n853), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n811), .A2(new_n817), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT53), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n858), .B(new_n859), .C1(new_n847), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT111), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n857), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(new_n857), .B2(new_n863), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n638), .A2(new_n726), .A3(new_n727), .A4(new_n678), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n771), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n707), .A2(new_n288), .A3(new_n189), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n767), .B(new_n868), .C1(new_n792), .C2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n868), .A2(new_n655), .A3(new_n693), .A4(new_n709), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT50), .Z(new_n872));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n709), .A2(new_n483), .A3(new_n767), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n691), .A3(new_n614), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n875), .A2(new_n625), .A3(new_n624), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n771), .A2(new_n732), .A3(new_n874), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n873), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(KEYINPUT114), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n870), .A2(new_n872), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n868), .A2(new_n719), .ZN(new_n887));
  INV_X1    g701(.A(G952), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(G953), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n887), .B(new_n889), .C1(new_n626), .C2(new_n875), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n825), .A2(new_n826), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n892), .A2(new_n771), .A3(new_n874), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT48), .ZN(new_n895));
  XNOR2_X1  g709(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n896));
  AOI211_X1 g710(.A(new_n890), .B(new_n895), .C1(new_n893), .C2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n870), .A2(new_n882), .A3(new_n872), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n886), .B(new_n897), .C1(new_n898), .C2(KEYINPUT51), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n865), .A2(new_n866), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(G952), .A2(G953), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n802), .B1(new_n900), .B2(new_n901), .ZN(G75));
  OR2_X1    g716(.A1(new_n847), .A2(new_n861), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(new_n858), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n275), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n905), .B2(G210), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n329), .B1(new_n341), .B2(new_n343), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n338), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n906), .A2(new_n909), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n191), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n910), .A2(KEYINPUT116), .A3(new_n911), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(G51));
  AND2_X1   g732(.A1(new_n284), .A2(new_n287), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n904), .B2(new_n859), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n862), .B(KEYINPUT117), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n903), .A2(new_n858), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n276), .B(KEYINPUT57), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n919), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n904), .A2(new_n275), .A3(new_n782), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n927), .B2(new_n928), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n912), .B1(new_n929), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  INV_X1    g747(.A(new_n493), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n933), .A2(KEYINPUT120), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n913), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT120), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(G60));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  AND2_X1   g754(.A1(new_n851), .A2(new_n855), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n848), .A2(new_n849), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n859), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT111), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n862), .B(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT112), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n857), .A2(new_n863), .A3(new_n864), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n621), .A2(new_n622), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT121), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT122), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n940), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n865), .B2(new_n866), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT122), .ZN(new_n954));
  INV_X1    g768(.A(new_n950), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n940), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n912), .B1(new_n925), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n951), .A2(new_n956), .A3(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n904), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n603), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(new_n912), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT61), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n962), .A2(new_n668), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(G66));
  INV_X1    g783(.A(G224), .ZN(new_n970));
  OAI21_X1  g784(.A(G953), .B1(new_n486), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n811), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(G953), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n907), .B1(G898), .B2(new_n191), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT124), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n973), .B(new_n975), .ZN(G69));
  NOR2_X1   g790(.A1(new_n191), .A2(G900), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT126), .ZN(new_n978));
  INV_X1    g792(.A(new_n762), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n786), .A2(new_n697), .A3(new_n729), .A4(new_n892), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n839), .A2(new_n704), .A3(new_n842), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n979), .A2(new_n980), .A3(new_n764), .A4(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n788), .A2(new_n796), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n978), .B1(new_n983), .B2(new_n191), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n534), .B(new_n490), .Z(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(G227), .A2(G900), .ZN(new_n987));
  OAI22_X1  g801(.A1(new_n986), .A2(KEYINPUT125), .B1(new_n191), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n981), .A2(new_n701), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT62), .Z(new_n990));
  INV_X1    g804(.A(new_n698), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n766), .B1(new_n626), .B2(new_n807), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n991), .B(new_n992), .C1(new_n615), .C2(new_n616), .ZN(new_n993));
  AND4_X1   g807(.A1(new_n788), .A2(new_n990), .A3(new_n796), .A4(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n985), .B1(new_n994), .B2(G953), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n985), .B2(new_n984), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n988), .B(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n994), .B2(new_n972), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n983), .A2(new_n811), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1002), .A2(new_n1000), .ZN(new_n1003));
  OAI221_X1 g817(.A(new_n913), .B1(new_n1001), .B2(new_n685), .C1(new_n1003), .C2(new_n554), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n685), .A2(new_n554), .A3(new_n999), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n941), .B2(new_n942), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1006), .A2(KEYINPUT127), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(KEYINPUT127), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(G57));
endmodule


