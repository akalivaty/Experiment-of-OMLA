//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G101), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT81), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(KEYINPUT81), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(new_n194), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n191), .A2(G107), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT81), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT3), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n201), .A3(new_n192), .A4(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT66), .A3(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n215), .A3(G143), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n212), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT1), .B1(new_n210), .B2(G146), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n212), .A2(new_n216), .B1(G128), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n196), .B(new_n206), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT82), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT10), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n222), .B2(new_n224), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n203), .A2(KEYINPUT3), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n204), .B1(new_n202), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n192), .B1(new_n194), .B2(new_n198), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT64), .B1(new_n210), .B2(G146), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n208), .A3(G143), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT65), .B(G146), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n233), .B(new_n235), .C1(new_n236), .C2(G143), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n236), .A2(G143), .B1(new_n209), .B2(new_n211), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n237), .A2(new_n240), .B1(new_n241), .B2(new_n238), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(G101), .C1(new_n229), .C2(new_n230), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n232), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT83), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n206), .A2(new_n246), .A3(new_n196), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n246), .B1(new_n206), .B2(new_n196), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n212), .A2(new_n216), .A3(new_n218), .ZN(new_n250));
  AOI21_X1  g064(.A(G143), .B1(new_n213), .B2(new_n215), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n233), .A2(new_n235), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n217), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT10), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n245), .B1(new_n249), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G137), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(G137), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT11), .A3(G134), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G131), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n260), .A2(new_n263), .A3(new_n266), .A4(new_n261), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n227), .A2(new_n257), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n206), .A2(new_n196), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n222), .B1(new_n255), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT12), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n274), .A3(new_n268), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n190), .B1(new_n269), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n268), .B1(new_n227), .B2(new_n257), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n232), .A2(new_n244), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n206), .A2(new_n196), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT83), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n206), .A2(new_n246), .A3(new_n196), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n236), .B2(G143), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n237), .B1(new_n286), .B2(new_n217), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n224), .B1(new_n287), .B2(new_n250), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n242), .A2(new_n280), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n222), .A2(new_n224), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT82), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n268), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n289), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n190), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n279), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n277), .A2(new_n278), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n278), .B1(new_n277), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g113(.A(G469), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G469), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n295), .A2(new_n296), .A3(new_n273), .A4(new_n275), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n296), .B1(new_n279), .B2(new_n295), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(KEYINPUT85), .B(new_n296), .C1(new_n279), .C2(new_n295), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n301), .B(new_n302), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(G469), .A2(G902), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n300), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT86), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT86), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G217), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(G234), .B2(new_n302), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT78), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT22), .B(G137), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  AOI21_X1  g143(.A(G146), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n329), .A3(G146), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(KEYINPUT75), .A3(new_n332), .ZN(new_n333));
  AOI211_X1 g147(.A(KEYINPUT75), .B(G146), .C1(new_n328), .C2(new_n329), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G119), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(G128), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(KEYINPUT74), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n217), .A2(KEYINPUT74), .A3(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(G128), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT24), .B(G110), .Z(new_n343));
  NAND3_X1  g157(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n340), .B(new_n344), .C1(new_n337), .C2(KEYINPUT23), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n342), .A2(new_n343), .B1(new_n345), .B2(G110), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n333), .A2(new_n335), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT76), .B(G110), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n342), .A2(new_n343), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G125), .B(G140), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n236), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT77), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n236), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n349), .A2(new_n355), .A3(new_n332), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n323), .B1(new_n357), .B2(KEYINPUT79), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n347), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n347), .A2(new_n359), .A3(new_n356), .A4(new_n323), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT25), .B1(new_n363), .B2(new_n302), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n365), .B(G902), .C1(new_n361), .C2(new_n362), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n319), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n319), .A2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT80), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n367), .A2(new_n372), .A3(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT26), .B(G101), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT70), .ZN(new_n376));
  NOR2_X1   g190(.A1(G237), .A2(G953), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(G210), .A3(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n375), .A2(KEYINPUT70), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(G210), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n375), .A2(KEYINPUT70), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n378), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n383), .B1(new_n378), .B2(new_n382), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT2), .A2(G113), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT2), .ZN(new_n389));
  INV_X1    g203(.A(G113), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT67), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT67), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(KEYINPUT2), .B2(G113), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n388), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n336), .A2(G116), .ZN(new_n395));
  INV_X1    g209(.A(G116), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G119), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT68), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n391), .A2(new_n393), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n387), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(new_n397), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(KEYINPUT68), .A3(new_n402), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n261), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n259), .A2(G137), .ZN(new_n408));
  OAI21_X1  g222(.A(G131), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n267), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n287), .B2(new_n250), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n241), .A2(new_n238), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n240), .B1(new_n251), .B2(new_n252), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n268), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT30), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n242), .A2(new_n268), .ZN(new_n416));
  INV_X1    g230(.A(new_n410), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n255), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n406), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n416), .A2(new_n418), .A3(new_n406), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n386), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n268), .A2(new_n242), .B1(new_n255), .B2(new_n417), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT28), .B1(new_n427), .B2(new_n406), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n406), .B1(new_n416), .B2(new_n418), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT71), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n394), .A2(new_n398), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n399), .B(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n411), .B2(new_n414), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT71), .A3(new_n422), .ZN(new_n436));
  AOI211_X1 g250(.A(new_n386), .B(new_n428), .C1(new_n432), .C2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT72), .B1(new_n426), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n428), .B1(new_n432), .B2(new_n436), .ZN(new_n439));
  INV_X1    g253(.A(new_n386), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n441), .A2(new_n442), .A3(new_n425), .A4(new_n424), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n435), .A2(new_n422), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n428), .B1(new_n444), .B2(KEYINPUT28), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n386), .A2(new_n425), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n438), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G472), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT73), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT73), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n451), .A3(G472), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n415), .A2(new_n420), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n423), .B1(new_n454), .B2(new_n434), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT31), .B1(new_n455), .B2(new_n440), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT31), .ZN(new_n457));
  NOR4_X1   g271(.A1(new_n421), .A2(new_n457), .A3(new_n386), .A4(new_n423), .ZN(new_n458));
  OAI22_X1  g272(.A1(new_n456), .A2(new_n458), .B1(new_n440), .B2(new_n439), .ZN(new_n459));
  INV_X1    g273(.A(G472), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n302), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT32), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n459), .A2(new_n463), .A3(new_n460), .A4(new_n302), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n374), .B1(new_n453), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G210), .B1(G237), .B2(G902), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n469), .B(KEYINPUT91), .Z(new_n470));
  XOR2_X1   g284(.A(G110), .B(G122), .Z(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT87), .A2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(KEYINPUT87), .A2(KEYINPUT5), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n395), .B(new_n397), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  OR2_X1    g289(.A1(KEYINPUT87), .A2(KEYINPUT5), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n476), .A2(G116), .A3(new_n336), .A4(new_n472), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n477), .A3(G113), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT88), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n394), .A2(new_n398), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n475), .A2(new_n477), .A3(new_n481), .A4(G113), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n282), .B2(new_n283), .ZN(new_n484));
  AND4_X1   g298(.A1(new_n405), .A2(new_n232), .A3(new_n404), .A4(new_n244), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n471), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n232), .A2(new_n404), .A3(new_n405), .A4(new_n244), .ZN(new_n487));
  INV_X1    g301(.A(new_n471), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n487), .B(new_n488), .C1(new_n249), .C2(new_n483), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(KEYINPUT6), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n491), .B(new_n471), .C1(new_n484), .C2(new_n485), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n412), .A2(new_n413), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G125), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(G125), .B2(new_n255), .ZN(new_n495));
  INV_X1    g309(.A(G224), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G953), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n495), .B(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT89), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n490), .A2(KEYINPUT89), .A3(new_n492), .A4(new_n498), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT7), .B1(new_n496), .B2(G953), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n495), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n503), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n494), .B(new_n505), .C1(G125), .C2(new_n255), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT5), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n477), .B(G113), .C1(new_n507), .C2(new_n402), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n480), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n270), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n471), .B(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n512), .C1(new_n270), .C2(new_n483), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n504), .A2(new_n506), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(G902), .B1(new_n514), .B2(new_n489), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n502), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n470), .B1(new_n501), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n499), .A2(new_n500), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n518), .A2(new_n469), .A3(new_n502), .A4(new_n515), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n468), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G237), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n188), .A3(G214), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n210), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n377), .A2(G143), .A3(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT18), .A2(G131), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n524), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(KEYINPUT18), .A3(G131), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n352), .A2(new_n354), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n350), .A2(new_n208), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n526), .B(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G113), .B(G122), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(new_n191), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(KEYINPUT17), .A3(G131), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(new_n330), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n534), .B1(new_n536), .B2(new_n334), .ZN(new_n537));
  AND4_X1   g351(.A1(G143), .A2(new_n521), .A3(new_n188), .A4(G214), .ZN(new_n538));
  AOI21_X1  g352(.A(G143), .B1(new_n377), .B2(G214), .ZN(new_n539));
  OAI21_X1  g353(.A(G131), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n523), .A2(new_n266), .A3(new_n524), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT93), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n540), .A2(new_n542), .A3(KEYINPUT93), .A4(new_n541), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n531), .B(new_n533), .C1(new_n537), .C2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n333), .A2(new_n335), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n550), .A2(new_n534), .A3(new_n545), .A4(new_n546), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n533), .B1(new_n551), .B2(new_n531), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n302), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G475), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT94), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT19), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n350), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n236), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n332), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n540), .A2(new_n542), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n528), .A2(new_n526), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n530), .B1(new_n352), .B2(new_n354), .ZN(new_n563));
  OAI22_X1  g377(.A1(new_n560), .A2(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n533), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n548), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(G475), .A2(G902), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n556), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  AOI211_X1 g384(.A(KEYINPUT20), .B(new_n570), .C1(new_n548), .C2(new_n566), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n554), .B(new_n555), .C1(new_n569), .C2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n531), .B1(new_n537), .B2(new_n547), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n565), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n574), .B2(new_n548), .ZN(new_n575));
  INV_X1    g389(.A(G475), .ZN(new_n576));
  OAI22_X1  g390(.A1(new_n569), .A2(new_n571), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT94), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n217), .A2(G143), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n217), .B2(G143), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n210), .A2(KEYINPUT96), .A3(G128), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n259), .B(new_n580), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G122), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G116), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n396), .A2(G122), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(G107), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n193), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n584), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n592));
  OAI21_X1  g406(.A(KEYINPUT97), .B1(new_n592), .B2(new_n580), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n579), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n580), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n582), .A2(new_n583), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n593), .A2(new_n596), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n591), .B1(new_n599), .B2(G134), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n580), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G134), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n584), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n193), .B1(new_n586), .B2(KEYINPUT14), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n605), .A2(new_n589), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n589), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n311), .A2(new_n318), .A3(G953), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n601), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n611), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n608), .B1(new_n603), .B2(new_n584), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n613), .B1(new_n614), .B2(new_n600), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G478), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(KEYINPUT15), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n616), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(G234), .A2(G237), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n620), .A2(G952), .A3(new_n188), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n620), .A2(G902), .A3(G953), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT21), .B(G898), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AND4_X1   g439(.A1(new_n572), .A2(new_n578), .A3(new_n619), .A4(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n520), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n317), .A2(new_n466), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  NAND2_X1  g443(.A1(new_n459), .A2(new_n302), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G472), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n461), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n374), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n317), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n611), .B1(new_n601), .B2(new_n610), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n614), .A2(new_n600), .A3(new_n613), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n302), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(KEYINPUT98), .A3(new_n617), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n616), .B2(G478), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT33), .B1(new_n636), .B2(new_n637), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n612), .A2(new_n615), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n617), .A2(G902), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n639), .A2(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI211_X1 g461(.A(new_n624), .B(new_n647), .C1(new_n578), .C2(new_n572), .ZN(new_n648));
  INV_X1    g462(.A(new_n469), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n501), .B2(new_n516), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n468), .B1(new_n650), .B2(new_n519), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n635), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  AOI21_X1  g469(.A(new_n570), .B1(new_n548), .B2(new_n566), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n556), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT99), .B1(new_n658), .B2(new_n569), .ZN(new_n659));
  INV_X1    g473(.A(new_n569), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n661), .A3(new_n657), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n638), .B(new_n618), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n554), .A2(new_n659), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n651), .A2(new_n625), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n635), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NOR2_X1   g482(.A1(new_n323), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n357), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n368), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n367), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n632), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n317), .A2(new_n627), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  AND3_X1   g491(.A1(new_n448), .A2(new_n451), .A3(G472), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n451), .B1(new_n448), .B2(G472), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n465), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n650), .A2(new_n519), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n467), .A3(new_n672), .ZN(new_n682));
  INV_X1    g496(.A(new_n621), .ZN(new_n683));
  INV_X1    g497(.A(new_n622), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n683), .B1(new_n684), .B2(G900), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT100), .Z(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n664), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n310), .A2(new_n315), .A3(new_n312), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n315), .B1(new_n310), .B2(new_n312), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n680), .B(new_n689), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  XOR2_X1   g507(.A(new_n686), .B(KEYINPUT39), .Z(new_n694));
  NAND2_X1  g508(.A1(new_n317), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n517), .A2(new_n519), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n698), .B(KEYINPUT38), .Z(new_n699));
  INV_X1    g513(.A(new_n455), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n440), .ZN(new_n701));
  INV_X1    g515(.A(new_n444), .ZN(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n702), .B2(new_n386), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n460), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n462), .B2(new_n464), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n578), .A2(new_n572), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n673), .A2(new_n467), .A3(new_n706), .A4(new_n663), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n699), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n696), .A2(new_n697), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  INV_X1    g524(.A(new_n647), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n706), .A2(new_n711), .A3(new_n687), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n682), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n680), .B(new_n713), .C1(new_n690), .C2(new_n691), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  INV_X1    g529(.A(new_n374), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n302), .B1(new_n306), .B2(new_n307), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G469), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n312), .A3(new_n308), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n680), .A2(new_n716), .A3(new_n652), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT101), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n721), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n665), .A2(new_n680), .A3(new_n716), .A4(new_n720), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND4_X1  g540(.A1(new_n626), .A2(new_n718), .A3(new_n312), .A4(new_n308), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n682), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n680), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NAND2_X1  g544(.A1(new_n651), .A2(new_n625), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n706), .B2(new_n663), .ZN(new_n734));
  AOI211_X1 g548(.A(KEYINPUT102), .B(new_n619), .C1(new_n578), .C2(new_n572), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n367), .A2(new_n369), .ZN(new_n737));
  OAI22_X1  g551(.A1(new_n456), .A2(new_n458), .B1(new_n440), .B2(new_n445), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n460), .A3(new_n302), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n631), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n732), .A2(new_n736), .A3(new_n741), .A4(new_n720), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND2_X1  g557(.A1(new_n681), .A2(new_n467), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n719), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n631), .A2(new_n739), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n746), .A2(new_n712), .A3(new_n673), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NAND2_X1  g563(.A1(new_n465), .A2(KEYINPUT106), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n462), .A2(new_n751), .A3(new_n464), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n453), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n737), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n517), .A2(new_n467), .A3(new_n519), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n297), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n279), .A2(new_n295), .A3(KEYINPUT104), .A4(new_n296), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n277), .A2(KEYINPUT103), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n761), .B(new_n190), .C1(new_n269), .C2(new_n276), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n759), .A2(G469), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n308), .A2(new_n763), .A3(new_n309), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n755), .A2(new_n312), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n712), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(KEYINPUT42), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n754), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n765), .A2(new_n680), .A3(new_n716), .A4(new_n766), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT105), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n773), .A3(new_n770), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n768), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n266), .ZN(G33));
  XOR2_X1   g590(.A(new_n688), .B(KEYINPUT107), .Z(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n466), .A3(new_n765), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  OR3_X1    g593(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT45), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n759), .A2(KEYINPUT45), .A3(new_n760), .A4(new_n762), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n781), .A3(G469), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n782), .B2(new_n309), .ZN(new_n783));
  INV_X1    g597(.A(new_n308), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n309), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n312), .A3(new_n694), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n711), .A2(new_n572), .A3(new_n578), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT43), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(KEYINPUT43), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n632), .A3(new_n672), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(KEYINPUT44), .A3(new_n632), .A4(new_n672), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n755), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n789), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(new_n262), .ZN(G39));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n787), .A2(new_n786), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n783), .A3(new_n784), .ZN(new_n803));
  INV_X1    g617(.A(new_n312), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n788), .A2(KEYINPUT47), .A3(new_n312), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n755), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n680), .A2(new_n716), .A3(new_n808), .A4(new_n712), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NAND3_X1  g625(.A1(new_n737), .A2(new_n312), .A3(new_n467), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n718), .A2(new_n308), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n790), .B(new_n812), .C1(KEYINPUT49), .C2(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n813), .A2(KEYINPUT49), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n699), .A3(new_n705), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n793), .A2(new_n621), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n720), .A2(new_n755), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n754), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT48), .ZN(new_n822));
  INV_X1    g636(.A(G952), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n817), .A2(new_n740), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n823), .B(G953), .C1(new_n824), .C2(new_n745), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n706), .A2(new_n711), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n716), .A2(new_n621), .A3(new_n705), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(new_n818), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n822), .B(new_n825), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n828), .A2(new_n706), .A3(new_n711), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n819), .A2(new_n631), .A3(new_n672), .A4(new_n739), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n699), .A2(new_n468), .A3(new_n720), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT50), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n824), .A2(new_n832), .A3(KEYINPUT50), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n830), .B(new_n831), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n805), .B(new_n806), .C1(new_n312), .C2(new_n813), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n817), .A2(new_n740), .A3(new_n808), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n829), .B1(new_n838), .B2(KEYINPUT51), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(KEYINPUT51), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n659), .A2(new_n662), .A3(new_n554), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n663), .B(KEYINPUT110), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n755), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(new_n680), .C1(new_n690), .C2(new_n691), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n746), .A2(new_n826), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n765), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n673), .A2(new_n686), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n778), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n775), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT108), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n648), .A2(new_n520), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n856), .B1(new_n648), .B2(new_n520), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n317), .A2(new_n859), .A3(new_n633), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT109), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n860), .A2(new_n628), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n860), .B2(new_n628), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n846), .A2(new_n706), .ZN(new_n864));
  INV_X1    g678(.A(new_n520), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n864), .A2(new_n865), .A3(new_n624), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n675), .B1(new_n634), .B2(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n862), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n725), .A2(new_n729), .A3(new_n721), .A4(new_n742), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n367), .A2(new_n312), .A3(new_n671), .A4(new_n687), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n764), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n705), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n744), .A2(new_n734), .A3(new_n735), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n692), .A2(new_n714), .A3(new_n875), .A4(new_n748), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n873), .B2(new_n874), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n692), .A3(new_n714), .A4(new_n748), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n855), .A2(new_n868), .A3(new_n870), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n778), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n885), .A2(new_n862), .A3(new_n863), .A4(new_n867), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n879), .A2(new_n714), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n745), .A2(new_n747), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n450), .A2(new_n452), .B1(new_n462), .B2(new_n464), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n314), .B2(new_n316), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n890), .B2(new_n689), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT111), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n887), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n880), .A2(KEYINPUT111), .ZN(new_n894));
  AOI221_X4 g708(.A(KEYINPUT112), .B1(new_n877), .B2(new_n876), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT112), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n878), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n886), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT114), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n869), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n731), .A2(new_n740), .A3(new_n719), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n903), .A2(new_n736), .B1(new_n728), .B2(new_n680), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n904), .A2(KEYINPUT114), .A3(new_n721), .A4(new_n725), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n900), .B1(new_n906), .B2(new_n775), .ZN(new_n907));
  INV_X1    g721(.A(new_n774), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n773), .B1(new_n769), .B2(new_n770), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n908), .A2(new_n909), .B1(new_n754), .B2(new_n767), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(KEYINPUT115), .A3(new_n902), .A4(new_n905), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n844), .B(new_n884), .C1(new_n899), .C2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT113), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n882), .A2(KEYINPUT53), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n895), .A2(new_n898), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n855), .A2(new_n868), .A3(new_n883), .A4(new_n870), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n915), .B(KEYINPUT54), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n913), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n892), .B1(new_n887), .B2(new_n891), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n880), .A2(KEYINPUT111), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n878), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT112), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n897), .A2(new_n896), .A3(new_n878), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n855), .A2(new_n868), .A3(new_n870), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n883), .A3(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n927), .A2(KEYINPUT113), .A3(KEYINPUT54), .A4(new_n915), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n843), .B1(new_n919), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(G952), .A2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n816), .B1(new_n929), .B2(new_n930), .ZN(G75));
  NAND2_X1  g745(.A1(new_n490), .A2(new_n492), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n498), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT55), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n907), .A2(new_n911), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n925), .A2(new_n937), .A3(new_n886), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n302), .B1(new_n938), .B2(new_n884), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n470), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT117), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT117), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n942), .A3(new_n470), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n936), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n188), .A2(G952), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT56), .B1(new_n939), .B2(G210), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n934), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n944), .A2(new_n948), .ZN(G51));
  INV_X1    g763(.A(new_n782), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n939), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT118), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n913), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n844), .B1(new_n938), .B2(new_n884), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n309), .B(KEYINPUT57), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n956), .A2(new_n957), .B1(new_n307), .B2(new_n306), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n945), .B1(new_n953), .B2(new_n958), .ZN(G54));
  NAND2_X1  g773(.A1(KEYINPUT58), .A2(G475), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT119), .Z(new_n961));
  AND3_X1   g775(.A1(new_n939), .A2(new_n567), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n567), .B1(new_n939), .B2(new_n961), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n962), .A2(new_n963), .A3(new_n945), .ZN(G60));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT59), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n919), .A2(new_n928), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n645), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(new_n966), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n954), .B2(new_n955), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(KEYINPUT120), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT120), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n973), .B(new_n970), .C1(new_n954), .C2(new_n955), .ZN(new_n974));
  AOI221_X4 g788(.A(new_n945), .B1(new_n968), .B2(new_n969), .C1(new_n972), .C2(new_n974), .ZN(G63));
  NAND2_X1  g789(.A1(new_n938), .A2(new_n884), .ZN(new_n976));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT60), .Z(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n362), .A3(new_n361), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n976), .A2(new_n670), .A3(new_n978), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n946), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n980), .A2(KEYINPUT61), .A3(new_n946), .A4(new_n981), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G66));
  NAND2_X1  g800(.A1(new_n868), .A2(new_n870), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n188), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n623), .B2(new_n496), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(KEYINPUT121), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(KEYINPUT121), .B2(new_n988), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n932), .B1(G898), .B2(new_n188), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n991), .B(new_n992), .Z(G69));
  AND2_X1   g807(.A1(new_n891), .A2(new_n714), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n820), .A2(new_n874), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n789), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n799), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n810), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n910), .A2(new_n778), .ZN(new_n999));
  OR2_X1    g813(.A1(new_n999), .A2(KEYINPUT123), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(KEYINPUT123), .ZN(new_n1001));
  AOI211_X1 g815(.A(new_n996), .B(new_n998), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n188), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n454), .B(new_n558), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(G900), .B2(G953), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n799), .B1(new_n807), .B2(new_n809), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n808), .B1(new_n864), .B2(new_n826), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n317), .A2(new_n466), .A3(new_n694), .A4(new_n1008), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n709), .A2(KEYINPUT62), .A3(new_n994), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT62), .B1(new_n709), .B2(new_n994), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1007), .B(new_n1009), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n188), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT122), .B1(new_n1013), .B2(new_n1004), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1006), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G72));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n927), .A2(new_n915), .ZN(new_n1019));
  OAI21_X1  g833(.A(KEYINPUT125), .B1(new_n700), .B2(new_n386), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(new_n424), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT126), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1023), .B1(new_n1012), .B2(new_n987), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT124), .ZN(new_n1028));
  INV_X1    g842(.A(new_n701), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1028), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n1026), .B(new_n946), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n987), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1002), .A2(new_n1033), .ZN(new_n1034));
  AOI211_X1 g848(.A(new_n440), .B(new_n700), .C1(new_n1034), .C2(new_n1023), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1018), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1031), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1034), .A2(new_n1023), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1040), .A2(new_n386), .A3(new_n455), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n945), .B1(new_n1019), .B2(new_n1025), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n1039), .A2(new_n1041), .A3(KEYINPUT127), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1036), .A2(new_n1043), .ZN(G57));
endmodule


