//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT77), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G125), .ZN(new_n194));
  XOR2_X1   g008(.A(G125), .B(G140), .Z(new_n195));
  OAI211_X1 g009(.A(G146), .B(new_n194), .C1(new_n195), .C2(new_n192), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G110), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT24), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G110), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(new_n202), .B2(new_n204), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G128), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT69), .B(G119), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT76), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(KEYINPUT69), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G119), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(new_n216), .A3(G128), .ZN(new_n217));
  INV_X1    g031(.A(new_n210), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT76), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n219), .B(new_n220), .C1(new_n206), .C2(new_n207), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n213), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(new_n217), .B2(new_n218), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n214), .A2(new_n216), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT23), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n224), .A2(new_n227), .A3(G110), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n200), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n194), .B1(new_n195), .B2(new_n192), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n198), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n231), .A2(new_n196), .B1(new_n208), .B2(new_n212), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT75), .B1(new_n224), .B2(new_n227), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G110), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n224), .A2(new_n227), .A3(KEYINPUT75), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n229), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n229), .B2(new_n236), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n191), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G902), .ZN(new_n241));
  INV_X1    g055(.A(new_n191), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n229), .A2(new_n236), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(KEYINPUT78), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n240), .A2(KEYINPUT25), .A3(new_n241), .A4(new_n244), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT73), .B(G217), .Z(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G234), .B2(new_n241), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n240), .A2(new_n244), .ZN(new_n253));
  OR2_X1    g067(.A1(new_n253), .A2(KEYINPUT79), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(KEYINPUT79), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n251), .A2(G902), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n252), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n198), .A2(G143), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT65), .B(G143), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(new_n198), .ZN(new_n262));
  AND2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT66), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(G137), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT11), .A3(G134), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(G137), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G131), .ZN(new_n275));
  INV_X1    g089(.A(G131), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n270), .A2(new_n272), .A3(new_n276), .A4(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n279));
  OR2_X1    g093(.A1(KEYINPUT65), .A2(G143), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT65), .A2(G143), .ZN(new_n281));
  AOI21_X1  g095(.A(G146), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n279), .B(new_n265), .C1(new_n282), .C2(new_n260), .ZN(new_n283));
  INV_X1    g097(.A(G143), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G146), .ZN(new_n285));
  AND2_X1   g099(.A1(KEYINPUT65), .A2(G143), .ZN(new_n286));
  NOR2_X1   g100(.A1(KEYINPUT65), .A2(G143), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n285), .B1(new_n288), .B2(G146), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n263), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n267), .A2(new_n278), .A3(new_n283), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n198), .A2(G143), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n292), .B(new_n293), .C1(new_n261), .C2(new_n198), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n226), .B1(new_n292), .B2(KEYINPUT1), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n262), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT67), .B1(new_n269), .B2(G137), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n273), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n269), .A2(KEYINPUT67), .A3(G137), .ZN(new_n299));
  OAI21_X1  g113(.A(G131), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n277), .A3(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT2), .B(G113), .Z(new_n302));
  NAND3_X1  g116(.A1(new_n214), .A2(new_n216), .A3(G116), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n209), .A2(G116), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n291), .A2(new_n301), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n291), .A2(new_n301), .A3(new_n307), .A4(KEYINPUT70), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n291), .A2(new_n301), .ZN(new_n312));
  INV_X1    g126(.A(new_n307), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT28), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n317));
  INV_X1    g131(.A(G210), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n318), .A2(G237), .A3(G953), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n317), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G101), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n308), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n316), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n329));
  NAND2_X1  g143(.A1(new_n312), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT68), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n312), .A2(new_n332), .A3(new_n329), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n291), .A2(new_n301), .A3(KEYINPUT30), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n331), .A2(new_n313), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n310), .A2(new_n311), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n323), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n328), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n241), .B1(new_n326), .B2(new_n327), .ZN(new_n339));
  OAI21_X1  g153(.A(G472), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n323), .A3(new_n336), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT31), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n316), .A2(new_n325), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n322), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT31), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n335), .A2(new_n345), .A3(new_n323), .A4(new_n336), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(G472), .A2(G902), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(KEYINPUT32), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n340), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n348), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT32), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n347), .A2(KEYINPUT72), .A3(new_n348), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n259), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT9), .B(G234), .ZN(new_n359));
  OAI21_X1  g173(.A(G221), .B1(new_n359), .B2(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G140), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n187), .A2(G227), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(G107), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(G101), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n267), .A2(new_n283), .A3(new_n290), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(G101), .ZN(new_n375));
  INV_X1    g189(.A(G101), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n366), .A2(new_n369), .A3(new_n376), .A4(new_n370), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(KEYINPUT4), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT80), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n375), .A2(new_n380), .A3(KEYINPUT4), .A4(new_n377), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n374), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT1), .ZN(new_n384));
  OAI21_X1  g198(.A(G128), .B1(new_n285), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n282), .B2(new_n260), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n383), .B1(new_n386), .B2(new_n294), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n365), .A2(G107), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n368), .A2(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(G101), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n377), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n292), .B1(new_n261), .B2(new_n198), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n384), .B1(new_n261), .B2(new_n198), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n394), .B1(new_n395), .B2(new_n226), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n391), .B1(new_n396), .B2(new_n294), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n393), .B1(new_n397), .B2(KEYINPUT10), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n382), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n278), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n364), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n198), .B1(new_n286), .B2(new_n287), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n226), .B1(new_n402), .B2(KEYINPUT1), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n294), .B1(new_n403), .B2(new_n289), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n392), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n386), .A2(new_n391), .A3(new_n294), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT12), .B1(new_n407), .B2(new_n278), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT12), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n409), .B(new_n400), .C1(new_n405), .C2(new_n406), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n408), .A2(new_n410), .A3(KEYINPUT82), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n412));
  INV_X1    g226(.A(new_n406), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n278), .B1(new_n397), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n409), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n407), .A2(KEYINPUT12), .A3(new_n278), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n401), .B1(new_n411), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT81), .B1(new_n382), .B2(new_n398), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n405), .A2(new_n383), .B1(new_n392), .B2(new_n387), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n379), .A2(new_n381), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n422), .B(new_n423), .C1(new_n424), .C2(new_n374), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n425), .A3(new_n278), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n399), .A2(new_n400), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n364), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT82), .B1(new_n408), .B2(new_n410), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n415), .A2(new_n412), .A3(new_n416), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT83), .A3(new_n401), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n420), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G469), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n241), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(new_n241), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n415), .A2(new_n416), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n427), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n364), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n426), .A2(new_n401), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n437), .B1(new_n442), .B2(G469), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n361), .B1(new_n436), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G214), .B1(G237), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n267), .A2(G125), .A3(new_n283), .A4(new_n290), .ZN(new_n449));
  INV_X1    g263(.A(G125), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n296), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n187), .A2(G224), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT85), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT87), .ZN(new_n458));
  XNOR2_X1  g272(.A(G110), .B(G122), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT84), .B1(new_n303), .B2(KEYINPUT5), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n303), .A2(KEYINPUT5), .A3(new_n304), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT84), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT5), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n211), .A2(new_n462), .A3(new_n463), .A4(G116), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n460), .A2(new_n461), .A3(G113), .A4(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n305), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n392), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n373), .B1(new_n305), .B2(new_n306), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n459), .B(new_n467), .C1(new_n424), .C2(new_n468), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n452), .A2(new_n456), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n452), .A2(new_n471), .A3(new_n456), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n458), .A2(new_n469), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(new_n466), .A3(new_n391), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n459), .B(KEYINPUT8), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n461), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n460), .A2(G113), .A3(new_n464), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n479), .B2(new_n478), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n466), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n476), .B1(new_n482), .B2(new_n392), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n241), .B1(new_n473), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n459), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n468), .B1(new_n379), .B2(new_n381), .ZN(new_n486));
  INV_X1    g300(.A(new_n467), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n469), .A2(new_n488), .A3(KEYINPUT6), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n490), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n452), .B(new_n455), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n448), .B1(new_n484), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n483), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n458), .A2(new_n472), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n469), .A2(new_n470), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(new_n241), .A3(new_n499), .A4(new_n447), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n446), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n231), .A2(new_n196), .ZN(new_n502));
  INV_X1    g316(.A(G214), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n503), .A2(G237), .A3(G953), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT88), .B1(new_n261), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n506));
  INV_X1    g320(.A(G237), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n187), .A3(G214), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n288), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n508), .B2(new_n284), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(KEYINPUT89), .A3(G143), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n505), .A2(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n276), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n502), .B1(new_n514), .B2(KEYINPUT17), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n511), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n261), .A2(new_n504), .A3(KEYINPUT88), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n506), .B1(new_n288), .B2(new_n508), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G131), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n513), .A2(new_n276), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G113), .B(G122), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(new_n365), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT91), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n199), .B(G146), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(new_n276), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n528), .B1(new_n513), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n519), .A2(KEYINPUT18), .A3(G131), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n532), .B2(new_n533), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n524), .B(new_n527), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n528), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n519), .B2(new_n530), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n513), .A2(new_n529), .A3(new_n276), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT90), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n542), .A2(new_n535), .B1(new_n523), .B2(new_n515), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n538), .B1(new_n543), .B2(new_n526), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n241), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G475), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n520), .A2(new_n521), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n199), .B(KEYINPUT19), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n197), .B1(new_n198), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n542), .A2(new_n535), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n538), .B1(new_n550), .B2(new_n526), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT20), .ZN(new_n552));
  NOR2_X1   g366(.A1(G475), .A2(G902), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n546), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n288), .A2(G128), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n226), .A2(G143), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n269), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G116), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(new_n368), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n557), .A2(KEYINPUT13), .A3(new_n558), .ZN(new_n562));
  OAI21_X1  g376(.A(G134), .B1(new_n557), .B2(KEYINPUT13), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n559), .B(new_n561), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT14), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G122), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G116), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n368), .B1(new_n568), .B2(KEYINPUT14), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n566), .A2(new_n569), .B1(new_n368), .B2(new_n560), .ZN(new_n570));
  INV_X1    g384(.A(new_n559), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n269), .B1(new_n557), .B2(new_n558), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n250), .A2(G953), .A3(new_n359), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n564), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n564), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n241), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G478), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT15), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n580), .A2(KEYINPUT92), .A3(new_n581), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G952), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(KEYINPUT93), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(KEYINPUT93), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n187), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(G234), .B2(G237), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT94), .ZN(new_n592));
  NAND2_X1  g406(.A1(G234), .A2(G237), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(G902), .A3(G953), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT95), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT21), .B(G898), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n556), .A2(new_n586), .A3(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n444), .A2(new_n501), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n358), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  INV_X1    g416(.A(new_n251), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n247), .B2(new_n248), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n254), .A2(new_n255), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n604), .B1(new_n605), .B2(new_n257), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n444), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n347), .B2(new_n241), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n354), .A3(new_n356), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT96), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n551), .A2(new_n553), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT20), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n615), .A2(new_n616), .B1(G475), .B2(new_n545), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n578), .A2(new_n241), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n577), .B2(G478), .ZN(new_n620));
  OR3_X1    g434(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT33), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT33), .B1(new_n575), .B2(new_n576), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n620), .B1(new_n623), .B2(G478), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n446), .B(new_n598), .C1(new_n494), .C2(new_n500), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n613), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NAND2_X1  g446(.A1(new_n494), .A2(new_n500), .ZN(new_n633));
  INV_X1    g447(.A(new_n598), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n445), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n617), .A2(new_n586), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n613), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n242), .A2(KEYINPUT36), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n229), .B2(new_n236), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n229), .A2(new_n236), .A3(new_n642), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n645), .ZN(new_n647));
  INV_X1    g461(.A(new_n641), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n647), .A2(new_n648), .A3(new_n643), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n257), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n644), .A2(new_n641), .A3(new_n645), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n648), .B1(new_n647), .B2(new_n643), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(KEYINPUT98), .A3(new_n257), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n252), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  AND4_X1   g471(.A1(new_n501), .A2(new_n444), .A3(new_n599), .A4(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n611), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n436), .A2(new_n443), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n501), .A3(new_n360), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n357), .B2(new_n351), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n652), .A2(new_n656), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n604), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n595), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n592), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n667), .A2(new_n636), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XOR2_X1   g487(.A(new_n633), .B(KEYINPUT38), .Z(new_n674));
  NAND4_X1  g488(.A1(new_n667), .A2(new_n445), .A3(new_n556), .A4(new_n586), .ZN(new_n675));
  INV_X1    g489(.A(new_n444), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n670), .B(KEYINPUT39), .Z(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AOI211_X1 g494(.A(new_n674), .B(new_n675), .C1(new_n680), .C2(KEYINPUT40), .ZN(new_n681));
  INV_X1    g495(.A(new_n357), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n335), .A2(new_n336), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n322), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n241), .B1(new_n315), .B2(new_n323), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n349), .A2(new_n686), .ZN(new_n687));
  OAI221_X1 g501(.A(new_n681), .B1(KEYINPUT40), .B2(new_n680), .C1(new_n682), .C2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n261), .ZN(G45));
  NAND2_X1  g503(.A1(new_n351), .A2(new_n357), .ZN(new_n690));
  INV_X1    g504(.A(new_n670), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n556), .A2(new_n624), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n667), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n690), .A2(new_n501), .A3(new_n444), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  AND3_X1   g509(.A1(new_n432), .A2(KEYINPUT83), .A3(new_n401), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT83), .B1(new_n432), .B2(new_n401), .ZN(new_n697));
  INV_X1    g511(.A(new_n364), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n426), .B2(new_n427), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n360), .A3(new_n436), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n358), .A2(new_n703), .A3(new_n629), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND3_X1  g520(.A1(new_n358), .A2(new_n703), .A3(new_n637), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT99), .B(G116), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G18));
  AND3_X1   g523(.A1(new_n434), .A2(new_n435), .A3(new_n241), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n435), .B1(new_n434), .B2(new_n241), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT100), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n501), .A4(new_n360), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n701), .A2(new_n501), .A3(new_n360), .A4(new_n436), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT101), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n657), .A2(new_n599), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n357), .B2(new_n351), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n718), .B1(new_n717), .B2(new_n720), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n209), .ZN(G21));
  NAND3_X1  g538(.A1(new_n627), .A2(new_n556), .A3(new_n586), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n702), .ZN(new_n726));
  INV_X1    g540(.A(new_n352), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n259), .A2(new_n727), .A3(new_n609), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NOR2_X1   g544(.A1(new_n727), .A2(new_n609), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n693), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(new_n692), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n633), .A2(new_n446), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n444), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT32), .B1(new_n347), .B2(new_n348), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n606), .B(new_n741), .C1(new_n350), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n352), .A2(new_n355), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n349), .A3(new_n340), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n741), .B1(new_n746), .B2(new_n606), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n740), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n663), .A2(new_n360), .A3(new_n738), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n358), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n751));
  AOI22_X1  g565(.A1(KEYINPUT42), .A2(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  NOR2_X1   g567(.A1(new_n636), .A2(new_n670), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n358), .A2(new_n754), .A3(new_n749), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n625), .B1(new_n556), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n757), .B2(new_n556), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT43), .ZN(new_n760));
  OR3_X1    g574(.A1(new_n556), .A2(new_n625), .A3(KEYINPUT43), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n611), .A3(new_n657), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(KEYINPUT107), .A3(new_n763), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n761), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(KEYINPUT43), .B2(new_n759), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(KEYINPUT44), .A3(new_n611), .A4(new_n657), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n738), .B(KEYINPUT105), .Z(new_n772));
  AND3_X1   g586(.A1(new_n771), .A2(KEYINPUT106), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT106), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n768), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n768), .B(KEYINPUT108), .C1(new_n773), .C2(new_n774), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n442), .A2(KEYINPUT45), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n440), .A2(new_n441), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n435), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n437), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT103), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n437), .B1(new_n779), .B2(new_n782), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n710), .B1(new_n789), .B2(KEYINPUT46), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT103), .B1(new_n789), .B2(KEYINPUT46), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n360), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n678), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n777), .A2(new_n778), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  AND3_X1   g610(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n360), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT47), .B1(new_n792), .B2(new_n360), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n737), .A2(new_n259), .A3(new_n738), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n801));
  OR3_X1    g615(.A1(new_n690), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n690), .B2(new_n800), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n193), .ZN(G42));
  INV_X1    g620(.A(new_n592), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n770), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n808), .A2(new_n703), .A3(new_n738), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n744), .A2(new_n747), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT48), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n703), .A2(new_n606), .A3(new_n807), .A4(new_n738), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n682), .A3(new_n687), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n626), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n808), .A2(new_n728), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n590), .B1(new_n816), .B2(new_n717), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n812), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n703), .A2(new_n674), .A3(new_n446), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n808), .A2(new_n728), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n823));
  NAND2_X1  g637(.A1(new_n617), .A2(new_n625), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n822), .A2(new_n823), .B1(new_n814), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n667), .A2(new_n727), .A3(new_n609), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n821), .A2(new_n827), .B1(new_n809), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT115), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n798), .B(new_n797), .C1(new_n361), .C2(new_n712), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n816), .A2(KEYINPUT115), .A3(new_n772), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n831), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n826), .B2(new_n829), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT51), .B1(new_n839), .B2(new_n835), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n818), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n501), .A2(new_n556), .A3(new_n586), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n842), .A2(new_n657), .A3(new_n670), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n843), .B(new_n444), .C1(new_n687), .C2(new_n682), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n735), .A2(new_n672), .A3(new_n694), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT52), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n748), .A2(KEYINPUT42), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n731), .A2(new_n657), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n739), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n749), .A2(new_n828), .A3(KEYINPUT113), .A4(new_n737), .ZN(new_n856));
  INV_X1    g670(.A(new_n582), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n617), .A2(new_n857), .A3(new_n691), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n444), .A2(new_n859), .A3(new_n657), .A4(new_n738), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n855), .A2(new_n856), .B1(new_n690), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n358), .A2(new_n749), .A3(new_n751), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n852), .A2(new_n861), .A3(new_n862), .A4(new_n755), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n658), .A2(new_n659), .B1(new_n726), .B2(new_n728), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n358), .B(new_n703), .C1(new_n629), .C2(new_n637), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n546), .B(new_n582), .C1(new_n554), .C2(new_n555), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n635), .A2(KEYINPUT112), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n868));
  INV_X1    g682(.A(new_n866), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n627), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n628), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n612), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n864), .A2(new_n865), .A3(new_n601), .A4(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n863), .A2(new_n723), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT53), .B1(new_n851), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n845), .A2(new_n849), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n717), .A2(new_n732), .B1(new_n665), .B2(new_n671), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(KEYINPUT52), .A3(new_n694), .A4(new_n844), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n723), .A2(new_n873), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n852), .A2(new_n861), .A3(new_n862), .A4(new_n755), .ZN(new_n881));
  AND4_X1   g695(.A1(KEYINPUT53), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT54), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n851), .A2(new_n874), .A3(KEYINPUT53), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n876), .A2(new_n878), .ZN(new_n886));
  INV_X1    g700(.A(new_n873), .ZN(new_n887));
  INV_X1    g701(.A(new_n722), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n855), .A2(new_n856), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n860), .A2(new_n690), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n891), .A2(new_n755), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n887), .A2(new_n890), .A3(new_n752), .A4(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n885), .B1(new_n886), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n884), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n841), .A2(new_n883), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(G952), .B2(G953), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n759), .A2(new_n259), .A3(new_n446), .A4(new_n361), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n901), .A2(KEYINPUT110), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT49), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n674), .B1(new_n712), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n901), .B2(KEYINPUT110), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n682), .A2(new_n687), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n712), .A2(new_n903), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT111), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n902), .A2(new_n905), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n899), .A2(new_n909), .ZN(G75));
  NAND2_X1  g724(.A1(new_n489), .A2(new_n491), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n492), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT55), .Z(new_n913));
  AOI21_X1  g727(.A(new_n241), .B1(new_n884), .B2(new_n895), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(G210), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n915), .B2(KEYINPUT56), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n187), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n915), .A2(KEYINPUT56), .A3(new_n913), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(G51));
  XNOR2_X1  g735(.A(new_n434), .B(KEYINPUT117), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n849), .B1(new_n845), .B2(new_n846), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n925), .A2(new_n885), .A3(new_n894), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT53), .B1(new_n874), .B2(new_n879), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT54), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n897), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n437), .B(KEYINPUT57), .Z(new_n931));
  OAI21_X1  g745(.A(new_n922), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n241), .B(new_n783), .C1(new_n884), .C2(new_n895), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT118), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n917), .B1(new_n932), .B2(new_n934), .ZN(G54));
  AND2_X1   g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n914), .A2(new_n551), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n551), .B1(new_n914), .B2(new_n936), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n917), .ZN(G60));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n618), .B(KEYINPUT59), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n883), .B2(new_n897), .ZN(new_n942));
  INV_X1    g756(.A(new_n623), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n623), .A2(new_n941), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT119), .B1(new_n929), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT119), .ZN(new_n947));
  INV_X1    g761(.A(new_n945), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n947), .B(new_n948), .C1(new_n928), .C2(new_n897), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n944), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n941), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n884), .A2(new_n895), .A3(new_n896), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n885), .B1(new_n925), .B2(new_n894), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n874), .A2(KEYINPUT53), .A3(new_n879), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n896), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n951), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(KEYINPUT120), .A3(new_n623), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n918), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n950), .A2(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(new_n884), .A2(new_n895), .ZN(new_n960));
  XOR2_X1   g774(.A(KEYINPUT121), .B(KEYINPUT60), .Z(new_n961));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n917), .B1(new_n964), .B2(new_n256), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n655), .B(KEYINPUT122), .Z(new_n967));
  NAND4_X1  g781(.A1(new_n960), .A2(new_n966), .A3(new_n963), .A4(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n960), .A2(new_n963), .A3(new_n967), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT123), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n965), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n965), .A2(new_n970), .A3(KEYINPUT61), .A4(new_n968), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(G66));
  INV_X1    g789(.A(G224), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n596), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n880), .B2(G953), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n911), .B1(G898), .B2(new_n187), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G69));
  NAND3_X1  g794(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(new_n548), .Z(new_n982));
  AOI21_X1  g796(.A(G227), .B1(new_n982), .B2(KEYINPUT126), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n983), .B2(new_n668), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(G227), .B2(new_n187), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n735), .A2(new_n672), .A3(new_n694), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT124), .ZN(new_n987));
  INV_X1    g801(.A(new_n805), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n793), .A2(new_n678), .A3(new_n842), .ZN(new_n989));
  AOI22_X1  g803(.A1(new_n989), .A2(new_n810), .B1(new_n754), .B2(new_n750), .ZN(new_n990));
  AND4_X1   g804(.A1(new_n752), .A2(new_n987), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n795), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n985), .B1(new_n992), .B2(new_n187), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n738), .B1(new_n626), .B2(new_n869), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n680), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n805), .B1(new_n358), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n795), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n987), .A2(KEYINPUT62), .A3(new_n688), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT62), .B1(new_n987), .B2(new_n688), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(KEYINPUT125), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1000), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n998), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT125), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1004), .A2(new_n1005), .A3(new_n795), .A4(new_n996), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n982), .A2(G953), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n993), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT126), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n984), .B1(new_n1009), .B2(new_n1010), .ZN(G72));
  AND2_X1   g825(.A1(new_n683), .A2(new_n322), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n795), .A2(new_n991), .A3(new_n880), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  AND3_X1   g830(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1014), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1012), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n953), .A2(new_n954), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1016), .ZN(new_n1021));
  INV_X1    g835(.A(new_n337), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1021), .B1(new_n1022), .B2(new_n341), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n917), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n684), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1002), .A2(new_n880), .A3(new_n1006), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1026), .B1(new_n1027), .B2(new_n1016), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1025), .A2(new_n1028), .ZN(G57));
endmodule


