//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n544,
    new_n545, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT68), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n461), .A2(KEYINPUT68), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n462), .B(new_n463), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT69), .B1(new_n468), .B2(G2105), .ZN(new_n471));
  OR2_X1    g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n473), .C1(new_n464), .C2(new_n465), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n475), .ZN(new_n477));
  INV_X1    g052(.A(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n476), .A2(new_n477), .B1(G101), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n472), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n466), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n466), .A2(new_n473), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NOR2_X1   g064(.A1(new_n473), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT71), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OR3_X1    g067(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT71), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n492), .A2(new_n493), .B1(new_n484), .B2(G126), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n473), .C1(new_n464), .C2(new_n465), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT4), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n494), .A2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G50), .ZN(new_n502));
  XOR2_X1   g077(.A(new_n502), .B(KEYINPUT72), .Z(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n498), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n503), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n513), .A2(new_n514), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n521), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n524), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n509), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n522), .A2(new_n532), .B1(new_n515), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(new_n501), .A2(G43), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n507), .A2(new_n521), .A3(G81), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n509), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  INV_X1    g121(.A(G91), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT75), .B1(new_n515), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n507), .A2(new_n521), .A3(new_n549), .A4(G91), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(KEYINPUT74), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n501), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n554), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n525), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n551), .A2(new_n558), .A3(new_n562), .ZN(G299));
  OR2_X1    g138(.A1(new_n531), .A2(new_n534), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  AOI22_X1  g140(.A1(new_n499), .A2(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G87), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT76), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n507), .A2(G74), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n501), .B2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n509), .ZN(new_n573));
  INV_X1    g148(.A(G48), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n522), .A2(new_n574), .B1(new_n515), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n566), .A2(G85), .B1(new_n501), .B2(G47), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n509), .B2(new_n580), .ZN(G290));
  INV_X1    g156(.A(G868), .ZN(new_n582));
  NOR2_X1   g157(.A1(G301), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G66), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n587), .C1(new_n513), .C2(new_n514), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n588), .A2(KEYINPUT78), .A3(new_n589), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n592), .A2(G651), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n521), .A2(G54), .A3(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n515), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n507), .A2(new_n521), .A3(KEYINPUT10), .A4(G92), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT79), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n583), .B1(new_n603), .B2(new_n582), .ZN(G284));
  AOI21_X1  g179(.A(new_n583), .B1(new_n603), .B2(new_n582), .ZN(G321));
  NAND2_X1  g180(.A1(G299), .A2(new_n582), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n582), .B2(G168), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n582), .B2(G168), .ZN(G280));
  XNOR2_X1  g183(.A(KEYINPUT80), .B(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n603), .B1(G860), .B2(new_n609), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT81), .Z(G148));
  NOR2_X1   g186(.A1(new_n539), .A2(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n603), .A2(new_n609), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT82), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n612), .B1(new_n615), .B2(G868), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g192(.A1(new_n464), .A2(new_n465), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n479), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT12), .Z(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT13), .Z(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n482), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n484), .A2(G123), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n623), .A2(new_n624), .A3(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n638), .ZN(new_n640));
  NAND4_X1  g215(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n639), .A2(new_n645), .A3(new_n641), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(G14), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n651), .A3(new_n648), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  OR3_X1    g237(.A1(new_n661), .A2(KEYINPUT85), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(KEYINPUT85), .B1(new_n661), .B2(new_n662), .ZN(new_n664));
  INV_X1    g239(.A(new_n659), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n660), .B(KEYINPUT17), .Z(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n664), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n662), .A2(new_n659), .A3(new_n660), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n662), .A3(new_n665), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT87), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT88), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(new_n680), .ZN(new_n685));
  MUX2_X1   g260(.A(new_n685), .B(new_n684), .S(new_n677), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT90), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT89), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n690), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT94), .Z(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G303), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1971), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT95), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n698), .A2(G23), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G288), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT33), .B(G1976), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT93), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G6), .A2(G16), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n577), .B2(G16), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n707), .A2(new_n709), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n710), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n704), .A2(new_n705), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G24), .B(G290), .S(G16), .Z(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1986), .Z(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n482), .A2(G131), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n484), .A2(G119), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n473), .A2(G107), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n724), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT91), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT92), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n723), .B1(new_n731), .B2(new_n722), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n721), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n732), .B2(new_n734), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n719), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n717), .A2(new_n718), .ZN(new_n738));
  OR3_X1    g313(.A1(new_n737), .A2(KEYINPUT36), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT36), .B1(new_n737), .B2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n722), .A2(G33), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT96), .B(KEYINPUT25), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n618), .A2(new_n473), .ZN(new_n747));
  INV_X1    g322(.A(G139), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND2_X1  g327(.A1(G115), .A2(G2104), .ZN(new_n753));
  INV_X1    g328(.A(G127), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n466), .B2(new_n754), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n751), .A2(new_n752), .B1(G2105), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n742), .B1(new_n756), .B2(new_n722), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G2072), .ZN(new_n758));
  INV_X1    g333(.A(G2090), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n722), .A2(G35), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n722), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT29), .Z(new_n762));
  OAI21_X1  g337(.A(new_n758), .B1(new_n759), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G2072), .B2(new_n757), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT31), .B(G11), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(G28), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n722), .B1(new_n766), .B2(G28), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n629), .A2(new_n722), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n765), .B1(new_n767), .B2(new_n768), .C1(new_n769), .C2(KEYINPUT101), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(KEYINPUT101), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g346(.A1(G168), .A2(new_n698), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n698), .B2(G21), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G5), .A2(G16), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G171), .B2(G16), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n774), .A2(G1966), .B1(G1961), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G1966), .ZN(new_n778));
  INV_X1    g353(.A(new_n776), .ZN(new_n779));
  INV_X1    g354(.A(G1961), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n773), .A2(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G19), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n540), .B2(G16), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1341), .Z(new_n784));
  NAND4_X1  g359(.A1(new_n771), .A2(new_n777), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(G164), .A2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G27), .B2(G29), .ZN(new_n787));
  INV_X1    g362(.A(G2078), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n722), .A2(G26), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n482), .A2(G140), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n484), .A2(G128), .ZN(new_n793));
  OR2_X1    g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n794), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n791), .B1(new_n797), .B2(new_n722), .ZN(new_n798));
  INV_X1    g373(.A(G2067), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n787), .A2(new_n788), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n785), .A2(new_n789), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n698), .A2(G4), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n603), .B2(new_n698), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  AND3_X1   g382(.A1(new_n764), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n722), .A2(G32), .ZN(new_n809));
  NAND3_X1  g384(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT99), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n482), .A2(G141), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n484), .A2(G129), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n479), .A2(G105), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT100), .ZN(new_n818));
  OR3_X1    g393(.A1(new_n813), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n813), .B2(new_n817), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n809), .B1(new_n822), .B2(new_n722), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT27), .Z(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(G1996), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n762), .A2(new_n759), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT102), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n698), .A2(G20), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT23), .Z(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G299), .B2(G16), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1956), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n832));
  INV_X1    g407(.A(G34), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n722), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  OAI22_X1  g410(.A1(G160), .A2(new_n722), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G2084), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n827), .A2(new_n831), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G1996), .B2(new_n824), .ZN(new_n840));
  AND4_X1   g415(.A1(new_n741), .A2(new_n808), .A3(new_n825), .A4(new_n840), .ZN(G311));
  NAND4_X1  g416(.A1(new_n741), .A2(new_n808), .A3(new_n825), .A4(new_n840), .ZN(G150));
  NAND2_X1  g417(.A1(new_n603), .A2(G559), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT38), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n501), .A2(G55), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n507), .A2(new_n521), .A3(G93), .ZN(new_n846));
  AND2_X1   g421(.A1(G80), .A2(G543), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n507), .B2(G67), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n845), .B(new_n846), .C1(new_n848), .C2(new_n509), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n539), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n539), .A2(new_n849), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n844), .B(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(KEYINPUT39), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n855), .A2(new_n856), .A3(G860), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n849), .A2(G860), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  INV_X1    g435(.A(new_n729), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n819), .A2(new_n797), .A3(new_n820), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n797), .B1(new_n819), .B2(new_n820), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n729), .A3(new_n862), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n484), .A2(G130), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT104), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G118), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n871), .A2(new_n872), .B1(new_n874), .B2(G2105), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n482), .A2(G142), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n620), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n751), .A2(new_n752), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n755), .A2(G2105), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n494), .A2(new_n496), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n756), .A2(G164), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n877), .B(new_n620), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n756), .A2(G164), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n868), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n865), .A2(new_n886), .A3(new_n867), .A4(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n488), .B(new_n629), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(KEYINPUT103), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n896), .A2(G160), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G160), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n892), .B(new_n893), .C1(new_n898), .C2(new_n899), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(G395));
  NAND2_X1  g481(.A1(new_n615), .A2(new_n853), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n614), .A2(new_n852), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n551), .A2(new_n558), .A3(new_n562), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n602), .ZN(new_n912));
  NAND3_X1  g487(.A1(G299), .A2(new_n594), .A3(new_n601), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(KEYINPUT107), .A3(new_n913), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n602), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n918), .B2(new_n910), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n912), .A2(new_n913), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n907), .A2(new_n908), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(G303), .B(G288), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n577), .B(G290), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n925), .B2(new_n926), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n920), .B(new_n923), .C1(new_n925), .C2(new_n926), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n928), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n928), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n849), .A2(new_n582), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(G295));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n937), .ZN(G331));
  NOR3_X1   g514(.A1(new_n850), .A2(new_n851), .A3(G171), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n538), .A2(new_n509), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n536), .A2(new_n537), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n507), .A2(G67), .ZN(new_n943));
  OAI21_X1  g518(.A(G651), .B1(new_n943), .B2(new_n847), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n566), .A2(G93), .B1(new_n501), .B2(G55), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n941), .A2(new_n942), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n539), .A2(new_n849), .ZN(new_n947));
  AOI21_X1  g522(.A(G301), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n940), .A2(new_n948), .A3(G286), .ZN(new_n949));
  OAI21_X1  g524(.A(G171), .B1(new_n850), .B2(new_n851), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(G301), .A3(new_n947), .ZN(new_n951));
  AOI21_X1  g526(.A(G168), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n921), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(G286), .B1(new_n940), .B2(new_n948), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(G168), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n919), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT109), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n953), .B(new_n959), .C1(new_n919), .C2(new_n956), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n931), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n962), .A3(new_n903), .ZN(new_n963));
  INV_X1    g538(.A(new_n931), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n957), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n962), .B1(new_n961), .B2(new_n903), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT43), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n964), .B2(new_n957), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n922), .B1(new_n956), .B2(new_n910), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n910), .B1(new_n915), .B2(new_n917), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n955), .B(new_n954), .C1(new_n973), .C2(KEYINPUT111), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n973), .A2(KEYINPUT111), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n931), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT44), .B1(new_n970), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n966), .B2(new_n968), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(new_n986), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n883), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n480), .B(G40), .C1(new_n470), .C2(new_n471), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n822), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n796), .B(G2067), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n993), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n729), .B(new_n733), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n993), .A2(new_n994), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT112), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n822), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1002), .A2(KEYINPUT113), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(KEYINPUT113), .ZN(new_n1004));
  OAI221_X1 g579(.A(new_n997), .B1(new_n998), .B2(new_n999), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(G290), .B(G1986), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n993), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT125), .ZN(new_n1008));
  INV_X1    g583(.A(G1971), .ZN(new_n1009));
  INV_X1    g584(.A(new_n992), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n883), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n991), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1009), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n989), .A2(KEYINPUT114), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n883), .A2(new_n1017), .A3(new_n988), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n992), .B1(KEYINPUT50), .B2(new_n989), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1014), .B1(new_n1021), .B2(G2090), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1025), .A3(G8), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1010), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n568), .A2(G1976), .A3(new_n570), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(G8), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n577), .B(G1981), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n577), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1033), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1027), .A2(new_n1032), .A3(new_n1037), .A4(G8), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT115), .B(G1976), .Z(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(G288), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1027), .A2(G8), .A3(new_n1028), .A4(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1026), .A2(new_n1030), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n989), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n992), .B1(new_n1044), .B2(new_n1016), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1017), .B1(new_n883), .B2(new_n988), .ZN(new_n1046));
  AOI211_X1 g621(.A(KEYINPUT114), .B(G1384), .C1(new_n494), .C2(new_n496), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT50), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1048), .A3(new_n759), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1014), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1025), .B1(new_n1050), .B2(G8), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1008), .B1(new_n1043), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1042), .A2(new_n1030), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1051), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(KEYINPUT125), .A4(new_n1026), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT53), .B1(new_n1057), .B2(new_n788), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n780), .B2(new_n1021), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1012), .B1(new_n1060), .B2(new_n990), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n788), .A2(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(G301), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1052), .A2(new_n1056), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(KEYINPUT124), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1019), .A2(new_n1020), .A3(new_n837), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1069), .B(G168), .C1(new_n1061), .C2(G1966), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1068), .B1(new_n1070), .B2(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(G8), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT124), .B(KEYINPUT51), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1012), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n990), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1966), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1069), .ZN(new_n1079));
  OAI211_X1 g654(.A(G8), .B(G286), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1069), .B1(new_n1061), .B2(G1966), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(KEYINPUT123), .A3(G8), .A4(G286), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1075), .A2(KEYINPUT62), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT62), .B1(new_n1075), .B2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1065), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(G288), .A2(G1976), .ZN(new_n1089));
  XOR2_X1   g664(.A(new_n1089), .B(KEYINPUT116), .Z(new_n1090));
  AOI21_X1  g665(.A(new_n1034), .B1(new_n1090), .B2(new_n1038), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1027), .A2(G8), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1053), .A2(new_n1026), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1083), .A2(G8), .A3(G168), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT63), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1025), .B1(new_n1022), .B2(G8), .ZN(new_n1096));
  OR3_X1    g671(.A1(new_n1095), .A2(new_n1043), .A3(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1054), .A2(new_n1055), .A3(new_n1094), .A4(new_n1026), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1093), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1088), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1071), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1070), .A2(G8), .A3(new_n1074), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1085), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1106));
  XNOR2_X1  g681(.A(G301), .B(KEYINPUT54), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n468), .A2(G2105), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n480), .A2(G40), .A3(new_n1108), .A4(new_n1062), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1013), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1110), .B2(new_n1011), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1106), .A2(new_n1107), .B1(new_n1059), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1105), .A2(new_n1052), .A3(new_n1112), .A4(new_n1056), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1021), .A2(new_n806), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(G2067), .B2(new_n1027), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n602), .A2(KEYINPUT122), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n602), .A2(KEYINPUT122), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1120), .B(new_n1121), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  OAI21_X1  g699(.A(G299), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1076), .A2(new_n991), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1956), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1128), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1057), .A2(new_n1129), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1133), .B(new_n1127), .C1(G1956), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT121), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1136), .A2(KEYINPUT121), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1057), .A2(new_n994), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(G1341), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1027), .A2(KEYINPUT119), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT119), .B1(new_n1027), .B2(new_n1145), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT120), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1148), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n1143), .A4(new_n1146), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1142), .B1(new_n1153), .B2(new_n540), .ZN(new_n1154));
  AOI211_X1 g729(.A(KEYINPUT59), .B(new_n539), .C1(new_n1149), .C2(new_n1152), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1122), .B(new_n1141), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1115), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1132), .B1(new_n1157), .B2(new_n602), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1135), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1113), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1007), .B1(new_n1102), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT46), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1001), .B(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n993), .B1(new_n821), .B2(new_n996), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1165), .A2(KEYINPUT47), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(KEYINPUT47), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n998), .A2(G1986), .A3(G290), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT48), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1166), .A2(new_n1167), .B1(new_n1005), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n730), .A2(new_n734), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n997), .B(new_n1171), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n797), .A2(new_n799), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n998), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1161), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n1178));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1179));
  NOR2_X1   g753(.A1(G227), .A2(new_n459), .ZN(new_n1180));
  INV_X1    g754(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g755(.A(new_n1179), .B1(G401), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g756(.A(new_n657), .ZN(new_n1183));
  NOR2_X1   g757(.A1(new_n1183), .A2(new_n655), .ZN(new_n1184));
  OAI211_X1 g758(.A(KEYINPUT126), .B(new_n1180), .C1(new_n1184), .C2(new_n652), .ZN(new_n1185));
  NAND4_X1  g759(.A1(new_n904), .A2(new_n1182), .A3(new_n696), .A4(new_n1185), .ZN(new_n1186));
  INV_X1    g760(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n1178), .B1(new_n985), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g762(.A(KEYINPUT127), .B(new_n1186), .C1(new_n982), .C2(new_n984), .ZN(new_n1189));
  NOR2_X1   g763(.A1(new_n1188), .A2(new_n1189), .ZN(G308));
  NAND2_X1  g764(.A1(new_n985), .A2(new_n1187), .ZN(G225));
endmodule


