//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n565, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT66), .A3(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n462), .A2(new_n477), .A3(new_n463), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT65), .B1(new_n467), .B2(new_n468), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n466), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n476), .A2(new_n482), .ZN(G160));
  AOI21_X1  g058(.A(new_n466), .B1(new_n462), .B2(new_n463), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n464), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(KEYINPUT4), .B(G138), .C1(new_n467), .C2(new_n468), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G126), .B1(new_n467), .B2(new_n468), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n466), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n478), .A2(new_n479), .A3(G138), .A4(new_n466), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(G543), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n504), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  AND2_X1   g086(.A1(G75), .A2(G543), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n503), .B(G651), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT69), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n515), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n510), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n513), .A2(new_n516), .A3(new_n525), .A4(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n524), .A2(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n527), .A2(G51), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n510), .A2(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n531), .A2(new_n532), .A3(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n523), .A2(new_n540), .B1(new_n526), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n515), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(G171));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n523), .A2(new_n546), .B1(new_n526), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n515), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(new_n510), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n524), .B2(G91), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n522), .A2(G53), .A3(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G299));
  OR2_X1    g139(.A1(new_n542), .A2(new_n544), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT70), .ZN(G301));
  NAND3_X1  g141(.A1(new_n510), .A2(new_n522), .A3(G87), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n510), .A2(G74), .ZN(new_n570));
  AOI22_X1  g145(.A1(G49), .A2(new_n527), .B1(new_n570), .B2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G288));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  INV_X1    g148(.A(G48), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n523), .A2(new_n573), .B1(new_n526), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n510), .A2(G61), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n515), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(G305));
  XNOR2_X1  g156(.A(KEYINPUT74), .B(G85), .ZN(new_n582));
  XOR2_X1   g157(.A(KEYINPUT73), .B(G47), .Z(new_n583));
  OAI22_X1  g158(.A1(new_n523), .A2(new_n582), .B1(new_n526), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n515), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND3_X1  g163(.A1(new_n510), .A2(new_n522), .A3(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n558), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n527), .B2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(G868), .ZN(new_n597));
  XNOR2_X1  g172(.A(G171), .B(KEYINPUT70), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G284));
  AOI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G286), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(G299), .B(KEYINPUT75), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G297));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G280));
  INV_X1    g180(.A(new_n596), .ZN(new_n606));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G860), .ZN(G148));
  INV_X1    g183(.A(new_n551), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(new_n601), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n596), .A2(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n601), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g188(.A1(G123), .A2(new_n484), .B1(new_n464), .B2(G135), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n466), .A2(G111), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n473), .B1(new_n615), .B2(KEYINPUT76), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT76), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n616), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  AND2_X1   g196(.A1(new_n478), .A2(new_n479), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n622), .A2(G2104), .A3(new_n466), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT12), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n621), .B1(new_n625), .B2(G2100), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(G2100), .B2(new_n625), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT77), .ZN(G156));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  AOI21_X1  g208(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT80), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n643), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(G401));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NOR2_X1   g222(.A1(G2072), .A2(G2078), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n442), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n650), .B2(KEYINPUT81), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(KEYINPUT81), .B2(new_n650), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n649), .B(KEYINPUT17), .ZN(new_n655));
  INV_X1    g230(.A(new_n647), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n652), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n650), .A2(new_n647), .A3(new_n653), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n656), .A3(new_n653), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g248(.A(new_n673), .B(new_n672), .S(new_n665), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G6), .A2(G16), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n579), .B(KEYINPUT72), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(G16), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT32), .B(G1981), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G22), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT84), .Z(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G303), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(G1971), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(G23), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n569), .A2(new_n571), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n690), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT33), .B(G1976), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n700), .A2(new_n701), .B1(new_n694), .B2(new_n693), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n689), .A2(new_n695), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(KEYINPUT34), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n689), .A2(new_n705), .A3(new_n702), .A4(new_n695), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n690), .A2(G24), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT83), .Z(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n587), .B2(new_n690), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1986), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n464), .A2(G131), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n484), .A2(G119), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n466), .A2(G107), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n711), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G25), .B(new_n715), .S(G29), .Z(new_n716));
  XOR2_X1   g291(.A(KEYINPUT35), .B(G1991), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n710), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g295(.A1(new_n706), .A2(KEYINPUT85), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(KEYINPUT85), .B1(new_n706), .B2(new_n720), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n704), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT36), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n690), .A2(G19), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n551), .B2(new_n690), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1341), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n728), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G2090), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT90), .Z(new_n733));
  INV_X1    g308(.A(G1956), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n690), .A2(G20), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT91), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT23), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G299), .B2(G16), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n727), .B(new_n733), .C1(new_n734), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n690), .A2(G21), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G168), .B2(new_n690), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT88), .B(G1966), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n728), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n484), .A2(G128), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n464), .A2(G140), .ZN(new_n747));
  OR2_X1    g322(.A1(G104), .A2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G29), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(KEYINPUT86), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(KEYINPUT86), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n745), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2067), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n738), .A2(new_n734), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n739), .A2(new_n743), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n464), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n484), .A2(G129), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(new_n728), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n728), .B2(G32), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G1996), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G164), .A2(G29), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G27), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G2078), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT24), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n728), .B1(new_n778), .B2(G34), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n778), .B2(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G160), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n772), .A2(new_n776), .A3(new_n777), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G5), .A2(G16), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT89), .Z(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n565), .B2(new_n690), .ZN(new_n788));
  INV_X1    g363(.A(G1961), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT30), .B(G28), .ZN(new_n792));
  OR2_X1    g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  NAND2_X1  g368(.A1(KEYINPUT31), .A2(G11), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n792), .A2(new_n728), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n728), .A2(G33), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n622), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(new_n466), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT25), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n464), .A2(G139), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(new_n728), .ZN(new_n804));
  OAI221_X1 g379(.A(new_n795), .B1(new_n728), .B2(new_n620), .C1(new_n804), .C2(G2072), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n791), .B(new_n805), .C1(G2072), .C2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n690), .A2(G4), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n606), .B2(new_n690), .ZN(new_n808));
  INV_X1    g383(.A(G1348), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n731), .A2(G2090), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n788), .A2(new_n789), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G2084), .B2(new_n781), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n811), .B(new_n813), .C1(new_n770), .C2(new_n771), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n785), .A2(new_n806), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n758), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n724), .A2(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  NAND3_X1  g393(.A1(new_n510), .A2(new_n522), .A3(G93), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n522), .A2(G55), .A3(G543), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT93), .ZN(new_n821));
  AOI21_X1  g396(.A(KEYINPUT93), .B1(new_n819), .B2(new_n820), .ZN(new_n822));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n510), .B2(G67), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT92), .ZN(new_n826));
  OAI21_X1  g401(.A(G651), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI211_X1 g402(.A(KEYINPUT92), .B(new_n824), .C1(new_n510), .C2(G67), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n821), .A2(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT94), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n508), .A2(new_n509), .ZN(new_n831));
  INV_X1    g406(.A(new_n505), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n831), .A2(G67), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(new_n823), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT92), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n825), .A2(new_n826), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n836), .A3(G651), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n837), .B(new_n838), .C1(new_n822), .C2(new_n821), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n830), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND3_X1  g417(.A1(new_n830), .A2(new_n609), .A3(new_n839), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n829), .A2(new_n551), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n596), .A2(new_n607), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT38), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n848), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n853));
  INV_X1    g428(.A(G860), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n852), .B2(KEYINPUT39), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n842), .B1(new_n853), .B2(new_n855), .ZN(G145));
  XNOR2_X1  g431(.A(new_n620), .B(new_n489), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G160), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n464), .A2(G142), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n484), .A2(G130), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n466), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n860), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n624), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n715), .ZN(new_n866));
  INV_X1    g441(.A(new_n750), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n768), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n767), .A2(new_n750), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n501), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n497), .A2(KEYINPUT96), .A3(new_n500), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n868), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n803), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n803), .A3(new_n876), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n866), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT98), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n866), .A3(new_n880), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n859), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n883), .B(KEYINPUT97), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n858), .B(KEYINPUT99), .Z(new_n888));
  NOR2_X1   g463(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n886), .A2(KEYINPUT40), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT40), .B1(new_n886), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(G395));
  OAI21_X1  g468(.A(new_n611), .B1(new_n846), .B2(new_n847), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n843), .A2(new_n845), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT95), .ZN(new_n896));
  INV_X1    g471(.A(new_n611), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n596), .A2(G299), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n561), .A2(new_n591), .A3(new_n595), .A4(new_n563), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT41), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n904), .A3(new_n901), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(KEYINPUT100), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n907), .A3(KEYINPUT41), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n894), .A2(new_n899), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n902), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(new_n894), .B2(new_n899), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n894), .A2(new_n899), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n902), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n910), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n686), .B(G166), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n697), .A2(new_n587), .ZN(new_n920));
  NAND2_X1  g495(.A1(G290), .A2(G288), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(KEYINPUT101), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G305), .B(G166), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(KEYINPUT101), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n921), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n914), .A2(new_n918), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n914), .B2(new_n918), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n840), .A2(new_n601), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n911), .A2(new_n913), .A3(KEYINPUT42), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n917), .B1(new_n916), .B2(new_n910), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n930), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n601), .B1(new_n941), .B2(new_n932), .ZN(new_n942));
  INV_X1    g517(.A(new_n937), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT102), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n938), .A2(new_n944), .ZN(G295));
  NAND2_X1  g520(.A1(new_n935), .A2(new_n937), .ZN(G331));
  NOR2_X1   g521(.A1(G168), .A2(G171), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n598), .B2(G168), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n846), .B2(new_n847), .ZN(new_n949));
  INV_X1    g524(.A(new_n947), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(G301), .B2(G286), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n896), .A2(new_n898), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n952), .A3(new_n912), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n949), .A2(new_n952), .A3(KEYINPUT104), .A4(new_n912), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n949), .A2(new_n952), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n905), .A2(KEYINPUT103), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(new_n903), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n955), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n931), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n949), .A2(new_n952), .A3(new_n912), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n909), .B1(new_n949), .B2(new_n952), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n965), .B2(new_n930), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n962), .A2(new_n966), .A3(KEYINPUT105), .A4(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n953), .A2(new_n954), .B1(new_n957), .B2(new_n959), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n930), .B1(new_n970), .B2(new_n956), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n906), .A2(new_n908), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n846), .A2(new_n847), .A3(new_n948), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n951), .B1(new_n896), .B2(new_n898), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n930), .A3(new_n953), .ZN(new_n976));
  INV_X1    g551(.A(G37), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n967), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n969), .B1(new_n971), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n965), .A2(new_n930), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n976), .A2(new_n977), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n968), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT106), .B1(new_n971), .B2(new_n981), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n962), .A2(new_n966), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n988), .A3(KEYINPUT43), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n978), .A2(new_n980), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(new_n984), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n985), .A2(new_n992), .ZN(G397));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n875), .B2(G1384), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n872), .A2(KEYINPUT107), .A3(new_n997), .A4(new_n873), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n480), .A2(new_n481), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G2105), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n465), .A2(new_n471), .B1(G101), .B2(new_n474), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(G40), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n750), .B(G2067), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT109), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n715), .A2(new_n718), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n715), .A2(new_n718), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1004), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n767), .B(G1996), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1004), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1986), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n587), .B(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1013), .B1(new_n1004), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT112), .B(G8), .Z(new_n1017));
  NOR2_X1   g592(.A1(G168), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n497), .B2(new_n500), .ZN(new_n1022));
  INV_X1    g597(.A(new_n996), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1003), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1024), .B(new_n1025), .C1(KEYINPUT45), .C2(new_n1022), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n742), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n501), .A2(new_n997), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1022), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT114), .B(G2084), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1029), .A2(new_n1025), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1017), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT123), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1038), .A3(new_n1035), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1021), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1033), .ZN(new_n1041));
  INV_X1    g616(.A(new_n742), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1003), .B1(new_n1028), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1042), .B1(new_n1044), .B2(new_n1024), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT121), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1027), .A2(new_n1047), .A3(new_n1033), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT122), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1046), .A2(new_n1048), .A3(new_n1051), .A4(G8), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1019), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1040), .B1(new_n1053), .B2(KEYINPUT51), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1046), .A2(new_n1018), .A3(new_n1048), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT62), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1018), .B1(new_n1049), .B2(KEYINPUT122), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1020), .B1(new_n1059), .B2(new_n1052), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1058), .B(new_n1055), .C1(new_n1060), .C2(new_n1040), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1035), .B1(new_n1028), .B2(new_n1003), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  OAI21_X1  g639(.A(G1981), .B1(new_n575), .B2(new_n578), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n575), .A2(new_n578), .A3(G1981), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1067), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT49), .A3(new_n1065), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1063), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n569), .A2(G1976), .A3(new_n571), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT113), .B(G1976), .Z(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1063), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT52), .B1(new_n1062), .B2(new_n1072), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1071), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G8), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n872), .A2(KEYINPUT45), .A3(new_n997), .A4(new_n873), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1028), .A2(new_n996), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1025), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n694), .ZN(new_n1083));
  OAI211_X1 g658(.A(G160), .B(G40), .C1(new_n1022), .C2(new_n1030), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1031), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT110), .B(G2090), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1079), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT111), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT111), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G303), .A2(G8), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1094), .B1(new_n1097), .B2(new_n1090), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1078), .B1(new_n1089), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n694), .A2(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n1017), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1080), .A2(new_n775), .A3(new_n1025), .A4(new_n1081), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1029), .A2(new_n1025), .A3(new_n1031), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1105), .A2(new_n1106), .B1(new_n789), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n775), .A2(KEYINPUT53), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1044), .A2(new_n1024), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n598), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1104), .A2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1057), .A2(new_n1061), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1107), .A2(new_n809), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1025), .A2(new_n1022), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(G2067), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1025), .A2(KEYINPUT118), .A3(new_n755), .A4(new_n1022), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1116), .A2(KEYINPUT60), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n606), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1116), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n596), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1122), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1107), .A2(new_n734), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1080), .A2(new_n1025), .A3(new_n1081), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(KEYINPUT119), .A3(new_n1129), .ZN(new_n1133));
  NAND3_X1  g708(.A1(G299), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n1134));
  NAND2_X1  g709(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1135));
  OR2_X1    g710(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n561), .A2(new_n563), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1132), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1138), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1141), .A2(KEYINPUT61), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1996), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1080), .A2(new_n1144), .A3(new_n1025), .A4(new_n1081), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  NAND3_X1  g721(.A1(new_n1118), .A2(KEYINPUT120), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1146), .B1(new_n1028), .B2(new_n1003), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1145), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n551), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1154), .A3(new_n551), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1141), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1140), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1126), .A2(new_n1143), .A3(new_n1156), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1139), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1123), .A2(new_n606), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1141), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1108), .A2(G301), .A3(new_n1111), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT54), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n999), .A2(new_n1025), .A3(new_n1110), .A4(new_n1080), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n565), .B1(new_n1168), .B2(new_n1108), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(G301), .A3(new_n1108), .ZN(new_n1171));
  AOI21_X1  g746(.A(KEYINPUT54), .B1(new_n1113), .B2(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1170), .A2(new_n1172), .A3(new_n1104), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1165), .B(new_n1173), .C1(new_n1056), .C2(new_n1054), .ZN(new_n1174));
  NOR2_X1   g749(.A1(G288), .A2(G1976), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1071), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1063), .B1(new_n1176), .B2(new_n1067), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1089), .A2(new_n1099), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n1078), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1036), .A2(new_n1180), .A3(G286), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1101), .B1(new_n1089), .B2(KEYINPUT115), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT115), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1102), .A2(new_n1183), .A3(new_n1079), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1100), .B(new_n1181), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT116), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1078), .ZN(new_n1187));
  AOI211_X1 g762(.A(G286), .B(new_n1017), .C1(new_n1027), .C2(new_n1033), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1178), .A2(new_n1103), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1185), .A2(new_n1186), .B1(new_n1180), .B2(new_n1189), .ZN(new_n1190));
  OR2_X1    g765(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1191), .A2(KEYINPUT116), .A3(new_n1100), .A4(new_n1181), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1179), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1174), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1016), .B1(new_n1115), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1004), .B1(new_n767), .B2(new_n1005), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT126), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT47), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1004), .A2(new_n1144), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT46), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1198), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1004), .A2(new_n1014), .A3(new_n587), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1203), .B(KEYINPUT48), .Z(new_n1204));
  OAI22_X1  g779(.A1(new_n1201), .A2(new_n1202), .B1(new_n1013), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1007), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n867), .A2(new_n755), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1206), .B1(new_n1209), .B2(new_n1004), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1004), .ZN(new_n1211));
  AOI211_X1 g786(.A(KEYINPUT125), .B(new_n1211), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1205), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1195), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g789(.A1(new_n886), .A2(new_n890), .ZN(new_n1216));
  NOR3_X1   g790(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1217));
  OAI21_X1  g791(.A(new_n1217), .B1(new_n681), .B2(new_n682), .ZN(new_n1218));
  XNOR2_X1  g792(.A(new_n1218), .B(KEYINPUT127), .ZN(new_n1219));
  AND3_X1   g793(.A1(new_n983), .A2(new_n1216), .A3(new_n1219), .ZN(G308));
  NAND3_X1  g794(.A1(new_n983), .A2(new_n1216), .A3(new_n1219), .ZN(G225));
endmodule


