//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT23), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n193), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n195), .A2(KEYINPUT77), .A3(new_n197), .A4(new_n199), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(G110), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n202), .A2(KEYINPUT78), .A3(G110), .A4(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(G125), .ZN(new_n212));
  INV_X1    g026(.A(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n211), .B1(new_n215), .B2(new_n209), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(G146), .B(new_n211), .C1(new_n215), .C2(new_n209), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT24), .B(G110), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(KEYINPUT75), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n197), .A2(KEYINPUT74), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n197), .A2(KEYINPUT74), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n192), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n220), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n208), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n225), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(G110), .B2(new_n200), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n212), .A2(new_n214), .A3(new_n217), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n219), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT22), .B(G137), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n233), .B(new_n235), .Z(new_n236));
  NAND3_X1  g050(.A1(new_n228), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n236), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n226), .B1(new_n206), .B2(new_n207), .ZN(new_n239));
  INV_X1    g053(.A(new_n232), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n241), .A3(new_n188), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n237), .A2(new_n241), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n190), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n237), .A2(new_n241), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n189), .A2(G902), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G116), .B(G119), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT2), .B(G113), .Z(new_n252));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n252), .A2(KEYINPUT68), .A3(new_n251), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n196), .A2(G116), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G119), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n259), .B1(new_n263), .B2(new_n255), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n267));
  INV_X1    g081(.A(G131), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT65), .B1(new_n269), .B2(G134), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(G134), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(KEYINPUT65), .A3(G134), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G137), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n268), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT64), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n275), .B2(G137), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT11), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n278), .B(KEYINPUT11), .C1(new_n275), .C2(G137), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n277), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n267), .B1(new_n274), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n217), .A2(G143), .ZN(new_n285));
  INV_X1    g099(.A(G143), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G146), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT1), .B1(new_n286), .B2(G146), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(G128), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n285), .B(new_n287), .C1(KEYINPUT1), .C2(new_n191), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n277), .ZN(new_n293));
  INV_X1    g107(.A(new_n282), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n269), .A2(G134), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT11), .B1(new_n295), .B2(new_n278), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n293), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(new_n275), .B2(G137), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n276), .A3(new_n273), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G131), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(KEYINPUT66), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n284), .A2(new_n292), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n271), .B1(new_n281), .B2(new_n282), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n297), .B1(new_n305), .B2(new_n268), .ZN(new_n306));
  AND2_X1   g120(.A1(KEYINPUT0), .A2(G128), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n285), .A2(new_n287), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G143), .B(G146), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT0), .B(G128), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n303), .A2(new_n304), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT69), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n308), .B(new_n315), .C1(new_n309), .C2(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(KEYINPUT69), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n306), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n292), .A2(new_n297), .A3(new_n301), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n304), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n266), .B1(new_n314), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT31), .ZN(new_n322));
  NOR2_X1   g136(.A1(G237), .A2(G953), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G210), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT27), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G101), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n256), .A2(new_n254), .B1(new_n258), .B2(new_n264), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n317), .A2(new_n316), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n276), .B1(new_n294), .B2(new_n296), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n283), .B1(new_n330), .B2(G131), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n319), .B(new_n328), .C1(new_n329), .C2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n321), .A2(new_n322), .A3(new_n327), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT70), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n321), .A2(new_n327), .A3(new_n332), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT31), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n339));
  INV_X1    g153(.A(new_n327), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT71), .ZN(new_n341));
  INV_X1    g155(.A(new_n332), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n328), .B1(new_n303), .B2(new_n313), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n341), .B(KEYINPUT28), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n342), .A2(KEYINPUT28), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n290), .A2(new_n291), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n297), .A2(new_n301), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(new_n267), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n349), .A2(new_n302), .B1(new_n306), .B2(new_n312), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n332), .B1(new_n350), .B2(new_n328), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n341), .B1(new_n351), .B2(KEYINPUT28), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n339), .B(new_n340), .C1(new_n346), .C2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT28), .B1(new_n342), .B2(new_n343), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT71), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n345), .A3(new_n344), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n339), .B1(new_n357), .B2(new_n340), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n337), .B(new_n338), .C1(new_n354), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G472), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n188), .A3(KEYINPUT73), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(G472), .B2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT32), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n364), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n366), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n342), .A2(KEYINPUT28), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n318), .A2(new_n319), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n266), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n332), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(KEYINPUT28), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT29), .A3(new_n327), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n321), .A2(new_n340), .A3(new_n332), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n357), .B2(new_n327), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n188), .B(new_n375), .C1(new_n377), .C2(KEYINPUT29), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n359), .A2(new_n369), .B1(new_n378), .B2(G472), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n250), .B1(new_n367), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n382));
  OAI211_X1 g196(.A(G104), .B(new_n381), .C1(new_n382), .C2(KEYINPUT80), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT81), .A3(G107), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n381), .B2(G104), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n382), .A2(KEYINPUT80), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n390), .A2(new_n391), .B1(G104), .B2(new_n381), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n388), .A2(new_n392), .A3(G101), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT84), .B1(new_n384), .B2(G107), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n381), .A3(G104), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n384), .A2(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G101), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(new_n292), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n384), .A2(G107), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n403), .A2(new_n390), .B1(new_n397), .B2(new_n386), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n381), .A2(G104), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n382), .A2(KEYINPUT80), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G101), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n404), .A2(new_n408), .A3(new_n409), .A4(new_n385), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n399), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n347), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n306), .B1(new_n402), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT12), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(KEYINPUT85), .A2(KEYINPUT10), .ZN(new_n416));
  NAND2_X1  g230(.A1(KEYINPUT85), .A2(KEYINPUT10), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(KEYINPUT85), .B(KEYINPUT10), .C1(new_n411), .C2(new_n347), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G101), .B1(new_n388), .B2(new_n392), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n410), .A2(new_n421), .A3(KEYINPUT4), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT82), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT82), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n410), .A2(new_n421), .A3(new_n424), .A4(KEYINPUT4), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n427), .B(G101), .C1(new_n388), .C2(new_n392), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n317), .A3(new_n316), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT83), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n432), .B(new_n429), .C1(new_n423), .C2(new_n425), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n420), .B(new_n331), .C1(new_n431), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n415), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n234), .A2(G227), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT79), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n439), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n434), .A2(KEYINPUT86), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n420), .B1(new_n431), .B2(new_n433), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n306), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT86), .B1(new_n434), .B2(new_n441), .ZN(new_n446));
  OAI211_X1 g260(.A(G469), .B(new_n440), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G469), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n441), .B1(new_n444), .B2(new_n434), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n415), .A2(new_n434), .A3(new_n441), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n448), .B(new_n188), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(G469), .A2(G902), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G221), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT9), .B(G234), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n456), .B2(new_n188), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G214), .B1(G237), .B2(G902), .ZN(new_n460));
  INV_X1    g274(.A(G237), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n234), .A3(G214), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n463), .A3(new_n286), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n323), .B(G214), .C1(KEYINPUT94), .C2(G143), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT18), .A2(G131), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT95), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n215), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT95), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(G146), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT96), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n472), .A2(new_n473), .A3(new_n231), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n472), .B2(new_n231), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(G113), .B(G122), .Z(new_n477));
  XOR2_X1   g291(.A(KEYINPUT97), .B(G104), .Z(new_n478));
  XOR2_X1   g292(.A(new_n477), .B(new_n478), .Z(new_n479));
  NOR2_X1   g293(.A1(new_n466), .A2(G131), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n268), .B1(new_n464), .B2(new_n465), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n480), .A2(KEYINPUT17), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(KEYINPUT17), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n219), .A3(new_n218), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n476), .B(new_n479), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n470), .A2(KEYINPUT19), .A3(new_n471), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n215), .A2(KEYINPUT19), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(new_n217), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(new_n219), .C1(new_n481), .C2(new_n480), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n476), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n485), .B1(new_n491), .B2(new_n479), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n493));
  NOR2_X1   g307(.A1(G475), .A2(G902), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n492), .B2(new_n494), .ZN(new_n497));
  INV_X1    g311(.A(G475), .ZN(new_n498));
  INV_X1    g312(.A(new_n479), .ZN(new_n499));
  INV_X1    g313(.A(new_n476), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n482), .A2(new_n484), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n502), .B2(new_n485), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(KEYINPUT98), .A2(G122), .ZN(new_n505));
  NOR2_X1   g319(.A1(KEYINPUT98), .A2(G122), .ZN(new_n506));
  OAI21_X1  g320(.A(G116), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n261), .A2(G122), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n381), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(KEYINPUT14), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n286), .A2(G128), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n191), .A2(G143), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n275), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT100), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(new_n513), .A3(new_n275), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n517), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT100), .B1(new_n519), .B2(new_n514), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n507), .B(new_n508), .C1(KEYINPUT14), .C2(new_n381), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n511), .A2(new_n518), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n286), .A2(KEYINPUT13), .A3(G128), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n513), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT13), .B1(new_n286), .B2(G128), .ZN(new_n525));
  OAI21_X1  g339(.A(G134), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT99), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n507), .A2(new_n381), .A3(new_n508), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n517), .B1(new_n529), .B2(new_n509), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n522), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n455), .A2(new_n187), .A3(G953), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n522), .B(new_n532), .C1(new_n528), .C2(new_n530), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT101), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT101), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(new_n537), .A3(new_n533), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n188), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT102), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT102), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n536), .A2(new_n541), .A3(new_n188), .A4(new_n538), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT15), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n540), .A2(new_n542), .B1(new_n543), .B2(G478), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n542), .A2(new_n543), .A3(G478), .ZN(new_n545));
  INV_X1    g359(.A(G952), .ZN(new_n546));
  AOI211_X1 g360(.A(G953), .B(new_n546), .C1(G234), .C2(G237), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n188), .B(new_n234), .C1(G234), .C2(G237), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT21), .B(G898), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR4_X1   g364(.A1(new_n504), .A2(new_n544), .A3(new_n545), .A4(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G122), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G110), .ZN(new_n553));
  INV_X1    g367(.A(G110), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(G122), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT87), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n553), .B2(new_n555), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n266), .A2(new_n428), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n425), .B2(new_n423), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n563));
  INV_X1    g377(.A(G113), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n260), .A2(new_n262), .A3(KEYINPUT5), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n401), .A2(new_n265), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n560), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n428), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n328), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n388), .A2(new_n392), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n427), .B1(new_n573), .B2(new_n409), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n424), .B1(new_n574), .B2(new_n421), .ZN(new_n575));
  INV_X1    g389(.A(new_n425), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n560), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n568), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n570), .A2(new_n579), .A3(KEYINPUT6), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT6), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n581), .B(new_n560), .C1(new_n562), .C2(new_n569), .ZN(new_n582));
  AOI21_X1  g396(.A(G125), .B1(new_n290), .B2(new_n291), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT88), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n583), .A2(new_n584), .B1(G125), .B2(new_n311), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT88), .B1(new_n292), .B2(G125), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G224), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G953), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n587), .B(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(new_n582), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT8), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n553), .A2(new_n555), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT87), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT89), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n557), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n595), .B1(new_n594), .B2(new_n557), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n592), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n265), .B(new_n567), .C1(new_n393), .C2(new_n400), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT89), .B1(new_n558), .B2(new_n559), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n596), .A3(KEYINPUT8), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT90), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n251), .A2(new_n605), .A3(KEYINPUT5), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n565), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n265), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT91), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n265), .A2(new_n607), .A3(KEYINPUT91), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n401), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT7), .B1(new_n588), .B2(G953), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n347), .A2(new_n584), .A3(new_n213), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n311), .A2(G125), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n583), .A2(new_n584), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n585), .A2(new_n586), .A3(new_n613), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n603), .A2(new_n612), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n579), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT92), .B1(new_n622), .B2(new_n188), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT92), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n624), .B(G902), .C1(new_n621), .C2(new_n579), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n591), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(G210), .B1(G237), .B2(G902), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n627), .B(new_n591), .C1(new_n623), .C2(new_n625), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(KEYINPUT93), .A3(new_n630), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n630), .A2(KEYINPUT93), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n460), .A2(new_n551), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n380), .A2(new_n459), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G101), .ZN(G3));
  NAND2_X1  g449(.A1(new_n359), .A2(new_n188), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n337), .A2(new_n338), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n340), .B1(new_n346), .B2(new_n352), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT72), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n353), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n368), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n360), .B1(new_n359), .B2(new_n188), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(KEYINPUT103), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n453), .A2(new_n458), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n250), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n562), .A2(new_n569), .A3(new_n560), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n610), .A2(new_n401), .A3(new_n611), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n617), .A2(new_n618), .A3(new_n614), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n613), .B1(new_n585), .B2(new_n586), .ZN(new_n655));
  OAI22_X1  g469(.A1(new_n652), .A2(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n188), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n624), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n622), .A2(KEYINPUT92), .A3(new_n188), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n627), .B1(new_n660), .B2(new_n591), .ZN(new_n661));
  INV_X1    g475(.A(new_n630), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n460), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n550), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT33), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n536), .A2(new_n667), .A3(new_n538), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n534), .A2(KEYINPUT33), .A3(new_n535), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(G478), .A3(new_n188), .A4(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(G478), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n539), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n504), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n629), .A2(new_n630), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(KEYINPUT104), .A3(new_n460), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n665), .A2(new_n666), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n678), .A2(KEYINPUT105), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(KEYINPUT105), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n648), .B(new_n650), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G104), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT106), .B(KEYINPUT34), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G6));
  NAND2_X1  g498(.A1(new_n502), .A2(new_n485), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n498), .B1(new_n685), .B2(new_n188), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n492), .A2(new_n494), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT20), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n688), .B2(new_n495), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n544), .B2(new_n545), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n665), .A2(new_n666), .A3(new_n677), .A4(new_n691), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n647), .A2(new_n692), .A3(new_n250), .A4(new_n649), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT35), .B(G107), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  NAND2_X1  g509(.A1(new_n633), .A2(new_n459), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n228), .A2(new_n232), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n238), .A2(KEYINPUT36), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n248), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n246), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n639), .A2(new_n646), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n696), .B1(new_n703), .B2(KEYINPUT107), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n639), .A2(new_n646), .A3(new_n705), .A4(new_n702), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT37), .B(G110), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT108), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n707), .B(new_n709), .ZN(G12));
  NAND3_X1  g524(.A1(new_n459), .A2(new_n665), .A3(new_n677), .ZN(new_n711));
  INV_X1    g525(.A(G900), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n548), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n547), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n689), .B(new_n715), .C1(new_n544), .C2(new_n545), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n246), .A2(new_n701), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n354), .A2(new_n358), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n337), .A2(new_n338), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n369), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n378), .A2(G472), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT32), .B1(new_n359), .B2(new_n364), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n718), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT109), .B1(new_n711), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n716), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n702), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n367), .B2(new_n379), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT104), .B1(new_n676), .B2(new_n460), .ZN(new_n731));
  INV_X1    g545(.A(new_n460), .ZN(new_n732));
  AOI211_X1 g546(.A(new_n664), .B(new_n732), .C1(new_n629), .C2(new_n630), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n729), .A2(new_n730), .A3(new_n459), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n726), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT110), .B(G128), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G30));
  AND2_X1   g552(.A1(new_n321), .A2(new_n332), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n739), .A2(new_n340), .ZN(new_n740));
  INV_X1    g554(.A(new_n373), .ZN(new_n741));
  AOI21_X1  g555(.A(G902), .B1(new_n741), .B2(new_n340), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n360), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n359), .B2(new_n369), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n367), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n544), .A2(new_n545), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n504), .ZN(new_n747));
  NOR4_X1   g561(.A1(new_n745), .A2(new_n732), .A3(new_n702), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n715), .B(KEYINPUT39), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n459), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT40), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n631), .A2(new_n632), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT38), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n748), .A2(new_n752), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G143), .ZN(G45));
  INV_X1    g572(.A(new_n715), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n674), .A2(new_n759), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n459), .A2(new_n665), .A3(new_n677), .A4(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n717), .B1(new_n367), .B2(new_n379), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G146), .ZN(G48));
  OAI21_X1  g578(.A(new_n188), .B1(new_n449), .B2(new_n450), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(G469), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n766), .A2(new_n458), .A3(new_n451), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n249), .B(new_n767), .C1(new_n723), .C2(new_n724), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n678), .A2(KEYINPUT105), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n734), .A2(new_n770), .A3(new_n666), .A4(new_n675), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT41), .B(G113), .Z(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G15));
  NOR3_X1   g588(.A1(new_n731), .A2(new_n733), .A3(new_n550), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(new_n380), .A3(new_n691), .A4(new_n767), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G116), .ZN(G18));
  NAND3_X1  g591(.A1(new_n766), .A2(new_n458), .A3(new_n451), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n731), .A2(new_n733), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n762), .A3(new_n551), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G119), .ZN(G21));
  INV_X1    g595(.A(new_n747), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n665), .A2(new_n666), .A3(new_n677), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n364), .B(KEYINPUT111), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n336), .B1(new_n327), .B2(new_n374), .ZN(new_n785));
  INV_X1    g599(.A(new_n333), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n637), .A2(new_n767), .A3(new_n249), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n552), .ZN(G24));
  NAND4_X1  g604(.A1(new_n637), .A2(new_n702), .A3(new_n760), .A4(new_n787), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n665), .A2(new_n767), .A3(new_n677), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n213), .ZN(G27));
  INV_X1    g608(.A(KEYINPUT42), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n721), .B(new_n722), .C1(new_n644), .C2(KEYINPUT32), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n732), .B1(new_n631), .B2(new_n632), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n249), .A3(new_n459), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n760), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n754), .A2(new_n458), .A3(new_n453), .A4(new_n460), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT42), .A3(new_n380), .A4(new_n760), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G131), .ZN(G33));
  OAI21_X1  g619(.A(new_n249), .B1(new_n723), .B2(new_n724), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n806), .A2(new_n801), .A3(new_n716), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(new_n275), .ZN(G36));
  AND2_X1   g622(.A1(new_n689), .A2(new_n673), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT43), .B1(new_n689), .B2(KEYINPUT113), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n809), .B(new_n810), .Z(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n702), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT44), .B1(new_n812), .B2(new_n647), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n440), .B1(new_n445), .B2(new_n446), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(G469), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n452), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT46), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n451), .A2(new_n452), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT46), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n457), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n749), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT112), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n827), .A3(new_n749), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n813), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n812), .A2(KEYINPUT44), .A3(new_n647), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n797), .B1(new_n830), .B2(new_n831), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT115), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n830), .A2(new_n831), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n797), .A4(new_n832), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n829), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G137), .ZN(G39));
  INV_X1    g654(.A(KEYINPUT47), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT116), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT116), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n824), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n820), .A2(new_n823), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(KEYINPUT116), .A3(new_n841), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n796), .A2(new_n249), .A3(new_n799), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n797), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G140), .ZN(G42));
  AND2_X1   g664(.A1(new_n745), .A2(new_n249), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n766), .A2(new_n451), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n852), .A2(KEYINPUT49), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(KEYINPUT49), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n809), .A2(new_n458), .A3(new_n460), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n851), .A2(new_n755), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  INV_X1    g672(.A(new_n793), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n731), .A2(new_n733), .A3(new_n747), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n715), .B(KEYINPUT117), .Z(new_n861));
  NOR3_X1   g675(.A1(new_n246), .A2(new_n701), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n453), .A2(new_n458), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n367), .B2(new_n744), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n761), .A2(new_n762), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(KEYINPUT52), .A2(new_n736), .A3(new_n859), .A4(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n793), .B1(new_n726), .B2(new_n735), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT52), .B1(new_n867), .B2(new_n865), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(G902), .B1(new_n640), .B2(new_n643), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n249), .B(new_n787), .C1(new_n870), .C2(new_n360), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n860), .A2(new_n666), .A3(new_n872), .A4(new_n767), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n776), .A2(new_n873), .A3(new_n780), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n772), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n631), .A2(new_n460), .A3(new_n632), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n690), .A2(new_n674), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n666), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n639), .A2(new_n879), .A3(new_n646), .A4(new_n650), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n634), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n706), .B2(new_n704), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n746), .A2(new_n504), .A3(new_n759), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n702), .B(new_n883), .C1(new_n723), .C2(new_n724), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n801), .B1(new_n884), .B2(new_n791), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n807), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n875), .A2(new_n882), .A3(new_n804), .A4(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n858), .B1(new_n869), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n551), .B(new_n702), .C1(new_n723), .C2(new_n724), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n692), .A2(new_n768), .B1(new_n889), .B2(new_n792), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n789), .ZN(new_n891));
  INV_X1    g705(.A(new_n768), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n679), .B2(new_n680), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n891), .A2(new_n893), .A3(new_n804), .A4(new_n886), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n707), .A2(new_n634), .A3(new_n880), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n736), .A2(new_n865), .A3(new_n859), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT52), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n867), .A2(KEYINPUT52), .A3(new_n865), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n896), .A2(new_n901), .A3(KEYINPUT53), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n888), .A2(KEYINPUT54), .A3(new_n902), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n811), .A2(new_n547), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n732), .A3(new_n755), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n788), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT50), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n908), .A2(new_n872), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n852), .A2(new_n458), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n797), .B(new_n912), .C1(new_n847), .C2(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n797), .A2(new_n767), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n851), .A2(new_n547), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n504), .A2(new_n673), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n908), .A2(new_n915), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n637), .A2(new_n702), .A3(new_n787), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n911), .A2(new_n914), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT51), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n912), .A2(new_n779), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT118), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n918), .A2(new_n380), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT48), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n546), .B(G953), .C1(new_n916), .C2(new_n675), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n923), .A2(new_n924), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n907), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(G952), .A2(G953), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n857), .B1(new_n932), .B2(new_n933), .ZN(G75));
  NOR2_X1   g748(.A1(new_n234), .A2(G952), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n188), .B1(new_n888), .B2(new_n902), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT56), .B1(new_n937), .B2(G210), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n580), .A2(new_n582), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n590), .ZN(new_n940));
  XOR2_X1   g754(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n936), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n903), .B2(G902), .ZN(new_n945));
  AOI211_X1 g759(.A(KEYINPUT120), .B(new_n188), .C1(new_n888), .C2(new_n902), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n628), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n943), .B1(new_n948), .B2(new_n950), .ZN(G51));
  INV_X1    g765(.A(new_n818), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n452), .B(KEYINPUT57), .Z(new_n954));
  NAND3_X1  g768(.A1(new_n905), .A2(new_n906), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n449), .A2(new_n450), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT121), .Z(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n935), .B1(new_n953), .B2(new_n958), .ZN(G54));
  AND2_X1   g773(.A1(KEYINPUT58), .A2(G475), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n492), .B1(new_n947), .B2(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n869), .A2(new_n887), .A3(new_n858), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT53), .B1(new_n896), .B2(new_n901), .ZN(new_n963));
  OAI21_X1  g777(.A(G902), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT120), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n937), .A2(new_n944), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n492), .A2(new_n960), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n936), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n961), .A2(new_n969), .ZN(G60));
  AND2_X1   g784(.A1(new_n668), .A2(new_n669), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n671), .A2(new_n188), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n971), .B1(new_n907), .B2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n905), .A2(new_n971), .A3(new_n906), .A4(new_n974), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n936), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n975), .A2(new_n977), .ZN(G63));
  NAND2_X1  g792(.A1(G217), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT60), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n903), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n247), .B(KEYINPUT123), .Z(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT124), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n980), .B1(new_n888), .B2(new_n902), .ZN(new_n986));
  INV_X1    g800(.A(new_n699), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n935), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT124), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n982), .A2(new_n989), .A3(new_n983), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n985), .A2(KEYINPUT61), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n984), .A2(new_n988), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT61), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n991), .A2(new_n994), .ZN(G66));
  OAI21_X1  g809(.A(G953), .B1(new_n549), .B2(new_n588), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n875), .A2(new_n882), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n996), .B1(new_n998), .B2(G953), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n939), .B1(G898), .B2(new_n234), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(G69));
  NOR2_X1   g815(.A1(new_n314), .A2(new_n320), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n486), .A2(new_n488), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1002), .B(new_n1003), .Z(new_n1004));
  NAND2_X1  g818(.A1(G900), .A2(G953), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n826), .A2(new_n828), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n380), .A3(new_n860), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n867), .A2(new_n763), .ZN(new_n1008));
  INV_X1    g822(.A(new_n807), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1008), .A2(new_n804), .A3(new_n1009), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n839), .A2(new_n849), .A3(new_n1007), .A4(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1004), .B(new_n1005), .C1(new_n1011), .C2(G953), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1008), .A2(new_n757), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1008), .A2(KEYINPUT62), .A3(new_n757), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n877), .B(KEYINPUT125), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n750), .A2(new_n380), .A3(new_n797), .A4(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT126), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n849), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1017), .A2(new_n839), .A3(new_n1021), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1022), .A2(new_n234), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1012), .B1(new_n1023), .B2(new_n1004), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n234), .B1(G227), .B2(G900), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1025), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1012), .B(new_n1027), .C1(new_n1023), .C2(new_n1004), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1026), .A2(new_n1028), .ZN(G72));
  NAND4_X1  g843(.A1(new_n1017), .A2(new_n839), .A3(new_n998), .A4(new_n1021), .ZN(new_n1030));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  NAND2_X1  g846(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n740), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n935), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1032), .B1(new_n1011), .B2(new_n997), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n376), .ZN(new_n1037));
  INV_X1    g851(.A(new_n376), .ZN(new_n1038));
  AND3_X1   g852(.A1(new_n740), .A2(new_n1038), .A3(new_n1032), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n903), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1040), .A2(KEYINPUT127), .ZN(new_n1041));
  AND2_X1   g855(.A1(new_n1040), .A2(KEYINPUT127), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1035), .B(new_n1037), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(G57));
endmodule


