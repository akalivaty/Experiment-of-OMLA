

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582;

  INV_X1 U319 ( .A(KEYINPUT93), .ZN(n392) );
  INV_X1 U320 ( .A(KEYINPUT32), .ZN(n329) );
  XNOR2_X1 U321 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U322 ( .A(n381), .B(n331), .ZN(n335) );
  INV_X1 U323 ( .A(n395), .ZN(n397) );
  XNOR2_X1 U324 ( .A(n515), .B(KEYINPUT27), .ZN(n395) );
  XNOR2_X1 U325 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U326 ( .A(KEYINPUT48), .B(KEYINPUT111), .ZN(n462) );
  XNOR2_X1 U327 ( .A(KEYINPUT37), .B(KEYINPUT99), .ZN(n441) );
  XNOR2_X1 U328 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U329 ( .A(n463), .B(n462), .ZN(n541) );
  XNOR2_X1 U330 ( .A(n442), .B(n441), .ZN(n511) );
  XNOR2_X1 U331 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U332 ( .A(n377), .B(n376), .ZN(n464) );
  INV_X1 U333 ( .A(G43GAT), .ZN(n445) );
  XNOR2_X1 U334 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U335 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U336 ( .A(n477), .B(n476), .ZN(G1349GAT) );
  XNOR2_X1 U337 ( .A(n448), .B(n447), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(G176GAT), .B(KEYINPUT86), .Z(n288) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(G99GAT), .ZN(n287) );
  XNOR2_X1 U340 ( .A(n288), .B(n287), .ZN(n289) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G71GAT), .Z(n339) );
  XOR2_X1 U342 ( .A(n289), .B(n339), .Z(n291) );
  XNOR2_X1 U343 ( .A(G169GAT), .B(G15GAT), .ZN(n290) );
  XNOR2_X1 U344 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U345 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n293) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U347 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U348 ( .A(n295), .B(n294), .Z(n301) );
  XNOR2_X1 U349 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n296), .B(KEYINPUT19), .ZN(n297) );
  XOR2_X1 U351 ( .A(n297), .B(KEYINPUT17), .Z(n299) );
  XNOR2_X1 U352 ( .A(G183GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n375) );
  XNOR2_X1 U354 ( .A(n375), .B(KEYINPUT83), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U356 ( .A(KEYINPUT82), .B(G134GAT), .Z(n303) );
  XNOR2_X1 U357 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U359 ( .A(G113GAT), .B(n304), .Z(n353) );
  XOR2_X1 U360 ( .A(n305), .B(n353), .Z(n524) );
  INV_X1 U361 ( .A(n524), .ZN(n517) );
  XOR2_X1 U362 ( .A(G43GAT), .B(G29GAT), .Z(n307) );
  XNOR2_X1 U363 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U365 ( .A(n308), .B(KEYINPUT8), .Z(n310) );
  XNOR2_X1 U366 ( .A(G36GAT), .B(KEYINPUT70), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n437) );
  XOR2_X1 U368 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n312) );
  XNOR2_X1 U369 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n437), .B(n313), .ZN(n322) );
  XOR2_X1 U372 ( .A(G141GAT), .B(G22GAT), .Z(n386) );
  XOR2_X1 U373 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n315) );
  XNOR2_X1 U374 ( .A(G15GAT), .B(G1GAT), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n315), .B(n314), .ZN(n415) );
  XOR2_X1 U376 ( .A(n386), .B(n415), .Z(n317) );
  NAND2_X1 U377 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U379 ( .A(G169GAT), .B(G8GAT), .Z(n373) );
  XOR2_X1 U380 ( .A(n318), .B(n373), .Z(n320) );
  XNOR2_X1 U381 ( .A(G113GAT), .B(G197GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n566) );
  XNOR2_X1 U384 ( .A(n566), .B(KEYINPUT73), .ZN(n556) );
  INV_X1 U385 ( .A(G148GAT), .ZN(n323) );
  NAND2_X1 U386 ( .A1(G78GAT), .A2(n323), .ZN(n326) );
  INV_X1 U387 ( .A(G78GAT), .ZN(n324) );
  NAND2_X1 U388 ( .A1(n324), .A2(G148GAT), .ZN(n325) );
  NAND2_X1 U389 ( .A1(n326), .A2(n325), .ZN(n328) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n328), .B(n327), .ZN(n381) );
  NAND2_X1 U392 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  XOR2_X1 U393 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n333) );
  XNOR2_X1 U394 ( .A(KEYINPUT31), .B(KEYINPUT77), .ZN(n332) );
  XOR2_X1 U395 ( .A(n333), .B(n332), .Z(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n342) );
  XOR2_X1 U397 ( .A(G64GAT), .B(G92GAT), .Z(n337) );
  XNOR2_X1 U398 ( .A(G176GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n369) );
  XNOR2_X1 U400 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n338), .B(KEYINPUT74), .ZN(n414) );
  XNOR2_X1 U402 ( .A(n369), .B(n414), .ZN(n340) );
  XNOR2_X1 U403 ( .A(G99GAT), .B(G85GAT), .ZN(n427) );
  XOR2_X1 U404 ( .A(n343), .B(n427), .Z(n449) );
  NAND2_X1 U405 ( .A1(n556), .A2(n449), .ZN(n344) );
  XOR2_X1 U406 ( .A(KEYINPUT78), .B(n344), .Z(n482) );
  XOR2_X1 U407 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n346) );
  XNOR2_X1 U408 ( .A(KEYINPUT6), .B(KEYINPUT88), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n363) );
  XOR2_X1 U410 ( .A(G85GAT), .B(G148GAT), .Z(n348) );
  XNOR2_X1 U411 ( .A(G29GAT), .B(G120GAT), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U413 ( .A(G57GAT), .B(KEYINPUT4), .Z(n350) );
  XNOR2_X1 U414 ( .A(G141GAT), .B(G1GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U416 ( .A(n352), .B(n351), .Z(n361) );
  INV_X1 U417 ( .A(n353), .ZN(n359) );
  XOR2_X1 U418 ( .A(G155GAT), .B(KEYINPUT3), .Z(n355) );
  XNOR2_X1 U419 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n382) );
  XOR2_X1 U421 ( .A(n382), .B(KEYINPUT87), .Z(n357) );
  NAND2_X1 U422 ( .A1(G225GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U424 ( .A(n359), .B(n358), .Z(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n540) );
  XOR2_X1 U427 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n365) );
  NAND2_X1 U428 ( .A1(G226GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U430 ( .A(n366), .B(KEYINPUT92), .Z(n371) );
  XOR2_X1 U431 ( .A(G211GAT), .B(KEYINPUT21), .Z(n368) );
  XNOR2_X1 U432 ( .A(G197GAT), .B(G218GAT), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n390) );
  XNOR2_X1 U434 ( .A(n369), .B(n390), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U436 ( .A(n372), .B(KEYINPUT91), .Z(n377) );
  XNOR2_X1 U437 ( .A(G36GAT), .B(n373), .ZN(n374) );
  INV_X1 U438 ( .A(n464), .ZN(n515) );
  NOR2_X1 U439 ( .A1(n540), .A2(n395), .ZN(n391) );
  XOR2_X1 U440 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n379) );
  NAND2_X1 U441 ( .A1(G228GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U443 ( .A(n380), .B(KEYINPUT24), .Z(n384) );
  XNOR2_X1 U444 ( .A(n381), .B(n382), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U446 ( .A(n385), .B(G204GAT), .Z(n388) );
  XNOR2_X1 U447 ( .A(G50GAT), .B(n386), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n469) );
  XNOR2_X1 U450 ( .A(KEYINPUT28), .B(n469), .ZN(n520) );
  NAND2_X1 U451 ( .A1(n391), .A2(n520), .ZN(n526) );
  XNOR2_X1 U452 ( .A(n526), .B(n392), .ZN(n393) );
  NOR2_X1 U453 ( .A1(n524), .A2(n393), .ZN(n394) );
  XOR2_X1 U454 ( .A(KEYINPUT94), .B(n394), .Z(n405) );
  NOR2_X1 U455 ( .A1(n469), .A2(n524), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n396), .B(KEYINPUT26), .ZN(n564) );
  NAND2_X1 U457 ( .A1(n397), .A2(n564), .ZN(n539) );
  XOR2_X1 U458 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n401) );
  NAND2_X1 U459 ( .A1(n524), .A2(n464), .ZN(n398) );
  XOR2_X1 U460 ( .A(KEYINPUT95), .B(n398), .Z(n399) );
  NAND2_X1 U461 ( .A1(n399), .A2(n469), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n402) );
  NAND2_X1 U463 ( .A1(n539), .A2(n402), .ZN(n403) );
  NAND2_X1 U464 ( .A1(n403), .A2(n540), .ZN(n404) );
  NAND2_X1 U465 ( .A1(n405), .A2(n404), .ZN(n479) );
  XOR2_X1 U466 ( .A(KEYINPUT81), .B(G64GAT), .Z(n407) );
  XNOR2_X1 U467 ( .A(G8GAT), .B(G22GAT), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n423) );
  XOR2_X1 U469 ( .A(G155GAT), .B(G78GAT), .Z(n409) );
  XNOR2_X1 U470 ( .A(G183GAT), .B(G211GAT), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U472 ( .A(G127GAT), .B(G71GAT), .Z(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n419) );
  XNOR2_X1 U474 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n412), .B(KEYINPUT12), .ZN(n413) );
  XOR2_X1 U476 ( .A(n413), .B(KEYINPUT80), .Z(n417) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n421) );
  NAND2_X1 U480 ( .A1(G231GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U482 ( .A(n423), .B(n422), .Z(n575) );
  NAND2_X1 U483 ( .A1(n479), .A2(n575), .ZN(n440) );
  XOR2_X1 U484 ( .A(G92GAT), .B(G162GAT), .Z(n425) );
  XNOR2_X1 U485 ( .A(G218GAT), .B(G106GAT), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U487 ( .A(n427), .B(n426), .ZN(n429) );
  NAND2_X1 U488 ( .A1(G232GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U490 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n431) );
  XNOR2_X1 U491 ( .A(G190GAT), .B(KEYINPUT11), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n439) );
  XOR2_X1 U494 ( .A(KEYINPUT67), .B(KEYINPUT79), .Z(n435) );
  XNOR2_X1 U495 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n560) );
  XOR2_X1 U499 ( .A(KEYINPUT36), .B(n560), .Z(n579) );
  NOR2_X1 U500 ( .A1(n440), .A2(n579), .ZN(n442) );
  NAND2_X1 U501 ( .A1(n482), .A2(n511), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n443), .B(KEYINPUT38), .ZN(n444) );
  XNOR2_X1 U503 ( .A(KEYINPUT100), .B(n444), .ZN(n495) );
  NOR2_X1 U504 ( .A1(n517), .A2(n495), .ZN(n448) );
  XNOR2_X1 U505 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n446) );
  INV_X1 U506 ( .A(KEYINPUT41), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n473) );
  NOR2_X1 U508 ( .A1(n566), .A2(n473), .ZN(n452) );
  INV_X1 U509 ( .A(KEYINPUT46), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n452), .B(n451), .ZN(n454) );
  INV_X1 U511 ( .A(n560), .ZN(n553) );
  AND2_X1 U512 ( .A1(n575), .A2(n553), .ZN(n453) );
  NAND2_X1 U513 ( .A1(n454), .A2(n453), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n455), .B(KEYINPUT47), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n457) );
  NOR2_X1 U516 ( .A1(n579), .A2(n575), .ZN(n456) );
  XOR2_X1 U517 ( .A(n457), .B(n456), .Z(n458) );
  NAND2_X1 U518 ( .A1(n449), .A2(n458), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n556), .A2(n459), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n461), .A2(n460), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n541), .A2(n464), .ZN(n466) );
  XOR2_X1 U522 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n465) );
  XNOR2_X1 U523 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n467), .A2(n540), .ZN(n468) );
  XOR2_X1 U525 ( .A(KEYINPUT64), .B(n468), .Z(n565) );
  NAND2_X1 U526 ( .A1(n565), .A2(n469), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT55), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n471), .A2(n524), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(KEYINPUT121), .ZN(n561) );
  INV_X1 U530 ( .A(n473), .ZN(n529) );
  NAND2_X1 U531 ( .A1(n561), .A2(n529), .ZN(n477) );
  XOR2_X1 U532 ( .A(G176GAT), .B(KEYINPUT56), .Z(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n575), .A2(n560), .ZN(n478) );
  XNOR2_X1 U535 ( .A(KEYINPUT16), .B(n478), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n481), .B(KEYINPUT97), .ZN(n498) );
  NAND2_X1 U538 ( .A1(n498), .A2(n482), .ZN(n489) );
  NOR2_X1 U539 ( .A1(n540), .A2(n489), .ZN(n484) );
  XNOR2_X1 U540 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U542 ( .A(G1GAT), .B(n485), .Z(G1324GAT) );
  NOR2_X1 U543 ( .A1(n515), .A2(n489), .ZN(n486) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  NOR2_X1 U545 ( .A1(n517), .A2(n489), .ZN(n488) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n520), .A2(n489), .ZN(n490) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n490), .Z(G1327GAT) );
  NOR2_X1 U550 ( .A1(n540), .A2(n495), .ZN(n493) );
  XOR2_X1 U551 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n491) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n491), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U554 ( .A1(n515), .A2(n495), .ZN(n494) );
  XOR2_X1 U555 ( .A(G36GAT), .B(n494), .Z(G1329GAT) );
  NOR2_X1 U556 ( .A1(n520), .A2(n495), .ZN(n496) );
  XOR2_X1 U557 ( .A(G50GAT), .B(n496), .Z(G1331GAT) );
  NAND2_X1 U558 ( .A1(n529), .A2(n566), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT103), .ZN(n512) );
  NAND2_X1 U560 ( .A1(n512), .A2(n498), .ZN(n505) );
  NOR2_X1 U561 ( .A1(n540), .A2(n505), .ZN(n499) );
  XOR2_X1 U562 ( .A(G57GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT42), .B(n500), .ZN(G1332GAT) );
  NOR2_X1 U564 ( .A1(n515), .A2(n505), .ZN(n501) );
  XOR2_X1 U565 ( .A(KEYINPUT104), .B(n501), .Z(n502) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U567 ( .A1(n517), .A2(n505), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(G1334GAT) );
  NOR2_X1 U570 ( .A1(n520), .A2(n505), .ZN(n510) );
  XOR2_X1 U571 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n507) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(KEYINPUT106), .B(n508), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n513) );
  XOR2_X1 U577 ( .A(KEYINPUT109), .B(n513), .Z(n519) );
  NOR2_X1 U578 ( .A1(n540), .A2(n519), .ZN(n514) );
  XOR2_X1 U579 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U580 ( .A1(n515), .A2(n519), .ZN(n516) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n517), .A2(n519), .ZN(n518) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U585 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U587 ( .A(G106GAT), .B(n523), .Z(G1339GAT) );
  NAND2_X1 U588 ( .A1(n524), .A2(n541), .ZN(n525) );
  NOR2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n556), .A2(n535), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(KEYINPUT112), .ZN(n528) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U594 ( .A1(n535), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U596 ( .A(G120GAT), .B(n532), .Z(G1341GAT) );
  INV_X1 U597 ( .A(n575), .ZN(n558) );
  NAND2_X1 U598 ( .A1(n558), .A2(n535), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U602 ( .A1(n535), .A2(n560), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U607 ( .A(KEYINPUT115), .B(n543), .Z(n552) );
  NOR2_X1 U608 ( .A1(n566), .A2(n552), .ZN(n544) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  NOR2_X1 U610 ( .A1(n473), .A2(n552), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT116), .B(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n575), .A2(n552), .ZN(n550) );
  XOR2_X1 U617 ( .A(KEYINPUT118), .B(n550), .Z(n551) );
  XNOR2_X1 U618 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n561), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n561), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n578) );
  NOR2_X1 U630 ( .A1(n578), .A2(n566), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n578), .A2(n449), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(n576), .Z(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

