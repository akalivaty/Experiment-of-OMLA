//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n545, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2106), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n462), .B1(new_n475), .B2(new_n476), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  MUX2_X1   g055(.A(G100), .B(G112), .S(G2105), .Z(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G138), .A4(new_n462), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G102), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2104), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT6), .B(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G50), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n500), .A2(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT66), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n509), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n508), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n500), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n503), .A2(new_n502), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n499), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n509), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT67), .B(G90), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n500), .A2(new_n531), .B1(new_n506), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n530), .A2(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  AOI22_X1  g110(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n509), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n500), .A2(new_n538), .B1(new_n506), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT68), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n543), .A2(new_n547), .ZN(G188));
  NOR3_X1   g123(.A1(new_n503), .A2(new_n502), .A3(KEYINPUT70), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n512), .B2(new_n513), .ZN(new_n551));
  OAI21_X1  g126(.A(G65), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT69), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n554), .A2(KEYINPUT69), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n552), .A2(new_n553), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT70), .B1(new_n503), .B2(new_n502), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n512), .A2(new_n550), .A3(new_n513), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n555), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT71), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(G651), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n500), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n505), .ZN(new_n567));
  NAND2_X1  g142(.A1(KEYINPUT6), .A2(G651), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n511), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n569), .A2(new_n570), .A3(G53), .ZN(new_n571));
  INV_X1    g146(.A(new_n506), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n566), .A2(new_n571), .B1(G91), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n564), .A2(new_n573), .ZN(G299));
  XNOR2_X1  g149(.A(G168), .B(KEYINPUT72), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n572), .A2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n569), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n506), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n514), .A2(new_n499), .A3(KEYINPUT73), .A4(G86), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n524), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G48), .B2(new_n569), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n509), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n500), .A2(new_n594), .B1(new_n506), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  XOR2_X1   g174(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n572), .A2(G92), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n600), .B1(new_n506), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n569), .A2(G54), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(G66), .B1(new_n549), .B2(new_n551), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n509), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(KEYINPUT75), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(KEYINPUT75), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n599), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n599), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(G299), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n617), .B2(new_n575), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(new_n617), .B2(new_n575), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  INV_X1    g197(.A(new_n541), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n611), .A2(new_n621), .A3(new_n612), .ZN(new_n624));
  MUX2_X1   g199(.A(new_n623), .B(new_n624), .S(G868), .Z(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n477), .A2(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(KEYINPUT13), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(KEYINPUT13), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n630), .B(new_n631), .C1(KEYINPUT77), .C2(G2100), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT77), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n630), .A2(KEYINPUT77), .A3(G2100), .A4(new_n631), .ZN(new_n636));
  MUX2_X1   g211(.A(G99), .B(G111), .S(G2105), .Z(new_n637));
  AOI22_X1  g212(.A1(G123), .A2(new_n479), .B1(new_n637), .B2(G2104), .ZN(new_n638));
  INV_X1    g213(.A(G135), .ZN(new_n639));
  INV_X1    g214(.A(new_n477), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n635), .A2(new_n636), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT78), .ZN(G156));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2443), .B(G2446), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n649), .B(KEYINPUT79), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(new_n652), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n647), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT80), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2430), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT14), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n654), .A2(new_n656), .A3(new_n647), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n658), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n666), .ZN(new_n669));
  INV_X1    g244(.A(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(new_n670), .B2(new_n657), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(new_n671), .A3(G14), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g249(.A1(new_n668), .A2(new_n671), .A3(KEYINPUT81), .A4(G14), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT82), .Z(G401));
  XOR2_X1   g252(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n678));
  NOR2_X1   g253(.A1(G2072), .A2(G2078), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n442), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n682), .B(KEYINPUT85), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(new_n680), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2084), .B(G2090), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT83), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n685), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT87), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n690), .A2(new_n681), .A3(new_n684), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n689), .B(new_n682), .C1(new_n442), .C2(new_n679), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n696), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n693), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n692), .A2(new_n642), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n642), .B1(new_n692), .B2(new_n699), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n634), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n702), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(G2100), .A3(new_n700), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(G227));
  XNOR2_X1  g281(.A(G1961), .B(G1966), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT88), .ZN(new_n708));
  XOR2_X1   g283(.A(G1956), .B(G2474), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1971), .B(G1976), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT19), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n708), .A2(new_n709), .ZN(new_n714));
  MUX2_X1   g289(.A(new_n713), .B(new_n712), .S(new_n714), .Z(new_n715));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n708), .A2(KEYINPUT89), .A3(new_n709), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n712), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n716), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI211_X1 g297(.A(KEYINPUT20), .B(new_n712), .C1(new_n718), .C2(new_n719), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n715), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n715), .B(new_n725), .C1(new_n722), .C2(new_n723), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(G1991), .B(G1996), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT90), .ZN(new_n731));
  XOR2_X1   g306(.A(G1981), .B(G1986), .Z(new_n732));
  XOR2_X1   g307(.A(new_n731), .B(new_n732), .Z(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n727), .A2(new_n728), .A3(new_n733), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(G229));
  MUX2_X1   g313(.A(G95), .B(G107), .S(G2105), .Z(new_n739));
  AOI22_X1  g314(.A1(G119), .A2(new_n479), .B1(new_n739), .B2(G2104), .ZN(new_n740));
  INV_X1    g315(.A(G131), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(new_n640), .ZN(new_n742));
  MUX2_X1   g317(.A(G25), .B(new_n742), .S(G29), .Z(new_n743));
  XOR2_X1   g318(.A(KEYINPUT35), .B(G1991), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G16), .A2(G24), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n597), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1986), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G6), .B(G305), .S(G16), .Z(new_n750));
  XOR2_X1   g325(.A(KEYINPUT32), .B(G1981), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G23), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT92), .ZN(new_n754));
  INV_X1    g329(.A(G16), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(G288), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT33), .B(G1976), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G16), .A2(G22), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G166), .B2(G16), .ZN(new_n760));
  INV_X1    g335(.A(G1971), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n752), .A2(new_n758), .A3(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n764));
  OAI211_X1 g339(.A(new_n745), .B(new_n749), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT36), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n470), .A2(G103), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT25), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n487), .A2(G127), .ZN(new_n770));
  INV_X1    g345(.A(G115), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n469), .ZN(new_n772));
  AOI21_X1  g347(.A(KEYINPUT95), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n769), .B(new_n773), .C1(G139), .C2(new_n477), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n772), .A2(KEYINPUT95), .A3(G2105), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G33), .B(new_n776), .S(G29), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2072), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n755), .A2(G19), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT93), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n623), .B2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(G164), .A2(G29), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G27), .B2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT99), .B(G28), .Z(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n787), .B2(KEYINPUT30), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(KEYINPUT30), .B2(new_n787), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT31), .B(G11), .ZN(new_n790));
  INV_X1    g365(.A(G29), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n789), .B(new_n790), .C1(new_n641), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G5), .A2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT101), .Z(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G301), .B2(new_n755), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n792), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n784), .A2(new_n785), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n782), .A2(new_n786), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G104), .B(G116), .S(G2105), .Z(new_n800));
  AOI22_X1  g375(.A1(G128), .A2(new_n479), .B1(new_n800), .B2(G2104), .ZN(new_n801));
  INV_X1    g376(.A(G140), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n640), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G29), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n791), .A2(G26), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT28), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT94), .Z(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(G2067), .ZN(new_n809));
  NAND2_X1  g384(.A1(G160), .A2(G29), .ZN(new_n810));
  AND2_X1   g385(.A1(KEYINPUT24), .A2(G34), .ZN(new_n811));
  NOR2_X1   g386(.A1(KEYINPUT24), .A2(G34), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n791), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G2084), .ZN(new_n815));
  INV_X1    g390(.A(G1966), .ZN(new_n816));
  NOR2_X1   g391(.A1(G168), .A2(new_n755), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n755), .B2(G21), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n815), .B1(new_n796), .B2(new_n795), .C1(new_n816), .C2(new_n818), .ZN(new_n819));
  NOR4_X1   g394(.A1(new_n778), .A2(new_n799), .A3(new_n809), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n816), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT100), .Z(new_n822));
  INV_X1    g397(.A(G2090), .ZN(new_n823));
  NOR2_X1   g398(.A1(G29), .A2(G35), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G162), .B2(G29), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT29), .Z(new_n826));
  AOI22_X1  g401(.A1(new_n808), .A2(G2067), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n822), .B(new_n827), .C1(new_n823), .C2(new_n826), .ZN(new_n828));
  NOR2_X1   g403(.A1(G29), .A2(G32), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n477), .A2(G141), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT96), .Z(new_n831));
  AND2_X1   g406(.A1(new_n470), .A2(G105), .ZN(new_n832));
  NAND3_X1  g407(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT26), .ZN(new_n834));
  AOI211_X1 g409(.A(new_n832), .B(new_n834), .C1(G129), .C2(new_n479), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n829), .B1(new_n838), .B2(G29), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT27), .B(G1996), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT98), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n839), .B(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n828), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n755), .A2(G20), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT102), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT23), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G299), .B2(G16), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G1956), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n755), .A2(G4), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n614), .B2(new_n755), .ZN(new_n850));
  INV_X1    g425(.A(G1348), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  AND4_X1   g427(.A1(new_n820), .A2(new_n843), .A3(new_n848), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n767), .A2(new_n853), .ZN(G150));
  INV_X1    g429(.A(G150), .ZN(G311));
  XNOR2_X1  g430(.A(KEYINPUT105), .B(G860), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n514), .A2(G67), .ZN(new_n857));
  NAND2_X1  g432(.A1(G80), .A2(G543), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n509), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n572), .A2(G93), .B1(G55), .B2(new_n569), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n859), .A2(new_n860), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n859), .A2(new_n860), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n623), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n541), .A3(new_n862), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n613), .A2(new_n621), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n856), .B(new_n874), .C1(new_n875), .C2(KEYINPUT104), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n875), .A2(KEYINPUT104), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n864), .B1(new_n876), .B2(new_n877), .ZN(G145));
  MUX2_X1   g453(.A(G106), .B(G118), .S(G2105), .Z(new_n879));
  AOI22_X1  g454(.A1(G130), .A2(new_n479), .B1(new_n879), .B2(G2104), .ZN(new_n880));
  INV_X1    g455(.A(G142), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n881), .B2(new_n640), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n742), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n629), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n488), .B1(new_n477), .B2(G138), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT106), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n496), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n803), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n883), .B(new_n629), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n836), .B(KEYINPUT107), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n898), .A2(new_n776), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n838), .A2(new_n776), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(G160), .B(new_n483), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(new_n641), .Z(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n894), .B(new_n896), .C1(new_n899), .C2(new_n900), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT108), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n902), .A2(new_n909), .A3(new_n905), .A4(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n902), .A2(new_n906), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n912), .B2(new_n904), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(KEYINPUT40), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT40), .B1(new_n911), .B2(new_n913), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(G395));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  OR2_X1    g494(.A1(new_n606), .A2(new_n609), .ZN(new_n920));
  NAND2_X1  g495(.A1(G299), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n610), .A2(new_n564), .A3(new_n573), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n922), .A3(new_n919), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI211_X1 g501(.A(KEYINPUT109), .B(new_n919), .C1(new_n921), .C2(new_n922), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n624), .B(new_n870), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n918), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G288), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(new_n597), .ZN(new_n932));
  XNOR2_X1  g507(.A(G305), .B(G166), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n932), .B(new_n933), .Z(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT42), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n614), .A2(new_n621), .A3(new_n870), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n624), .A2(new_n868), .A3(new_n869), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n938), .B(KEYINPUT110), .C1(new_n927), .C2(new_n926), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n921), .A2(new_n922), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n929), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n930), .A2(new_n935), .A3(new_n939), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT111), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n930), .A2(new_n939), .A3(new_n942), .ZN(new_n945));
  INV_X1    g520(.A(new_n935), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n943), .A2(KEYINPUT111), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n867), .A2(new_n617), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(G295));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n951), .ZN(G331));
  NAND2_X1  g528(.A1(G301), .A2(G168), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n575), .B2(G301), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(new_n870), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n941), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n957), .B(new_n934), .C1(new_n928), .C2(new_n956), .ZN(new_n958));
  INV_X1    g533(.A(G37), .ZN(new_n959));
  INV_X1    g534(.A(new_n934), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n870), .B(new_n954), .C1(G301), .C2(new_n575), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n868), .A3(new_n869), .ZN(new_n962));
  INV_X1    g537(.A(new_n923), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n961), .A2(new_n962), .B1(new_n963), .B2(new_n925), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n961), .A2(new_n962), .A3(new_n941), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n958), .A2(new_n959), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n957), .B1(new_n928), .B2(new_n956), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n960), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n971), .A2(KEYINPUT43), .A3(new_n959), .A4(new_n958), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT44), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n971), .A2(new_n968), .A3(new_n959), .A4(new_n958), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(KEYINPUT44), .B2(new_n976), .ZN(G397));
  XOR2_X1   g552(.A(KEYINPUT112), .B(G1384), .Z(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT45), .B1(new_n891), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n468), .A2(new_n471), .ZN(new_n981));
  INV_X1    g556(.A(G125), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n475), .B2(new_n476), .ZN(new_n983));
  INV_X1    g558(.A(new_n466), .ZN(new_n984));
  OAI21_X1  g559(.A(G2105), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n985), .A3(G40), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT113), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n988));
  NAND3_X1  g563(.A1(G160), .A2(new_n988), .A3(G40), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n980), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1996), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n838), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n803), .B(G2067), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(G1996), .B2(new_n836), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n991), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT114), .Z(new_n997));
  INV_X1    g572(.A(new_n991), .ZN(new_n998));
  INV_X1    g573(.A(new_n744), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n742), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n742), .A2(new_n999), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n597), .B(new_n748), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n891), .A2(KEYINPUT45), .A3(new_n979), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n490), .B2(new_n496), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1006), .A2(new_n1010), .A3(new_n785), .A4(new_n990), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n494), .A2(new_n495), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n490), .B2(new_n886), .ZN(new_n1015));
  AOI211_X1 g590(.A(KEYINPUT50), .B(G1384), .C1(new_n1015), .C2(new_n890), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n988), .B1(G160), .B2(G40), .ZN(new_n1017));
  AND4_X1   g592(.A1(new_n988), .A2(new_n981), .A3(new_n985), .A4(G40), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n1017), .A2(new_n1018), .B1(new_n1007), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n796), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n987), .A2(new_n989), .B1(new_n1007), .B2(KEYINPUT45), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1012), .A2(G2078), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1384), .B1(new_n1015), .B2(new_n890), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1022), .B(new_n1023), .C1(KEYINPUT45), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G171), .B1(new_n1013), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT123), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(KEYINPUT123), .B(G171), .C1(new_n1013), .C2(new_n1026), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n985), .A2(G40), .A3(new_n1023), .ZN(new_n1033));
  AND4_X1   g608(.A1(new_n1006), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n980), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1034), .A2(new_n1035), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n1021), .A2(KEYINPUT124), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1021), .A2(KEYINPUT124), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1036), .A2(new_n1037), .A3(G301), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1029), .A2(new_n1030), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT55), .B(G8), .C1(new_n508), .C2(new_n518), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1047));
  INV_X1    g622(.A(G1384), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n891), .A2(KEYINPUT50), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1008), .A2(new_n1019), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1006), .A2(new_n990), .A3(new_n1010), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n823), .A2(new_n1051), .B1(new_n1052), .B2(new_n761), .ZN(new_n1053));
  INV_X1    g628(.A(G8), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1046), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n761), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n891), .A2(new_n1019), .A3(new_n1048), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1008), .A2(KEYINPUT50), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n823), .A4(new_n990), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1046), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(G8), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1024), .A2(new_n990), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n931), .A2(G1976), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(G8), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT52), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1054), .B1(new_n1024), .B2(new_n990), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT49), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n569), .A2(G48), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n514), .A2(new_n499), .A3(G86), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1072), .B(new_n1073), .C1(new_n1074), .C2(new_n509), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(G1981), .ZN(new_n1077));
  INV_X1    g652(.A(G1981), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n586), .A2(new_n590), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1076), .B1(new_n1075), .B2(G1981), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1071), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1075), .A2(G1981), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1084), .A2(KEYINPUT49), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(new_n1067), .A3(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1066), .A2(new_n1070), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1055), .A2(new_n1062), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1013), .A2(new_n1026), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1041), .B1(new_n1091), .B2(G301), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1088), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT45), .B1(new_n891), .B2(new_n1048), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n1048), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n816), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G2084), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1057), .A2(new_n1058), .A3(new_n1098), .A4(new_n990), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G8), .ZN(new_n1101));
  OAI21_X1  g676(.A(G8), .B1(new_n523), .B2(new_n527), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT122), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(KEYINPUT51), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1054), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1103), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1100), .A2(new_n1107), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1042), .A2(new_n1093), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n564), .A2(new_n1112), .A3(new_n573), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n564), .B2(new_n573), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT118), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n564), .A2(new_n1112), .A3(new_n573), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT56), .B(G2072), .Z(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1006), .A2(new_n990), .A3(new_n1010), .A4(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1051), .B2(G1956), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1063), .A2(G2067), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n851), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n610), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1130));
  AOI21_X1  g705(.A(G1956), .B1(new_n1130), .B2(new_n990), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n1009), .B(new_n978), .C1(new_n1015), .C2(new_n890), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1017), .A2(new_n1018), .B1(new_n1007), .B2(KEYINPUT45), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1121), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1131), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1125), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1139));
  INV_X1    g714(.A(G1956), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1007), .A2(KEYINPUT50), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n1142), .B2(new_n1047), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1143), .B2(new_n1123), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1138), .B1(new_n1136), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(new_n1123), .A3(new_n1139), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1125), .A2(KEYINPUT61), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT58), .B(G1341), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT120), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1063), .A2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT119), .B(G1996), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1006), .A2(new_n1010), .A3(new_n990), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT59), .B1(new_n1153), .B2(new_n541), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1155), .B(new_n623), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1145), .A2(new_n1147), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1128), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n610), .B1(new_n1128), .B2(new_n1159), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1126), .A2(new_n1127), .A3(KEYINPUT60), .A4(new_n920), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1160), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1137), .B1(new_n1158), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1111), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1110), .A2(KEYINPUT62), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1088), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1104), .A2(new_n1108), .A3(new_n1173), .A4(new_n1109), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1054), .B(G286), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1054), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1176), .B(KEYINPUT63), .C1(new_n1061), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1087), .A2(new_n1062), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT117), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI211_X1 g755(.A(new_n1054), .B(new_n1046), .C1(new_n1056), .C2(new_n1059), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1066), .A2(new_n1070), .A3(new_n1086), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT117), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1177), .A2(new_n1061), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1106), .A2(KEYINPUT63), .A3(new_n575), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1055), .A2(new_n1087), .A3(new_n1062), .A4(new_n1176), .ZN(new_n1188));
  XOR2_X1   g763(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1180), .A2(new_n1187), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1086), .A2(new_n1068), .A3(new_n931), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1079), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1181), .A2(new_n1087), .B1(new_n1193), .B2(new_n1067), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1175), .A2(new_n1191), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1005), .B1(new_n1169), .B2(new_n1195), .ZN(new_n1196));
  OR3_X1    g771(.A1(new_n991), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1197));
  OAI21_X1  g772(.A(KEYINPUT46), .B1(new_n991), .B2(G1996), .ZN(new_n1198));
  OR2_X1    g773(.A1(new_n994), .A2(new_n836), .ZN(new_n1199));
  AOI22_X1  g774(.A1(new_n1197), .A2(new_n1198), .B1(new_n998), .B2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n991), .A2(G1986), .A3(G290), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT48), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1202), .B1(new_n1003), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n997), .A2(new_n1001), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n803), .A2(G2067), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n991), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1196), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g785(.A1(new_n703), .A2(new_n705), .A3(G319), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n1212), .A2(KEYINPUT127), .ZN(new_n1213));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n1214));
  NAND4_X1  g788(.A1(new_n703), .A2(new_n705), .A3(new_n1214), .A4(G319), .ZN(new_n1215));
  NAND4_X1  g789(.A1(new_n1213), .A2(new_n676), .A3(new_n737), .A4(new_n1215), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1216), .B1(new_n911), .B2(new_n913), .ZN(new_n1217));
  AND3_X1   g791(.A1(new_n1217), .A2(new_n969), .A3(new_n972), .ZN(G308));
  NAND3_X1  g792(.A1(new_n1217), .A2(new_n969), .A3(new_n972), .ZN(G225));
endmodule


