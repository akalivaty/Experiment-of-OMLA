//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT77), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT76), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n207));
  OR2_X1    g006(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(G190gat), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(G169gat), .A3(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n210), .A2(new_n215), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n219), .A2(G169gat), .A3(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n218), .B2(new_n219), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n207), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT66), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n231), .B(new_n207), .C1(new_n223), .C2(new_n228), .ZN(new_n232));
  INV_X1    g031(.A(new_n223), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n224), .A2(new_n207), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n230), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT27), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n221), .B1(KEYINPUT67), .B2(KEYINPUT28), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT68), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT27), .B(G183gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(G190gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n243), .A2(KEYINPUT67), .A3(new_n248), .A4(KEYINPUT28), .ZN(new_n249));
  NOR2_X1   g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT26), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n251), .A2(new_n215), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n243), .A2(new_n248), .ZN(new_n254));
  NAND2_X1  g053(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT29), .B1(new_n236), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G226gat), .ZN(new_n259));
  INV_X1    g058(.A(G233gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n206), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G197gat), .B(G204gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(G211gat), .A2(G218gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT22), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(G211gat), .A2(G218gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n264), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT75), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(KEYINPUT75), .A3(new_n264), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n268), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n272), .A2(new_n267), .A3(KEYINPUT74), .A4(new_n273), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n236), .A2(new_n257), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n261), .ZN(new_n281));
  INV_X1    g080(.A(new_n261), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n229), .A2(KEYINPUT66), .B1(new_n233), .B2(new_n234), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n283), .A2(new_n232), .B1(new_n253), .B2(new_n256), .ZN(new_n284));
  OAI211_X1 g083(.A(KEYINPUT76), .B(new_n282), .C1(new_n284), .C2(KEYINPUT29), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n262), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n258), .A2(new_n261), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n284), .A2(new_n282), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n279), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n205), .B1(new_n290), .B2(KEYINPUT37), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT37), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n292), .B1(new_n286), .B2(new_n289), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT38), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G1gat), .B(G29gat), .Z(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G57gat), .B(G85gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  NAND2_X1  g098(.A1(G225gat), .A2(G233gat), .ZN(new_n300));
  AND2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G141gat), .B(G148gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(G155gat), .B2(G162gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G141gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G148gat), .ZN(new_n309));
  INV_X1    g108(.A(G148gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G141gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G155gat), .B(G162gat), .ZN(new_n313));
  INV_X1    g112(.A(G155gat), .ZN(new_n314));
  INV_X1    g113(.A(G162gat), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT2), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G134gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G127gat), .ZN(new_n322));
  INV_X1    g121(.A(G127gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G134gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G113gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G120gat), .ZN(new_n331));
  INV_X1    g130(.A(G120gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G113gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n333), .A3(new_n328), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n325), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT71), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT1), .B1(new_n325), .B2(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(G113gat), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n331), .ZN(new_n342));
  XNOR2_X1  g141(.A(G127gat), .B(G134gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT71), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n338), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n336), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n307), .A2(new_n317), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n320), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT71), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT71), .B1(new_n322), .B2(new_n324), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT1), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n332), .A2(G113gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n330), .A2(G120gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT69), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n326), .A3(new_n334), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n353), .A2(new_n342), .B1(new_n357), .B2(new_n325), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n350), .B1(new_n358), .B2(new_n318), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n318), .A2(new_n336), .A3(new_n345), .A4(new_n350), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n300), .B(new_n349), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  AND3_X1   g161(.A1(new_n338), .A2(new_n342), .A3(new_n344), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n331), .A2(new_n333), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT1), .B1(new_n364), .B2(KEYINPUT69), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n343), .B1(new_n365), .B2(new_n334), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n347), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n318), .A2(new_n336), .A3(new_n345), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(KEYINPUT78), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n300), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n346), .A2(new_n371), .A3(new_n347), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n362), .A2(new_n373), .A3(KEYINPUT5), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n368), .A2(KEYINPUT4), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n360), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT5), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n300), .A4(new_n349), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n299), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT6), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n362), .A2(new_n373), .A3(KEYINPUT5), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n299), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n380), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n205), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n286), .A2(new_n289), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n280), .A2(new_n261), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n262), .A2(new_n390), .A3(new_n285), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT82), .B1(new_n391), .B2(new_n279), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n287), .A2(new_n279), .A3(new_n288), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(KEYINPUT82), .A3(new_n279), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n292), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT38), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n397), .B(new_n205), .C1(new_n290), .C2(KEYINPUT37), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n294), .B(new_n389), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n387), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n286), .A2(new_n289), .A3(KEYINPUT30), .A4(new_n386), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n290), .A2(new_n205), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n401), .A2(new_n403), .A3(KEYINPUT81), .A4(new_n402), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n300), .B1(new_n376), .B2(new_n349), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n370), .B1(new_n369), .B2(new_n372), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT39), .ZN(new_n410));
  OR3_X1    g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n410), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n411), .A2(KEYINPUT40), .A3(new_n299), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n374), .A2(new_n378), .ZN(new_n414));
  INV_X1    g213(.A(new_n299), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT40), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(new_n299), .A3(new_n412), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n406), .A2(new_n407), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n318), .B2(new_n319), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n278), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G228gat), .A2(G233gat), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT29), .B1(new_n274), .B2(new_n267), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n268), .A2(new_n272), .A3(new_n273), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT3), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n424), .B(new_n425), .C1(new_n318), .C2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT29), .B1(new_n276), .B2(new_n277), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n347), .B1(new_n432), .B2(KEYINPUT3), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n429), .B(new_n431), .C1(new_n434), .C2(new_n425), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n425), .B1(new_n424), .B2(new_n433), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n428), .A2(new_n318), .ZN(new_n437));
  INV_X1    g236(.A(new_n425), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n437), .A2(new_n423), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n430), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G22gat), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n435), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n435), .B2(new_n440), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n399), .A2(new_n421), .A3(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G15gat), .B(G43gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n236), .A2(new_n257), .A3(new_n346), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n346), .B1(new_n236), .B2(new_n257), .ZN(new_n452));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n450), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n280), .A2(new_n358), .ZN(new_n458));
  INV_X1    g257(.A(new_n453), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n236), .A2(new_n257), .A3(new_n346), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT72), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT32), .B1(new_n449), .B2(new_n455), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n462), .B1(new_n461), .B2(new_n464), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n457), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n458), .A2(new_n460), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(new_n453), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n468), .B(new_n453), .C1(new_n451), .C2(new_n452), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n470), .A2(new_n472), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT72), .B1(new_n454), .B2(new_n463), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n478), .B2(new_n457), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT73), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481));
  INV_X1    g280(.A(new_n456), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n449), .B1(new_n461), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n476), .B2(new_n477), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT73), .B1(new_n484), .B2(new_n475), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n445), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT80), .B1(new_n384), .B2(new_n379), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n378), .A2(new_n299), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT6), .B1(new_n490), .B2(new_n374), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n416), .A3(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n489), .A2(new_n493), .A3(new_n380), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n488), .B1(new_n494), .B2(new_n404), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n467), .A2(new_n473), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n475), .A3(new_n457), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n481), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n487), .A2(new_n495), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n446), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(new_n497), .A3(new_n445), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT83), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n494), .A2(new_n404), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n496), .A2(new_n445), .A3(new_n497), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(new_n496), .B2(new_n497), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n445), .A2(new_n385), .A3(new_n510), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n509), .A2(new_n511), .A3(new_n485), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n406), .A2(new_n407), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n507), .A2(KEYINPUT35), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n501), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G15gat), .B(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT16), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(G1gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G1gat), .B2(new_n516), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(G8gat), .Z(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR3_X1   g320(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT87), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n523), .B(KEYINPUT87), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT88), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n527), .A2(new_n529), .B1(G29gat), .B2(G36gat), .ZN(new_n530));
  INV_X1    g329(.A(G43gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(G50gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G50gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(G43gat), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n522), .A2(KEYINPUT90), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n522), .A2(KEYINPUT90), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n525), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT89), .B(G50gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(G43gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n533), .B1(new_n542), .B2(new_n532), .ZN(new_n543));
  NAND2_X1  g342(.A1(G29gat), .A2(G36gat), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n540), .A2(new_n543), .A3(new_n536), .A4(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT17), .B1(new_n537), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n548), .B(new_n545), .C1(new_n530), .C2(new_n536), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n521), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n537), .A2(new_n546), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(new_n520), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n551), .A2(KEYINPUT18), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n552), .B(new_n520), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n555), .B(KEYINPUT13), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n555), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n550), .A2(new_n553), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n556), .B(new_n559), .C1(new_n561), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n556), .A2(KEYINPUT92), .A3(new_n559), .ZN(new_n565));
  XNOR2_X1  g364(.A(G169gat), .B(G197gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT85), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G113gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT86), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n568), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT12), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n564), .A2(new_n565), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n561), .A2(new_n563), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n561), .A2(KEYINPUT18), .B1(new_n557), .B2(new_n558), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n576), .B(new_n577), .C1(KEYINPUT92), .C2(new_n573), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n515), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT93), .ZN(new_n583));
  NAND2_X1  g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n583), .A2(KEYINPUT9), .ZN(new_n587));
  OAI221_X1 g386(.A(new_n585), .B1(new_n583), .B2(new_n584), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT94), .B(G57gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(G64gat), .ZN(new_n590));
  INV_X1    g389(.A(G64gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(G57gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n584), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT95), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT95), .B1(new_n593), .B2(new_n595), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n588), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(KEYINPUT21), .ZN(new_n602));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  AOI21_X1  g403(.A(new_n521), .B1(new_n601), .B2(KEYINPUT21), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT97), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT96), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G183gat), .B(G211gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n606), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n552), .ZN(new_n618));
  NAND2_X1  g417(.A1(G85gat), .A2(G92gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT7), .ZN(new_n620));
  NAND2_X1  g419(.A1(G99gat), .A2(G106gat), .ZN(new_n621));
  INV_X1    g420(.A(G85gat), .ZN(new_n622));
  INV_X1    g421(.A(G92gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(KEYINPUT8), .A2(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G99gat), .B(G106gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n618), .A2(new_n627), .B1(KEYINPUT41), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n547), .A2(new_n549), .ZN(new_n630));
  INV_X1    g429(.A(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n617), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G134gat), .B(G162gat), .Z(new_n635));
  NOR2_X1   g434(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(KEYINPUT98), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n629), .A2(new_n632), .A3(new_n617), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n634), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n637), .B(KEYINPUT98), .Z(new_n641));
  INV_X1    g440(.A(new_n639), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n641), .B1(new_n642), .B2(new_n633), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n600), .A2(new_n631), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n627), .B(new_n588), .C1(new_n598), .C2(new_n599), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n627), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n650), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n647), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n662), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n654), .A2(new_n656), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n663), .A2(KEYINPUT101), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT101), .B1(new_n663), .B2(new_n665), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n615), .A2(new_n645), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n581), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n494), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT102), .B(G1gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1324gat));
  NOR2_X1   g475(.A1(new_n672), .A2(new_n513), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(KEYINPUT42), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(KEYINPUT104), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n678), .B(KEYINPUT103), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n677), .B1(KEYINPUT42), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n683), .B2(G8gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n679), .A2(KEYINPUT104), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n680), .A2(new_n684), .A3(new_n685), .ZN(G1325gat));
  NAND2_X1  g485(.A1(new_n496), .A2(new_n497), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n485), .B1(new_n687), .B2(KEYINPUT73), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n498), .B1(new_n688), .B2(new_n481), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n672), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n688), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(G15gat), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n690), .B1(new_n672), .B2(new_n692), .ZN(G1326gat));
  NOR2_X1   g492(.A1(new_n672), .A2(new_n445), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT43), .B(G22gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  NOR3_X1   g495(.A1(new_n670), .A2(new_n614), .A3(new_n644), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT105), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n581), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n699), .A2(G29gat), .A3(new_n673), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT45), .Z(new_n701));
  NAND2_X1  g500(.A1(new_n495), .A2(KEYINPUT107), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n703), .B(new_n488), .C1(new_n494), .C2(new_n404), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n399), .A2(new_n421), .A3(new_n445), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n705), .A2(new_n706), .A3(new_n689), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n645), .B1(new_n707), .B2(new_n514), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n644), .A2(new_n709), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n501), .B2(new_n514), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n669), .B(KEYINPUT106), .Z(new_n713));
  NOR3_X1   g512(.A1(new_n713), .A2(new_n580), .A3(new_n614), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n673), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n716), .ZN(G1328gat));
  NOR3_X1   g516(.A1(new_n699), .A2(G36gat), .A3(new_n513), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT46), .ZN(new_n719));
  OAI21_X1  g518(.A(G36gat), .B1(new_n715), .B2(new_n513), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1329gat));
  OAI21_X1  g520(.A(new_n531), .B1(new_n699), .B2(new_n691), .ZN(new_n722));
  INV_X1    g521(.A(new_n689), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G43gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n715), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g525(.A(new_n541), .B1(new_n699), .B2(new_n445), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n445), .A2(new_n541), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n715), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n615), .A2(new_n645), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n713), .A2(new_n580), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n507), .A2(KEYINPUT35), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n512), .A2(new_n513), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n705), .A2(new_n706), .A3(new_n689), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n494), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(new_n589), .Z(G1332gat));
  INV_X1    g538(.A(new_n513), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n741), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT108), .ZN(G1333gat));
  NAND2_X1  g545(.A1(new_n737), .A2(new_n723), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n691), .A2(G71gat), .ZN(new_n748));
  AOI22_X1  g547(.A1(new_n747), .A2(G71gat), .B1(new_n737), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n737), .A2(new_n488), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  OR3_X1    g553(.A1(new_n614), .A2(KEYINPUT110), .A3(new_n579), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT110), .B1(new_n614), .B2(new_n579), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n644), .B1(new_n736), .B2(new_n735), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI211_X1 g559(.A(KEYINPUT112), .B(new_n644), .C1(new_n736), .C2(new_n735), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n754), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n708), .A2(KEYINPUT112), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n758), .A2(new_n759), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n763), .A2(KEYINPUT51), .A3(new_n757), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n766), .A2(new_n622), .A3(new_n494), .A4(new_n670), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n669), .B1(new_n755), .B2(new_n756), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n710), .A2(new_n768), .A3(new_n712), .A4(new_n769), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n712), .B(new_n769), .C1(new_n758), .C2(KEYINPUT44), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT111), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n494), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n767), .B1(new_n774), .B2(new_n622), .ZN(G1336gat));
  INV_X1    g574(.A(new_n713), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n513), .A2(G92gat), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n776), .B(new_n778), .C1(new_n762), .C2(new_n765), .ZN(new_n779));
  INV_X1    g578(.A(new_n771), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n623), .B1(new_n780), .B2(new_n740), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n779), .A2(KEYINPUT52), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n770), .A2(new_n772), .A3(new_n740), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n783), .A2(new_n784), .A3(G92gat), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n783), .B2(G92gat), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n785), .A2(new_n786), .A3(new_n779), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(G1337gat));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n723), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G99gat), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n691), .A2(G99gat), .A3(new_n669), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n766), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1338gat));
  AOI21_X1  g593(.A(new_n776), .B1(new_n762), .B2(new_n765), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n445), .A2(G106gat), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n488), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT53), .B1(new_n798), .B2(G106gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n773), .A2(new_n488), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n801), .A2(G106gat), .B1(new_n795), .B2(new_n796), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(G1339gat));
  NOR2_X1   g603(.A1(new_n740), .A2(new_n673), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n555), .B1(new_n551), .B2(new_n554), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n557), .A2(new_n558), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n572), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI221_X1 g608(.A(new_n809), .B1(new_n574), .B2(new_n564), .C1(new_n667), .C2(new_n668), .ZN(new_n810));
  INV_X1    g609(.A(new_n665), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n651), .A2(new_n652), .A3(new_n647), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n664), .B1(new_n653), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n654), .A2(KEYINPUT114), .A3(KEYINPUT54), .A4(new_n812), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n811), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n818), .A4(new_n817), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n579), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n645), .B1(new_n810), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n809), .B1(new_n564), .B2(new_n574), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n644), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n822), .A3(new_n821), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n615), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n671), .A2(new_n580), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n806), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n503), .A2(new_n506), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n330), .B1(new_n833), .B2(new_n580), .ZN(new_n834));
  AOI211_X1 g633(.A(new_n488), .B(new_n691), .C1(new_n829), .C2(new_n830), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n805), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n579), .A2(G113gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT116), .ZN(G1340gat));
  OAI21_X1  g639(.A(G120gat), .B1(new_n837), .B2(new_n776), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n670), .A2(new_n339), .A3(new_n340), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n833), .B2(new_n842), .ZN(G1341gat));
  OAI21_X1  g642(.A(G127gat), .B1(new_n837), .B2(new_n615), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n614), .A2(new_n323), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n833), .B2(new_n845), .ZN(G1342gat));
  OAI21_X1  g645(.A(G134gat), .B1(new_n837), .B2(new_n644), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n833), .A2(G134gat), .A3(new_n644), .ZN(new_n848));
  XOR2_X1   g647(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n849));
  OR2_X1    g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(G1343gat));
  AND3_X1   g651(.A1(new_n831), .A2(new_n488), .A3(new_n689), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n580), .A2(G141gat), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(KEYINPUT118), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n806), .A2(new_n723), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n445), .B1(new_n829), .B2(new_n830), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT57), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(KEYINPUT57), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n579), .B(new_n858), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n857), .B1(G141gat), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n856), .A2(KEYINPUT118), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(G1344gat));
  NAND3_X1  g665(.A1(new_n853), .A2(new_n310), .A3(new_n670), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n861), .A2(new_n862), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n670), .A3(new_n858), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n869), .A2(new_n870), .A3(G148gat), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n810), .A2(new_n823), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n872), .B(new_n827), .C1(new_n873), .C2(new_n645), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT119), .B1(new_n824), .B2(new_n828), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n615), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n445), .B1(new_n876), .B2(new_n830), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n860), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n670), .A3(new_n858), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n870), .B1(new_n879), .B2(G148gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n867), .B1(new_n871), .B2(new_n880), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n853), .A2(new_n314), .A3(new_n614), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n868), .A2(new_n614), .A3(new_n858), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(new_n314), .ZN(G1346gat));
  NAND3_X1  g684(.A1(new_n853), .A2(new_n315), .A3(new_n645), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n645), .A3(new_n858), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G162gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n513), .A2(new_n494), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n832), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n829), .B2(new_n830), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n216), .A3(new_n579), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT121), .Z(new_n896));
  NAND2_X1  g695(.A1(new_n835), .A2(new_n892), .ZN(new_n897));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897), .B2(new_n580), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1348gat));
  OAI21_X1  g698(.A(G176gat), .B1(new_n897), .B2(new_n776), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n894), .A2(new_n217), .A3(new_n670), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1349gat));
  OAI21_X1  g701(.A(G183gat), .B1(new_n897), .B2(new_n615), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n894), .A2(new_n244), .A3(new_n614), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g705(.A1(new_n835), .A2(new_n645), .A3(new_n892), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G190gat), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n908), .A2(KEYINPUT123), .A3(KEYINPUT61), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(KEYINPUT61), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT123), .B1(new_n908), .B2(KEYINPUT61), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n909), .A2(new_n912), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n894), .A2(new_n221), .A3(new_n645), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1351gat));
  AND2_X1   g716(.A1(new_n689), .A2(new_n892), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n859), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(G197gat), .B1(new_n919), .B2(new_n579), .ZN(new_n920));
  INV_X1    g719(.A(new_n878), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n918), .B(KEYINPUT124), .Z(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n579), .A2(G197gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(G1352gat));
  INV_X1    g724(.A(G204gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n926), .A3(new_n670), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n927), .B(KEYINPUT62), .Z(new_n928));
  NOR3_X1   g727(.A1(new_n921), .A2(new_n776), .A3(new_n922), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n926), .B2(new_n929), .ZN(G1353gat));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n918), .A2(new_n614), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n878), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n878), .A2(new_n931), .A3(new_n933), .ZN(new_n936));
  NOR2_X1   g735(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n935), .A2(G211gat), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G211gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n859), .A2(new_n939), .A3(new_n933), .ZN(new_n940));
  INV_X1    g739(.A(new_n936), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n941), .A2(new_n934), .A3(new_n939), .ZN(new_n942));
  XNOR2_X1  g741(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n938), .B(new_n940), .C1(new_n942), .C2(new_n943), .ZN(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n919), .B2(new_n645), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n645), .A2(G218gat), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT127), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n945), .B1(new_n923), .B2(new_n947), .ZN(G1355gat));
endmodule


