

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  XNOR2_X1 U324 ( .A(n335), .B(n334), .ZN(n370) );
  XNOR2_X1 U325 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n331) );
  NOR2_X1 U326 ( .A1(n586), .A2(n414), .ZN(n416) );
  XNOR2_X1 U327 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U328 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U329 ( .A(n450), .B(KEYINPUT101), .ZN(n451) );
  INV_X1 U330 ( .A(KEYINPUT38), .ZN(n450) );
  XOR2_X1 U331 ( .A(G64GAT), .B(G204GAT), .Z(n292) );
  AND2_X1 U332 ( .A1(n563), .A2(n554), .ZN(n464) );
  INV_X1 U333 ( .A(KEYINPUT88), .ZN(n332) );
  XNOR2_X1 U334 ( .A(n436), .B(n435), .ZN(n438) );
  INV_X1 U335 ( .A(KEYINPUT77), .ZN(n340) );
  XNOR2_X1 U336 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U337 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U338 ( .A(KEYINPUT26), .B(n385), .ZN(n573) );
  XNOR2_X1 U339 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U340 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U341 ( .A(n579), .B(KEYINPUT41), .Z(n554) );
  XOR2_X1 U342 ( .A(n380), .B(n379), .Z(n477) );
  INV_X1 U343 ( .A(G190GAT), .ZN(n480) );
  XNOR2_X1 U344 ( .A(n452), .B(n451), .ZN(n500) );
  XNOR2_X1 U345 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U346 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U347 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n294) );
  XNOR2_X1 U350 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n308) );
  XNOR2_X1 U352 ( .A(G50GAT), .B(G162GAT), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n295), .B(KEYINPUT76), .ZN(n366) );
  XOR2_X1 U354 ( .A(G36GAT), .B(G190GAT), .Z(n337) );
  XOR2_X1 U355 ( .A(n366), .B(n337), .Z(n297) );
  NAND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U357 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U358 ( .A(G106GAT), .B(KEYINPUT65), .Z(n299) );
  XNOR2_X1 U359 ( .A(G134GAT), .B(G92GAT), .ZN(n298) );
  XNOR2_X1 U360 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U361 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U362 ( .A(G29GAT), .B(G43GAT), .Z(n303) );
  XNOR2_X1 U363 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n302) );
  XNOR2_X1 U364 ( .A(n303), .B(n302), .ZN(n422) );
  XNOR2_X1 U365 ( .A(G99GAT), .B(G85GAT), .ZN(n304) );
  XNOR2_X1 U366 ( .A(n304), .B(KEYINPUT73), .ZN(n439) );
  XNOR2_X1 U367 ( .A(n422), .B(n439), .ZN(n305) );
  XNOR2_X1 U368 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n561) );
  INV_X1 U370 ( .A(n561), .ZN(n485) );
  XNOR2_X1 U371 ( .A(KEYINPUT36), .B(n485), .ZN(n586) );
  XOR2_X1 U372 ( .A(G211GAT), .B(G155GAT), .Z(n310) );
  XNOR2_X1 U373 ( .A(G127GAT), .B(G183GAT), .ZN(n309) );
  XNOR2_X1 U374 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G64GAT), .Z(n312) );
  XNOR2_X1 U376 ( .A(G8GAT), .B(KEYINPUT77), .ZN(n311) );
  XNOR2_X1 U377 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U378 ( .A(n314), .B(n313), .Z(n319) );
  XOR2_X1 U379 ( .A(KEYINPUT78), .B(KEYINPUT80), .Z(n316) );
  NAND2_X1 U380 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U381 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U382 ( .A(KEYINPUT79), .B(n317), .ZN(n318) );
  XNOR2_X1 U383 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U384 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n321) );
  XNOR2_X1 U385 ( .A(G71GAT), .B(KEYINPUT14), .ZN(n320) );
  XNOR2_X1 U386 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U387 ( .A(n323), .B(n322), .Z(n327) );
  XNOR2_X1 U388 ( .A(G1GAT), .B(G22GAT), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n324), .B(G15GAT), .ZN(n417) );
  XNOR2_X1 U390 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n325) );
  XNOR2_X1 U391 ( .A(n325), .B(KEYINPUT13), .ZN(n446) );
  XNOR2_X1 U392 ( .A(n417), .B(n446), .ZN(n326) );
  XNOR2_X1 U393 ( .A(n327), .B(n326), .ZN(n484) );
  XOR2_X1 U394 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n329) );
  XNOR2_X1 U395 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n328) );
  XNOR2_X1 U396 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U397 ( .A(KEYINPUT18), .B(n330), .Z(n362) );
  XNOR2_X1 U398 ( .A(n331), .B(KEYINPUT89), .ZN(n335) );
  XNOR2_X1 U399 ( .A(G197GAT), .B(G218GAT), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n362), .B(n370), .ZN(n345) );
  XNOR2_X1 U401 ( .A(G176GAT), .B(G92GAT), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n292), .B(n336), .ZN(n447) );
  XOR2_X1 U403 ( .A(n337), .B(n447), .Z(n339) );
  NAND2_X1 U404 ( .A1(G226GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U406 ( .A(G169GAT), .B(G8GAT), .Z(n418) );
  XNOR2_X1 U407 ( .A(n418), .B(KEYINPUT92), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n507) );
  XNOR2_X1 U409 ( .A(G127GAT), .B(KEYINPUT81), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n346), .B(KEYINPUT0), .ZN(n347) );
  XOR2_X1 U411 ( .A(n347), .B(KEYINPUT82), .Z(n349) );
  XNOR2_X1 U412 ( .A(G113GAT), .B(G134GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n403) );
  XOR2_X1 U414 ( .A(G99GAT), .B(G190GAT), .Z(n351) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(G43GAT), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U417 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n353) );
  XNOR2_X1 U418 ( .A(G15GAT), .B(G176GAT), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U420 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U421 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XOR2_X1 U422 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n357) );
  NAND2_X1 U423 ( .A1(G227GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n434), .B(n358), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n403), .B(n361), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n534) );
  INV_X1 U429 ( .A(n534), .ZN(n509) );
  NOR2_X1 U430 ( .A1(n507), .A2(n509), .ZN(n381) );
  XOR2_X1 U431 ( .A(KEYINPUT72), .B(G78GAT), .Z(n365) );
  XNOR2_X1 U432 ( .A(G148GAT), .B(G106GAT), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n436) );
  XOR2_X1 U434 ( .A(n436), .B(n366), .Z(n372) );
  XOR2_X1 U435 ( .A(KEYINPUT90), .B(KEYINPUT3), .Z(n368) );
  XNOR2_X1 U436 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n367) );
  XNOR2_X1 U437 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U438 ( .A(G141GAT), .B(n369), .Z(n397) );
  XNOR2_X1 U439 ( .A(n397), .B(n370), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n372), .B(n371), .ZN(n380) );
  NAND2_X1 U441 ( .A1(G228GAT), .A2(G233GAT), .ZN(n378) );
  XOR2_X1 U442 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n374) );
  XNOR2_X1 U443 ( .A(KEYINPUT87), .B(KEYINPUT24), .ZN(n373) );
  XNOR2_X1 U444 ( .A(n374), .B(n373), .ZN(n376) );
  XOR2_X1 U445 ( .A(G22GAT), .B(G204GAT), .Z(n375) );
  XNOR2_X1 U446 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n378), .B(n377), .ZN(n379) );
  NOR2_X1 U448 ( .A1(n381), .A2(n477), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n382), .B(KEYINPUT25), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n383), .B(KEYINPUT95), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n507), .B(KEYINPUT27), .ZN(n407) );
  NAND2_X1 U452 ( .A1(n477), .A2(n509), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n384), .B(KEYINPUT94), .ZN(n385) );
  NOR2_X1 U454 ( .A1(n407), .A2(n573), .ZN(n386) );
  NOR2_X1 U455 ( .A1(n387), .A2(n386), .ZN(n404) );
  XOR2_X1 U456 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n389) );
  XNOR2_X1 U457 ( .A(G120GAT), .B(G148GAT), .ZN(n388) );
  XNOR2_X1 U458 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U459 ( .A(KEYINPUT91), .B(KEYINPUT4), .Z(n391) );
  XNOR2_X1 U460 ( .A(G1GAT), .B(G162GAT), .ZN(n390) );
  XNOR2_X1 U461 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U462 ( .A(n393), .B(n392), .ZN(n401) );
  XOR2_X1 U463 ( .A(G57GAT), .B(KEYINPUT5), .Z(n395) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U465 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U466 ( .A(n396), .B(G85GAT), .Z(n399) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(n397), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n503) );
  INV_X1 U471 ( .A(n503), .ZN(n517) );
  NOR2_X1 U472 ( .A1(n404), .A2(n517), .ZN(n406) );
  INV_X1 U473 ( .A(KEYINPUT96), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n406), .B(n405), .ZN(n412) );
  NOR2_X1 U475 ( .A1(n503), .A2(n407), .ZN(n529) );
  XOR2_X1 U476 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n408) );
  XNOR2_X1 U477 ( .A(n477), .B(n408), .ZN(n533) );
  NAND2_X1 U478 ( .A1(n529), .A2(n533), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n409), .B(KEYINPUT93), .ZN(n410) );
  NAND2_X1 U480 ( .A1(n410), .A2(n509), .ZN(n411) );
  NAND2_X1 U481 ( .A1(n412), .A2(n411), .ZN(n488) );
  NAND2_X1 U482 ( .A1(n484), .A2(n488), .ZN(n413) );
  XOR2_X1 U483 ( .A(KEYINPUT99), .B(n413), .Z(n414) );
  XOR2_X1 U484 ( .A(KEYINPUT37), .B(KEYINPUT100), .Z(n415) );
  XNOR2_X1 U485 ( .A(n416), .B(n415), .ZN(n515) );
  XOR2_X1 U486 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U487 ( .A1(G229GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U489 ( .A(n421), .B(KEYINPUT30), .Z(n424) );
  XNOR2_X1 U490 ( .A(n422), .B(KEYINPUT67), .ZN(n423) );
  XNOR2_X1 U491 ( .A(n424), .B(n423), .ZN(n432) );
  XOR2_X1 U492 ( .A(G113GAT), .B(G141GAT), .Z(n426) );
  XNOR2_X1 U493 ( .A(G36GAT), .B(G50GAT), .ZN(n425) );
  XNOR2_X1 U494 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U495 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n428) );
  XNOR2_X1 U496 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n427) );
  XNOR2_X1 U497 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U498 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U499 ( .A(n432), .B(n431), .ZN(n563) );
  INV_X1 U500 ( .A(n563), .ZN(n575) );
  AND2_X1 U501 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  INV_X1 U502 ( .A(KEYINPUT32), .ZN(n437) );
  XNOR2_X1 U503 ( .A(n438), .B(n437), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n439), .B(KEYINPUT75), .ZN(n443) );
  XOR2_X1 U505 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n441) );
  XNOR2_X1 U506 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n440) );
  XOR2_X1 U507 ( .A(n441), .B(n440), .Z(n442) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n579) );
  NOR2_X1 U510 ( .A1(n575), .A2(n579), .ZN(n489) );
  NAND2_X1 U511 ( .A1(n515), .A2(n489), .ZN(n452) );
  NOR2_X1 U512 ( .A1(n500), .A2(n509), .ZN(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n454) );
  INV_X1 U514 ( .A(G43GAT), .ZN(n453) );
  NOR2_X1 U515 ( .A1(n500), .A2(n503), .ZN(n458) );
  XNOR2_X1 U516 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n458), .B(n457), .ZN(G1328GAT) );
  INV_X1 U518 ( .A(KEYINPUT48), .ZN(n473) );
  NOR2_X1 U519 ( .A1(n484), .A2(n586), .ZN(n460) );
  XNOR2_X1 U520 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n459) );
  XNOR2_X1 U521 ( .A(n460), .B(n459), .ZN(n461) );
  NOR2_X1 U522 ( .A1(n461), .A2(n579), .ZN(n462) );
  XNOR2_X1 U523 ( .A(KEYINPUT112), .B(n462), .ZN(n463) );
  NAND2_X1 U524 ( .A1(n463), .A2(n575), .ZN(n471) );
  XOR2_X1 U525 ( .A(KEYINPUT47), .B(KEYINPUT110), .Z(n469) );
  XOR2_X1 U526 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(n464), .ZN(n466) );
  NOR2_X1 U528 ( .A1(n561), .A2(n466), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n467), .A2(n484), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n531) );
  NOR2_X1 U533 ( .A1(n531), .A2(n507), .ZN(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT54), .B(n474), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n475), .A2(n503), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(KEYINPUT64), .ZN(n572) );
  NOR2_X1 U537 ( .A1(n572), .A2(n477), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(KEYINPUT55), .ZN(n479) );
  NOR2_X2 U539 ( .A1(n509), .A2(n479), .ZN(n570) );
  NAND2_X1 U540 ( .A1(n570), .A2(n561), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n481) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n492) );
  INV_X1 U543 ( .A(n484), .ZN(n583) );
  NAND2_X1 U544 ( .A1(n485), .A2(n583), .ZN(n486) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(n486), .Z(n487) );
  AND2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n502) );
  NAND2_X1 U547 ( .A1(n489), .A2(n502), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT97), .B(n490), .ZN(n497) );
  NAND2_X1 U549 ( .A1(n517), .A2(n497), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(G1324GAT) );
  INV_X1 U551 ( .A(n507), .ZN(n520) );
  NAND2_X1 U552 ( .A1(n520), .A2(n497), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT98), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n494), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U556 ( .A1(n497), .A2(n534), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  INV_X1 U558 ( .A(n533), .ZN(n524) );
  NAND2_X1 U559 ( .A1(n524), .A2(n497), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U561 ( .A1(n507), .A2(n500), .ZN(n499) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  NOR2_X1 U563 ( .A1(n533), .A2(n500), .ZN(n501) );
  XOR2_X1 U564 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  XOR2_X1 U565 ( .A(n554), .B(KEYINPUT103), .Z(n566) );
  AND2_X1 U566 ( .A1(n575), .A2(n566), .ZN(n514) );
  NAND2_X1 U567 ( .A1(n514), .A2(n502), .ZN(n511) );
  NOR2_X1 U568 ( .A1(n503), .A2(n511), .ZN(n505) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n506), .Z(G1332GAT) );
  NOR2_X1 U572 ( .A1(n507), .A2(n511), .ZN(n508) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n508), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n509), .A2(n511), .ZN(n510) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n510), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n533), .A2(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(KEYINPUT105), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n525), .A2(n517), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT106), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n525), .A2(n520), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  XOR2_X1 U586 ( .A(G99GAT), .B(KEYINPUT107), .Z(n523) );
  NAND2_X1 U587 ( .A1(n525), .A2(n534), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n527) );
  NAND2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n528), .Z(G1339GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n537) );
  INV_X1 U594 ( .A(n529), .ZN(n530) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U596 ( .A(KEYINPUT113), .B(n532), .ZN(n549) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n549), .A2(n535), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n545), .A2(n563), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n540) );
  NAND2_X1 U603 ( .A1(n545), .A2(n566), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n543) );
  NAND2_X1 U607 ( .A1(n545), .A2(n583), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n547) );
  NAND2_X1 U611 ( .A1(n545), .A2(n561), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n548), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n573), .A2(n549), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT119), .B(n550), .Z(n560) );
  AND2_X1 U616 ( .A1(n563), .A2(n560), .ZN(n552) );
  XNOR2_X1 U617 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U621 ( .A1(n560), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n583), .A2(n560), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT122), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT123), .Z(n565) );
  NAND2_X1 U630 ( .A1(n570), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n570), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n583), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(KEYINPUT125), .ZN(n585) );
  NOR2_X1 U640 ( .A1(n575), .A2(n585), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  INV_X1 U645 ( .A(n585), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n582), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(G218GAT), .B(n589), .Z(G1355GAT) );
endmodule

