

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751;

  AND2_X1 U374 ( .A1(n621), .A2(n620), .ZN(n699) );
  AND2_X1 U375 ( .A1(n551), .A2(n662), .ZN(n355) );
  BUF_X1 U376 ( .A(G953), .Z(n351) );
  XNOR2_X1 U377 ( .A(n721), .B(n513), .ZN(n506) );
  XNOR2_X1 U378 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X2 U379 ( .A(KEYINPUT4), .B(KEYINPUT76), .ZN(n433) );
  XNOR2_X2 U380 ( .A(n590), .B(n400), .ZN(n582) );
  XOR2_X2 U381 ( .A(G110), .B(G104), .Z(n437) );
  XNOR2_X2 U382 ( .A(n382), .B(n459), .ZN(n531) );
  XNOR2_X2 U383 ( .A(G143), .B(G128), .ZN(n427) );
  XNOR2_X1 U384 ( .A(n418), .B(n499), .ZN(n736) );
  XNOR2_X1 U385 ( .A(n394), .B(G125), .ZN(n464) );
  BUF_X1 U386 ( .A(n696), .Z(n352) );
  BUF_X1 U387 ( .A(n590), .Z(n353) );
  INV_X1 U388 ( .A(n429), .ZN(n354) );
  XNOR2_X1 U389 ( .A(n427), .B(n426), .ZN(n467) );
  XNOR2_X2 U390 ( .A(n483), .B(n482), .ZN(n551) );
  NAND2_X1 U391 ( .A1(n565), .A2(n677), .ZN(n454) );
  XNOR2_X1 U392 ( .A(n450), .B(n449), .ZN(n565) );
  BUF_X1 U393 ( .A(n582), .Z(n356) );
  XNOR2_X2 U394 ( .A(n454), .B(KEYINPUT89), .ZN(n590) );
  INV_X1 U395 ( .A(G902), .ZN(n519) );
  NAND2_X1 U396 ( .A1(n533), .A2(n537), .ZN(n680) );
  INV_X1 U397 ( .A(KEYINPUT19), .ZN(n400) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n510) );
  XOR2_X1 U399 ( .A(KEYINPUT66), .B(G131), .Z(n500) );
  NOR2_X1 U400 ( .A1(n645), .A2(n649), .ZN(n682) );
  INV_X1 U401 ( .A(KEYINPUT88), .ZN(n407) );
  INV_X1 U402 ( .A(G237), .ZN(n446) );
  INV_X1 U403 ( .A(KEYINPUT79), .ZN(n426) );
  XNOR2_X1 U404 ( .A(n521), .B(n520), .ZN(n524) );
  XNOR2_X1 U405 ( .A(G113), .B(KEYINPUT68), .ZN(n440) );
  INV_X1 U406 ( .A(KEYINPUT7), .ZN(n469) );
  XOR2_X1 U407 ( .A(G122), .B(KEYINPUT9), .Z(n470) );
  NAND2_X1 U408 ( .A1(n540), .A2(n417), .ZN(n401) );
  NAND2_X1 U409 ( .A1(n532), .A2(KEYINPUT34), .ZN(n416) );
  XNOR2_X1 U410 ( .A(n466), .B(n395), .ZN(n537) );
  XNOR2_X1 U411 ( .A(n465), .B(n396), .ZN(n395) );
  INV_X1 U412 ( .A(G475), .ZN(n396) );
  INV_X1 U413 ( .A(KEYINPUT1), .ZN(n412) );
  BUF_X1 U414 ( .A(n524), .Z(n669) );
  NOR2_X1 U415 ( .A1(n751), .A2(n750), .ZN(n610) );
  XNOR2_X1 U416 ( .A(KEYINPUT65), .B(G101), .ZN(n513) );
  XOR2_X1 U417 ( .A(G146), .B(KEYINPUT5), .Z(n512) );
  INV_X1 U418 ( .A(G146), .ZN(n394) );
  XNOR2_X1 U419 ( .A(G143), .B(G113), .ZN(n389) );
  XNOR2_X1 U420 ( .A(G104), .B(G122), .ZN(n462) );
  XNOR2_X1 U421 ( .A(n463), .B(n500), .ZN(n392) );
  XNOR2_X1 U422 ( .A(n460), .B(n461), .ZN(n390) );
  XOR2_X1 U423 ( .A(KEYINPUT103), .B(KEYINPUT12), .Z(n461) );
  XNOR2_X1 U424 ( .A(KEYINPUT15), .B(G902), .ZN(n623) );
  XOR2_X1 U425 ( .A(G146), .B(G140), .Z(n504) );
  XNOR2_X1 U426 ( .A(n501), .B(G137), .ZN(n418) );
  XOR2_X1 U427 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n434) );
  NAND2_X1 U428 ( .A1(G234), .A2(G237), .ZN(n456) );
  XNOR2_X1 U429 ( .A(n385), .B(n384), .ZN(n621) );
  INV_X1 U430 ( .A(KEYINPUT48), .ZN(n384) );
  XNOR2_X1 U431 ( .A(n453), .B(n452), .ZN(n677) );
  XNOR2_X1 U432 ( .A(KEYINPUT64), .B(KEYINPUT0), .ZN(n459) );
  NOR2_X1 U433 ( .A1(n680), .A2(n479), .ZN(n480) );
  BUF_X1 U434 ( .A(n699), .Z(n739) );
  INV_X1 U435 ( .A(G107), .ZN(n436) );
  XNOR2_X1 U436 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n486) );
  XNOR2_X1 U437 ( .A(G137), .B(G128), .ZN(n484) );
  XNOR2_X1 U438 ( .A(n464), .B(n393), .ZN(n737) );
  XNOR2_X1 U439 ( .A(G140), .B(KEYINPUT10), .ZN(n393) );
  XNOR2_X1 U440 ( .A(n391), .B(n387), .ZN(n629) );
  XNOR2_X1 U441 ( .A(n390), .B(n388), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n737), .B(n392), .ZN(n391) );
  XNOR2_X1 U443 ( .A(n462), .B(n389), .ZN(n388) );
  INV_X1 U444 ( .A(n623), .ZN(n409) );
  XNOR2_X1 U445 ( .A(n419), .B(n736), .ZN(n712) );
  XNOR2_X1 U446 ( .A(n508), .B(n502), .ZN(n419) );
  XNOR2_X1 U447 ( .A(n735), .B(KEYINPUT74), .ZN(n502) );
  XNOR2_X1 U448 ( .A(n507), .B(n506), .ZN(n508) );
  NAND2_X1 U449 ( .A1(n614), .A2(n411), .ZN(n615) );
  XNOR2_X1 U450 ( .A(KEYINPUT16), .B(G122), .ZN(n442) );
  XNOR2_X1 U451 ( .A(G116), .B(G107), .ZN(n473) );
  NOR2_X1 U452 ( .A1(n592), .A2(n411), .ZN(n658) );
  XNOR2_X1 U453 ( .A(n535), .B(KEYINPUT35), .ZN(n749) );
  XNOR2_X1 U454 ( .A(n397), .B(n362), .ZN(n632) );
  NOR2_X2 U455 ( .A1(n604), .A2(n568), .ZN(n648) );
  XNOR2_X1 U456 ( .A(n536), .B(KEYINPUT105), .ZN(n645) );
  INV_X1 U457 ( .A(KEYINPUT109), .ZN(n422) );
  AND2_X1 U458 ( .A1(n549), .A2(n411), .ZN(n550) );
  INV_X1 U459 ( .A(KEYINPUT56), .ZN(n372) );
  XOR2_X1 U460 ( .A(n487), .B(n486), .Z(n357) );
  OR2_X1 U461 ( .A1(n458), .A2(n561), .ZN(n358) );
  XOR2_X1 U462 ( .A(n480), .B(KEYINPUT107), .Z(n359) );
  AND2_X1 U463 ( .A1(n416), .A2(n534), .ZN(n360) );
  AND2_X1 U464 ( .A1(n548), .A2(n527), .ZN(n666) );
  AND2_X1 U465 ( .A1(n423), .A2(n378), .ZN(G66) );
  XNOR2_X1 U466 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n362) );
  XOR2_X1 U467 ( .A(n624), .B(KEYINPUT124), .Z(n363) );
  XOR2_X1 U468 ( .A(n635), .B(n634), .Z(n364) );
  XNOR2_X1 U469 ( .A(n710), .B(n709), .ZN(n365) );
  XNOR2_X1 U470 ( .A(KEYINPUT59), .B(n629), .ZN(n366) );
  XNOR2_X1 U471 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n367) );
  XOR2_X1 U472 ( .A(KEYINPUT115), .B(KEYINPUT63), .Z(n368) );
  AND2_X1 U473 ( .A1(n626), .A2(n351), .ZN(n720) );
  INV_X1 U474 ( .A(n720), .ZN(n378) );
  XNOR2_X1 U475 ( .A(n696), .B(KEYINPUT2), .ZN(n369) );
  BUF_X1 U476 ( .A(n632), .Z(n370) );
  XNOR2_X1 U477 ( .A(n696), .B(KEYINPUT2), .ZN(n410) );
  AND2_X2 U478 ( .A1(n410), .A2(n409), .ZN(n371) );
  AND2_X2 U479 ( .A1(n369), .A2(n409), .ZN(n715) );
  BUF_X1 U480 ( .A(n708), .Z(n710) );
  BUF_X1 U481 ( .A(n698), .Z(n726) );
  XNOR2_X1 U482 ( .A(n373), .B(n372), .ZN(G51) );
  NAND2_X1 U483 ( .A1(n380), .A2(n378), .ZN(n373) );
  XNOR2_X1 U484 ( .A(n374), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U485 ( .A1(n377), .A2(n378), .ZN(n374) );
  XNOR2_X1 U486 ( .A(n375), .B(n367), .ZN(G60) );
  NAND2_X1 U487 ( .A1(n381), .A2(n378), .ZN(n375) );
  XNOR2_X1 U488 ( .A(n376), .B(n368), .ZN(G57) );
  NAND2_X1 U489 ( .A1(n379), .A2(n378), .ZN(n376) );
  XNOR2_X1 U490 ( .A(n625), .B(n363), .ZN(n377) );
  XNOR2_X1 U491 ( .A(n636), .B(n364), .ZN(n379) );
  XNOR2_X1 U492 ( .A(n711), .B(n365), .ZN(n380) );
  XNOR2_X1 U493 ( .A(n630), .B(n366), .ZN(n381) );
  NAND2_X1 U494 ( .A1(n582), .A2(n358), .ZN(n382) );
  NAND2_X1 U495 ( .A1(n383), .A2(n571), .ZN(n572) );
  XNOR2_X1 U496 ( .A(n648), .B(KEYINPUT85), .ZN(n383) );
  NAND2_X1 U497 ( .A1(n612), .A2(n611), .ZN(n385) );
  XNOR2_X1 U498 ( .A(n386), .B(n488), .ZN(n491) );
  XNOR2_X1 U499 ( .A(n490), .B(n357), .ZN(n386) );
  NAND2_X1 U500 ( .A1(n628), .A2(n632), .ZN(n526) );
  NAND2_X1 U501 ( .A1(n355), .A2(n425), .ZN(n397) );
  XNOR2_X2 U502 ( .A(n398), .B(n422), .ZN(n628) );
  NAND2_X1 U503 ( .A1(n399), .A2(n523), .ZN(n398) );
  AND2_X2 U504 ( .A1(n551), .A2(n662), .ZN(n399) );
  NAND2_X1 U505 ( .A1(n402), .A2(n401), .ZN(n415) );
  INV_X1 U506 ( .A(n676), .ZN(n402) );
  NAND2_X1 U507 ( .A1(n403), .A2(n553), .ZN(n554) );
  XNOR2_X1 U508 ( .A(n405), .B(n404), .ZN(n403) );
  INV_X1 U509 ( .A(KEYINPUT44), .ZN(n404) );
  NAND2_X1 U510 ( .A1(n406), .A2(n408), .ZN(n405) );
  XNOR2_X1 U511 ( .A(n526), .B(n407), .ZN(n406) );
  INV_X1 U512 ( .A(n749), .ZN(n408) );
  NAND2_X2 U513 ( .A1(n698), .A2(n699), .ZN(n696) );
  XNOR2_X2 U514 ( .A(n554), .B(KEYINPUT45), .ZN(n698) );
  NAND2_X1 U515 ( .A1(n665), .A2(n666), .ZN(n528) );
  INV_X1 U516 ( .A(n665), .ZN(n411) );
  XNOR2_X2 U517 ( .A(n580), .B(n412), .ZN(n665) );
  NAND2_X1 U518 ( .A1(n413), .A2(n360), .ZN(n535) );
  NAND2_X1 U519 ( .A1(n415), .A2(n414), .ZN(n413) );
  NAND2_X1 U520 ( .A1(n676), .A2(n417), .ZN(n414) );
  XNOR2_X1 U521 ( .A(n530), .B(n529), .ZN(n676) );
  INV_X1 U522 ( .A(KEYINPUT34), .ZN(n417) );
  XNOR2_X1 U523 ( .A(n421), .B(n420), .ZN(n438) );
  XNOR2_X1 U524 ( .A(n435), .B(n434), .ZN(n420) );
  NAND2_X1 U525 ( .A1(n431), .A2(n430), .ZN(n421) );
  XNOR2_X1 U526 ( .A(n424), .B(n719), .ZN(n423) );
  NAND2_X1 U527 ( .A1(n371), .A2(G217), .ZN(n424) );
  XNOR2_X2 U528 ( .A(n437), .B(n436), .ZN(n721) );
  XNOR2_X1 U529 ( .A(n736), .B(n518), .ZN(n635) );
  XNOR2_X1 U530 ( .A(n354), .B(G134), .ZN(n499) );
  AND2_X1 U531 ( .A1(n665), .A2(n586), .ZN(n425) );
  INV_X1 U532 ( .A(KEYINPUT83), .ZN(n569) );
  NOR2_X1 U533 ( .A1(n593), .A2(n658), .ZN(n598) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U535 ( .A1(n588), .A2(n577), .ZN(n578) );
  NOR2_X1 U536 ( .A1(G902), .A2(n624), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n581), .B(KEYINPUT112), .ZN(n600) );
  XNOR2_X1 U538 ( .A(n605), .B(KEYINPUT70), .ZN(n606) );
  XNOR2_X1 U539 ( .A(n607), .B(n606), .ZN(n613) );
  INV_X1 U540 ( .A(n467), .ZN(n429) );
  INV_X1 U541 ( .A(n464), .ZN(n428) );
  NAND2_X1 U542 ( .A1(n429), .A2(n428), .ZN(n431) );
  NAND2_X1 U543 ( .A1(n467), .A2(n464), .ZN(n430) );
  INV_X2 U544 ( .A(G953), .ZN(n741) );
  NAND2_X1 U545 ( .A1(G224), .A2(n741), .ZN(n432) );
  XNOR2_X1 U546 ( .A(n438), .B(n506), .ZN(n445) );
  XNOR2_X1 U547 ( .A(G119), .B(G116), .ZN(n439) );
  XNOR2_X1 U548 ( .A(n439), .B(KEYINPUT3), .ZN(n441) );
  XNOR2_X1 U549 ( .A(n441), .B(n440), .ZN(n516) );
  INV_X1 U550 ( .A(n516), .ZN(n444) );
  XNOR2_X1 U551 ( .A(n442), .B(KEYINPUT71), .ZN(n443) );
  XNOR2_X1 U552 ( .A(n444), .B(n443), .ZN(n722) );
  XNOR2_X1 U553 ( .A(n445), .B(n722), .ZN(n708) );
  NAND2_X1 U554 ( .A1(n708), .A2(n623), .ZN(n450) );
  NAND2_X1 U555 ( .A1(n519), .A2(n446), .ZN(n451) );
  NAND2_X1 U556 ( .A1(n451), .A2(G210), .ZN(n448) );
  INV_X1 U557 ( .A(KEYINPUT80), .ZN(n447) );
  XNOR2_X1 U558 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U559 ( .A1(n451), .A2(G214), .ZN(n453) );
  INV_X1 U560 ( .A(KEYINPUT91), .ZN(n452) );
  XOR2_X1 U561 ( .A(G898), .B(KEYINPUT92), .Z(n730) );
  NAND2_X1 U562 ( .A1(n730), .A2(n351), .ZN(n455) );
  XOR2_X1 U563 ( .A(KEYINPUT93), .B(n455), .Z(n724) );
  XNOR2_X1 U564 ( .A(n456), .B(KEYINPUT14), .ZN(n457) );
  NAND2_X1 U565 ( .A1(G902), .A2(n457), .ZN(n557) );
  NOR2_X1 U566 ( .A1(n724), .A2(n557), .ZN(n458) );
  NAND2_X1 U567 ( .A1(G952), .A2(n457), .ZN(n692) );
  NOR2_X1 U568 ( .A1(n692), .A2(n351), .ZN(n561) );
  INV_X1 U569 ( .A(n531), .ZN(n481) );
  NAND2_X1 U570 ( .A1(G214), .A2(n510), .ZN(n460) );
  XOR2_X1 U571 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n463) );
  NOR2_X1 U572 ( .A1(G902), .A2(n629), .ZN(n466) );
  XNOR2_X1 U573 ( .A(KEYINPUT13), .B(KEYINPUT104), .ZN(n465) );
  NAND2_X1 U574 ( .A1(G234), .A2(n741), .ZN(n468) );
  XOR2_X1 U575 ( .A(KEYINPUT8), .B(n468), .Z(n489) );
  NAND2_X1 U576 ( .A1(G217), .A2(n489), .ZN(n472) );
  XNOR2_X1 U577 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U578 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U579 ( .A(n499), .B(n475), .ZN(n624) );
  XOR2_X1 U580 ( .A(G478), .B(n476), .Z(n538) );
  INV_X1 U581 ( .A(n538), .ZN(n533) );
  NAND2_X1 U582 ( .A1(G234), .A2(n623), .ZN(n477) );
  XNOR2_X1 U583 ( .A(KEYINPUT20), .B(n477), .ZN(n492) );
  NAND2_X1 U584 ( .A1(n492), .A2(G221), .ZN(n478) );
  XNOR2_X1 U585 ( .A(n478), .B(KEYINPUT21), .ZN(n663) );
  XOR2_X1 U586 ( .A(n663), .B(KEYINPUT98), .Z(n527) );
  INV_X1 U587 ( .A(n527), .ZN(n479) );
  NAND2_X1 U588 ( .A1(n481), .A2(n359), .ZN(n483) );
  INV_X1 U589 ( .A(KEYINPUT22), .ZN(n482) );
  XOR2_X1 U590 ( .A(G110), .B(G119), .Z(n485) );
  XNOR2_X1 U591 ( .A(n485), .B(n484), .ZN(n488) );
  XOR2_X1 U592 ( .A(KEYINPUT23), .B(KEYINPUT95), .Z(n487) );
  NAND2_X1 U593 ( .A1(G221), .A2(n489), .ZN(n490) );
  XNOR2_X1 U594 ( .A(n491), .B(n737), .ZN(n719) );
  NAND2_X1 U595 ( .A1(n719), .A2(n519), .ZN(n498) );
  XOR2_X1 U596 ( .A(KEYINPUT73), .B(KEYINPUT97), .Z(n494) );
  NAND2_X1 U597 ( .A1(n492), .A2(G217), .ZN(n493) );
  XNOR2_X1 U598 ( .A(n494), .B(n493), .ZN(n496) );
  INV_X1 U599 ( .A(KEYINPUT25), .ZN(n495) );
  XNOR2_X1 U600 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n498), .B(n497), .ZN(n662) );
  XOR2_X1 U602 ( .A(n500), .B(KEYINPUT4), .Z(n501) );
  INV_X1 U603 ( .A(KEYINPUT94), .ZN(n735) );
  NAND2_X1 U604 ( .A1(G227), .A2(n741), .ZN(n503) );
  XNOR2_X1 U605 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U606 ( .A(n505), .B(KEYINPUT75), .Z(n507) );
  NOR2_X1 U607 ( .A1(n712), .A2(G902), .ZN(n509) );
  XNOR2_X2 U608 ( .A(n509), .B(G469), .ZN(n580) );
  NAND2_X1 U609 ( .A1(n510), .A2(G210), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n512), .B(n511), .ZN(n515) );
  XNOR2_X1 U611 ( .A(n513), .B(KEYINPUT99), .ZN(n514) );
  XNOR2_X1 U612 ( .A(n515), .B(n514), .ZN(n517) );
  XNOR2_X1 U613 ( .A(n517), .B(n516), .ZN(n518) );
  NAND2_X1 U614 ( .A1(n635), .A2(n519), .ZN(n521) );
  XOR2_X1 U615 ( .A(G472), .B(KEYINPUT100), .Z(n520) );
  INV_X1 U616 ( .A(KEYINPUT108), .ZN(n522) );
  XNOR2_X1 U617 ( .A(n524), .B(n522), .ZN(n576) );
  NOR2_X1 U618 ( .A1(n665), .A2(n576), .ZN(n523) );
  INV_X1 U619 ( .A(KEYINPUT6), .ZN(n525) );
  XNOR2_X1 U620 ( .A(n669), .B(n525), .ZN(n586) );
  INV_X1 U621 ( .A(n662), .ZN(n548) );
  INV_X1 U622 ( .A(n666), .ZN(n542) );
  XNOR2_X1 U623 ( .A(n528), .B(KEYINPUT72), .ZN(n539) );
  NOR2_X1 U624 ( .A1(n586), .A2(n539), .ZN(n530) );
  XOR2_X1 U625 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n529) );
  BUF_X1 U626 ( .A(n531), .Z(n532) );
  NOR2_X1 U627 ( .A1(n537), .A2(n533), .ZN(n567) );
  XOR2_X1 U628 ( .A(n567), .B(KEYINPUT77), .Z(n534) );
  NAND2_X1 U629 ( .A1(n538), .A2(n537), .ZN(n536) );
  NOR2_X1 U630 ( .A1(n538), .A2(n537), .ZN(n649) );
  XOR2_X1 U631 ( .A(KEYINPUT84), .B(n682), .Z(n595) );
  NOR2_X1 U632 ( .A1(n539), .A2(n669), .ZN(n673) );
  INV_X1 U633 ( .A(n532), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n673), .A2(n540), .ZN(n541) );
  XOR2_X1 U635 ( .A(KEYINPUT31), .B(n541), .Z(n655) );
  OR2_X1 U636 ( .A1(n580), .A2(n542), .ZN(n562) );
  INV_X1 U637 ( .A(n562), .ZN(n543) );
  NAND2_X1 U638 ( .A1(n543), .A2(n669), .ZN(n544) );
  NOR2_X1 U639 ( .A1(n532), .A2(n544), .ZN(n545) );
  XNOR2_X1 U640 ( .A(KEYINPUT101), .B(n545), .ZN(n640) );
  NAND2_X1 U641 ( .A1(n655), .A2(n640), .ZN(n546) );
  NAND2_X1 U642 ( .A1(n595), .A2(n546), .ZN(n547) );
  XOR2_X1 U643 ( .A(KEYINPUT106), .B(n547), .Z(n552) );
  AND2_X1 U644 ( .A1(n586), .A2(n548), .ZN(n549) );
  AND2_X1 U645 ( .A1(n551), .A2(n550), .ZN(n637) );
  NOR2_X1 U646 ( .A1(n552), .A2(n637), .ZN(n553) );
  NAND2_X1 U647 ( .A1(n576), .A2(n677), .ZN(n556) );
  XNOR2_X1 U648 ( .A(KEYINPUT30), .B(KEYINPUT111), .ZN(n555) );
  XNOR2_X1 U649 ( .A(n556), .B(n555), .ZN(n564) );
  NOR2_X1 U650 ( .A1(G900), .A2(n557), .ZN(n558) );
  NAND2_X1 U651 ( .A1(n351), .A2(n558), .ZN(n559) );
  XOR2_X1 U652 ( .A(KEYINPUT110), .B(n559), .Z(n560) );
  NOR2_X1 U653 ( .A1(n561), .A2(n560), .ZN(n573) );
  NOR2_X1 U654 ( .A1(n573), .A2(n562), .ZN(n563) );
  NAND2_X1 U655 ( .A1(n564), .A2(n563), .ZN(n604) );
  BUF_X1 U656 ( .A(n565), .Z(n566) );
  NAND2_X1 U657 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U658 ( .A1(KEYINPUT47), .A2(n682), .ZN(n570) );
  XNOR2_X1 U659 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U660 ( .A(n572), .B(KEYINPUT81), .ZN(n584) );
  NOR2_X1 U661 ( .A1(n663), .A2(n573), .ZN(n574) );
  XOR2_X1 U662 ( .A(KEYINPUT67), .B(n574), .Z(n575) );
  NAND2_X1 U663 ( .A1(n662), .A2(n575), .ZN(n588) );
  INV_X1 U664 ( .A(n576), .ZN(n577) );
  XOR2_X1 U665 ( .A(KEYINPUT28), .B(n578), .Z(n579) );
  NOR2_X1 U666 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U667 ( .A1(n600), .A2(n356), .ZN(n594) );
  NAND2_X1 U668 ( .A1(n594), .A2(KEYINPUT47), .ZN(n583) );
  NAND2_X1 U669 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U670 ( .A(KEYINPUT82), .B(n585), .ZN(n593) );
  INV_X1 U671 ( .A(n586), .ZN(n587) );
  NAND2_X1 U672 ( .A1(n649), .A2(n587), .ZN(n589) );
  NOR2_X1 U673 ( .A1(n589), .A2(n588), .ZN(n614) );
  NAND2_X1 U674 ( .A1(n614), .A2(n353), .ZN(n591) );
  XNOR2_X1 U675 ( .A(n591), .B(KEYINPUT36), .ZN(n592) );
  INV_X1 U676 ( .A(n594), .ZN(n650) );
  NAND2_X1 U677 ( .A1(n650), .A2(n595), .ZN(n596) );
  OR2_X1 U678 ( .A1(KEYINPUT47), .A2(n596), .ZN(n597) );
  AND2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n612) );
  XNOR2_X1 U680 ( .A(n566), .B(KEYINPUT38), .ZN(n603) );
  INV_X1 U681 ( .A(n603), .ZN(n678) );
  NAND2_X1 U682 ( .A1(n678), .A2(n677), .ZN(n681) );
  NOR2_X1 U683 ( .A1(n681), .A2(n680), .ZN(n599) );
  XNOR2_X1 U684 ( .A(KEYINPUT41), .B(n599), .ZN(n693) );
  INV_X1 U685 ( .A(n600), .ZN(n601) );
  NOR2_X1 U686 ( .A1(n693), .A2(n601), .ZN(n602) );
  XNOR2_X1 U687 ( .A(n602), .B(KEYINPUT42), .ZN(n751) );
  NOR2_X1 U688 ( .A1(n604), .A2(n603), .ZN(n607) );
  XNOR2_X1 U689 ( .A(KEYINPUT87), .B(KEYINPUT39), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n649), .A2(n613), .ZN(n609) );
  XNOR2_X1 U691 ( .A(KEYINPUT113), .B(KEYINPUT40), .ZN(n608) );
  XNOR2_X1 U692 ( .A(n609), .B(n608), .ZN(n750) );
  XNOR2_X1 U693 ( .A(n610), .B(KEYINPUT46), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n645), .A2(n613), .ZN(n661) );
  INV_X1 U695 ( .A(n677), .ZN(n616) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U697 ( .A(n617), .B(KEYINPUT43), .Z(n619) );
  INV_X1 U698 ( .A(n566), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n627) );
  AND2_X1 U700 ( .A1(n661), .A2(n627), .ZN(n620) );
  INV_X1 U701 ( .A(KEYINPUT2), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n371), .A2(G478), .ZN(n625) );
  INV_X1 U703 ( .A(G952), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n627), .B(G140), .ZN(G42) );
  XNOR2_X1 U705 ( .A(n628), .B(G110), .ZN(G12) );
  NAND2_X1 U706 ( .A1(n715), .A2(G475), .ZN(n630) );
  XOR2_X1 U707 ( .A(G119), .B(KEYINPUT127), .Z(n631) );
  XNOR2_X1 U708 ( .A(n370), .B(n631), .ZN(G21) );
  NAND2_X1 U709 ( .A1(n715), .A2(G472), .ZN(n636) );
  XOR2_X1 U710 ( .A(KEYINPUT90), .B(KEYINPUT114), .Z(n633) );
  XNOR2_X1 U711 ( .A(n633), .B(KEYINPUT62), .ZN(n634) );
  XOR2_X1 U712 ( .A(G101), .B(n637), .Z(G3) );
  INV_X1 U713 ( .A(n649), .ZN(n652) );
  NOR2_X1 U714 ( .A1(n652), .A2(n640), .ZN(n638) );
  XOR2_X1 U715 ( .A(G104), .B(n638), .Z(n639) );
  XNOR2_X1 U716 ( .A(KEYINPUT116), .B(n639), .ZN(G6) );
  INV_X1 U717 ( .A(n645), .ZN(n656) );
  NOR2_X1 U718 ( .A1(n640), .A2(n656), .ZN(n644) );
  XOR2_X1 U719 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n642) );
  XNOR2_X1 U720 ( .A(G107), .B(KEYINPUT26), .ZN(n641) );
  XNOR2_X1 U721 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n644), .B(n643), .ZN(G9) );
  XOR2_X1 U723 ( .A(G128), .B(KEYINPUT29), .Z(n647) );
  NAND2_X1 U724 ( .A1(n650), .A2(n645), .ZN(n646) );
  XNOR2_X1 U725 ( .A(n647), .B(n646), .ZN(G30) );
  XOR2_X1 U726 ( .A(G143), .B(n648), .Z(G45) );
  NAND2_X1 U727 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n651), .B(G146), .ZN(G48) );
  NOR2_X1 U729 ( .A1(n652), .A2(n655), .ZN(n653) );
  XOR2_X1 U730 ( .A(KEYINPUT118), .B(n653), .Z(n654) );
  XNOR2_X1 U731 ( .A(G113), .B(n654), .ZN(G15) );
  NOR2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U733 ( .A(G116), .B(n657), .Z(G18) );
  XOR2_X1 U734 ( .A(KEYINPUT119), .B(KEYINPUT37), .Z(n660) );
  XNOR2_X1 U735 ( .A(G125), .B(n658), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n660), .B(n659), .ZN(G27) );
  XNOR2_X1 U737 ( .A(G134), .B(n661), .ZN(G36) );
  NAND2_X1 U738 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n664), .B(KEYINPUT49), .ZN(n671) );
  NOR2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U741 ( .A(KEYINPUT50), .B(n667), .Z(n668) );
  NAND2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U745 ( .A(KEYINPUT51), .B(n674), .Z(n675) );
  NOR2_X1 U746 ( .A1(n693), .A2(n675), .ZN(n689) );
  NOR2_X1 U747 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n685), .B(KEYINPUT120), .ZN(n686) );
  NOR2_X1 U752 ( .A1(n676), .A2(n686), .ZN(n687) );
  XOR2_X1 U753 ( .A(KEYINPUT121), .B(n687), .Z(n688) );
  NOR2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n690), .B(KEYINPUT52), .ZN(n691) );
  NOR2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U757 ( .A1(n676), .A2(n693), .ZN(n694) );
  NOR2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n705) );
  NAND2_X1 U759 ( .A1(n352), .A2(KEYINPUT86), .ZN(n697) );
  NAND2_X1 U760 ( .A1(n697), .A2(KEYINPUT2), .ZN(n703) );
  XNOR2_X1 U761 ( .A(n739), .B(KEYINPUT86), .ZN(n700) );
  NAND2_X1 U762 ( .A1(n726), .A2(n700), .ZN(n701) );
  NAND2_X1 U763 ( .A1(n701), .A2(n622), .ZN(n702) );
  NAND2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U765 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U766 ( .A1(n706), .A2(n351), .ZN(n707) );
  XNOR2_X1 U767 ( .A(n707), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U768 ( .A1(n715), .A2(G210), .ZN(n711) );
  XOR2_X1 U769 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n709) );
  XNOR2_X1 U770 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n714) );
  XNOR2_X1 U771 ( .A(n712), .B(KEYINPUT57), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n714), .B(n713), .ZN(n717) );
  NAND2_X1 U773 ( .A1(n371), .A2(G469), .ZN(n716) );
  XOR2_X1 U774 ( .A(n717), .B(n716), .Z(n718) );
  NOR2_X1 U775 ( .A1(n720), .A2(n718), .ZN(G54) );
  XOR2_X1 U776 ( .A(n721), .B(G101), .Z(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n725), .A2(n724), .ZN(n734) );
  INV_X1 U779 ( .A(n726), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n727), .A2(n351), .ZN(n732) );
  NAND2_X1 U781 ( .A1(n351), .A2(G224), .ZN(n728) );
  XOR2_X1 U782 ( .A(KEYINPUT61), .B(n728), .Z(n729) );
  NOR2_X1 U783 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n734), .B(n733), .ZN(G69) );
  XNOR2_X1 U786 ( .A(n736), .B(n735), .ZN(n738) );
  XOR2_X1 U787 ( .A(n738), .B(n737), .Z(n743) );
  INV_X1 U788 ( .A(n743), .ZN(n740) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n748) );
  XNOR2_X1 U791 ( .A(G227), .B(n743), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n744), .A2(G900), .ZN(n745) );
  XNOR2_X1 U793 ( .A(KEYINPUT126), .B(n745), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(n351), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U796 ( .A(n749), .B(G122), .Z(G24) );
  XOR2_X1 U797 ( .A(G131), .B(n750), .Z(G33) );
  XOR2_X1 U798 ( .A(G137), .B(n751), .Z(G39) );
endmodule

