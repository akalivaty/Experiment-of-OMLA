//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  XOR2_X1   g006(.A(new_n206), .B(new_n207), .Z(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n209), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT25), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT23), .B1(new_n218), .B2(KEYINPUT64), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n220), .B(new_n221), .C1(G169gat), .C2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n211), .A2(new_n225), .A3(new_n212), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n217), .A2(new_n224), .B1(new_n227), .B2(KEYINPUT25), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT27), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT27), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G183gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT28), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n233), .A2(new_n234), .A3(G190gat), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT66), .B1(new_n230), .B2(new_n232), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT66), .B1(new_n231), .B2(G183gat), .ZN(new_n237));
  INV_X1    g036(.A(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n234), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT67), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n242), .B(new_n234), .C1(new_n236), .C2(new_n239), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n235), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT26), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n218), .B1(new_n245), .B2(new_n223), .ZN(new_n246));
  NOR3_X1   g045(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n209), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n228), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT72), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n228), .B(KEYINPUT72), .C1(new_n244), .C2(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n249), .A2(new_n257), .A3(new_n254), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n208), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G8gat), .B(G36gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n251), .A2(new_n257), .A3(new_n252), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n254), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n263), .A2(KEYINPUT73), .A3(new_n254), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n255), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT74), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT74), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n270), .A3(new_n255), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  AOI211_X1 g072(.A(new_n259), .B(new_n262), .C1(new_n273), .C2(new_n208), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT30), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n208), .ZN(new_n276));
  INV_X1    g075(.A(new_n259), .ZN(new_n277));
  INV_X1    g076(.A(new_n262), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT30), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n263), .A2(KEYINPUT73), .A3(new_n254), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT73), .B1(new_n263), .B2(new_n254), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n269), .A2(new_n271), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n208), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n277), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT75), .B1(new_n287), .B2(new_n262), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n259), .B1(new_n273), .B2(new_n208), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n289), .A2(new_n290), .A3(new_n278), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n275), .B(new_n281), .C1(new_n288), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT84), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(new_n289), .B2(new_n278), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n283), .A2(new_n284), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n286), .B1(new_n295), .B2(new_n267), .ZN(new_n296));
  OAI211_X1 g095(.A(KEYINPUT75), .B(new_n262), .C1(new_n296), .C2(new_n259), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n294), .A2(new_n297), .B1(KEYINPUT30), .B2(new_n274), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT84), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(new_n281), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G1gat), .B(G29gat), .Z(new_n302));
  XNOR2_X1  g101(.A(G57gat), .B(G85gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G120gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(G120gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(KEYINPUT69), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(KEYINPUT69), .B2(new_n308), .ZN(new_n311));
  XOR2_X1   g110(.A(G127gat), .B(G134gat), .Z(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT1), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G120gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G113gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(new_n308), .A3(KEYINPUT68), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT68), .B1(new_n316), .B2(new_n308), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n312), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G155gat), .B(G162gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G155gat), .ZN(new_n326));
  INV_X1    g125(.A(G162gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT2), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G141gat), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(G148gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n330), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT78), .B(G148gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(new_n331), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n323), .A2(new_n328), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n325), .A2(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n325), .A2(new_n333), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n336), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n314), .A2(new_n321), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT39), .B1(new_n348), .B2(KEYINPUT85), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(KEYINPUT85), .B2(new_n348), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n322), .B2(new_n338), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n322), .A2(new_n351), .A3(new_n338), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n352), .A2(new_n353), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n340), .B2(new_n341), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT79), .B1(new_n338), .B2(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n338), .A2(new_n358), .ZN(new_n363));
  AND4_X1   g162(.A1(new_n361), .A2(new_n362), .A3(new_n343), .A4(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n347), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n306), .B1(new_n350), .B2(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n365), .A2(KEYINPUT39), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(KEYINPUT40), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT86), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT40), .B1(new_n366), .B2(new_n367), .ZN(new_n370));
  INV_X1    g169(.A(new_n306), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n361), .A2(new_n362), .A3(new_n343), .A4(new_n363), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n347), .A2(KEYINPUT5), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n372), .B(new_n373), .C1(new_n355), .C2(new_n356), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT5), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(new_n345), .B2(new_n347), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT4), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n346), .B1(new_n377), .B2(new_n352), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n364), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n371), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n370), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n369), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n301), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT37), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n276), .A2(new_n385), .A3(new_n277), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n262), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n289), .A2(new_n385), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT38), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n273), .A2(new_n286), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n256), .A2(new_n258), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n385), .B1(new_n391), .B2(new_n208), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT38), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(new_n262), .A3(new_n386), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n374), .A2(new_n379), .A3(new_n371), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n397), .A2(new_n380), .A3(KEYINPUT6), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n399));
  AOI211_X1 g198(.A(new_n399), .B(new_n371), .C1(new_n374), .C2(new_n379), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n279), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n393), .A2(new_n386), .A3(KEYINPUT87), .A4(new_n262), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n396), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT3), .B1(new_n286), .B2(new_n257), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n338), .B2(new_n358), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n406), .A2(new_n338), .B1(new_n286), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G50gat), .ZN(new_n413));
  XOR2_X1   g212(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  MUX2_X1   g214(.A(new_n411), .B(G22gat), .S(new_n415), .Z(new_n416));
  XNOR2_X1  g215(.A(new_n410), .B(new_n416), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n405), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n384), .A2(new_n418), .A3(KEYINPUT88), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n382), .B1(new_n293), .B2(new_n300), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n417), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n417), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n401), .B1(new_n280), .B2(new_n279), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n298), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n294), .A2(new_n297), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n428), .A2(new_n426), .A3(new_n275), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n424), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G15gat), .B(G43gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n249), .B(new_n322), .ZN(new_n434));
  INV_X1    g233(.A(G227gat), .ZN(new_n435));
  INV_X1    g234(.A(G233gat), .ZN(new_n436));
  OR3_X1    g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n438));
  AOI21_X1  g237(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(KEYINPUT32), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n437), .B(KEYINPUT32), .C1(new_n438), .C2(new_n433), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n444));
  XOR2_X1   g243(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(new_n446), .A3(new_n442), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT36), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n430), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n419), .A2(new_n423), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n301), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n449), .A3(new_n417), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n456), .A2(KEYINPUT35), .A3(new_n401), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n298), .A2(new_n426), .ZN(new_n459));
  INV_X1    g258(.A(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n298), .A2(new_n426), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .A4(new_n425), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n454), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT18), .ZN(new_n466));
  INV_X1    g265(.A(G29gat), .ZN(new_n467));
  INV_X1    g266(.A(G36gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(KEYINPUT14), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT89), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT89), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(KEYINPUT14), .B2(new_n469), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n471), .A2(new_n474), .B1(G29gat), .B2(G36gat), .ZN(new_n475));
  INV_X1    g274(.A(G50gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G43gat), .ZN(new_n477));
  INV_X1    g276(.A(G43gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G50gat), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT15), .ZN(new_n480));
  INV_X1    g279(.A(new_n472), .ZN(new_n481));
  OAI221_X1 g280(.A(new_n480), .B1(new_n467), .B2(new_n468), .C1(new_n470), .C2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT90), .B(G50gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n478), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT15), .B1(new_n484), .B2(new_n477), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n475), .A2(new_n480), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT17), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT16), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(G1gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(KEYINPUT92), .C1(G1gat), .C2(new_n491), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(G8gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT93), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n486), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(KEYINPUT95), .B(new_n466), .C1(new_n502), .C2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n495), .A2(new_n486), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT96), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n501), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n503), .B(KEYINPUT13), .Z(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT95), .B1(new_n502), .B2(new_n504), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT18), .ZN(new_n514));
  XOR2_X1   g313(.A(G113gat), .B(G141gat), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT11), .ZN(new_n516));
  INV_X1    g315(.A(G169gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G197gat), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n519), .B(KEYINPUT12), .Z(new_n520));
  NAND3_X1  g319(.A1(new_n512), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT97), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n512), .A2(KEYINPUT97), .A3(new_n514), .A4(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n512), .A2(new_n514), .ZN(new_n526));
  INV_X1    g325(.A(new_n520), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT10), .ZN(new_n530));
  XNOR2_X1  g329(.A(G57gat), .B(G64gat), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(G71gat), .B(G78gat), .Z(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G99gat), .B(G106gat), .Z(new_n538));
  NAND2_X1  g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  INV_X1    g341(.A(G85gat), .ZN(new_n543));
  INV_X1    g342(.A(G92gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(KEYINPUT8), .A2(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n537), .B1(new_n538), .B2(new_n546), .ZN(new_n547));
  OR3_X1    g346(.A1(new_n546), .A2(KEYINPUT101), .A3(new_n538), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT101), .B1(new_n546), .B2(new_n538), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT102), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n548), .A2(KEYINPUT102), .A3(new_n549), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n553), .A2(new_n554), .B1(new_n538), .B2(new_n546), .ZN(new_n555));
  INV_X1    g354(.A(new_n537), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n530), .B(new_n551), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n554), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT10), .A3(new_n547), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n563));
  INV_X1    g362(.A(new_n561), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n565), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n564), .B1(new_n557), .B2(new_n559), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n529), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n555), .A2(new_n486), .B1(KEYINPUT41), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n546), .A2(new_n538), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n490), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT103), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT103), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n586), .A3(new_n583), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n582), .A2(new_n583), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n577), .A2(KEYINPUT41), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT99), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n585), .A2(new_n588), .A3(new_n587), .A4(new_n590), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n594), .B1(new_n592), .B2(new_n595), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n556), .A2(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT98), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n603), .B(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n495), .B1(KEYINPUT21), .B2(new_n556), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n576), .A2(new_n598), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n465), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n401), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G1gat), .ZN(G1324gat));
  INV_X1    g413(.A(new_n612), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n455), .ZN(new_n616));
  INV_X1    g415(.A(G8gat), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT42), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT16), .B(G8gat), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  MUX2_X1   g419(.A(KEYINPUT42), .B(new_n618), .S(new_n620), .Z(G1325gat));
  OR3_X1    g420(.A1(new_n615), .A2(G15gat), .A3(new_n450), .ZN(new_n622));
  OAI21_X1  g421(.A(G15gat), .B1(new_n615), .B2(new_n452), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(G1326gat));
  NAND2_X1  g423(.A1(new_n612), .A2(new_n424), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT43), .B(G22gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(G1327gat));
  AOI22_X1  g426(.A1(new_n455), .A2(new_n457), .B1(new_n462), .B2(KEYINPUT35), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n430), .A2(new_n452), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n421), .A2(new_n422), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(KEYINPUT88), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n628), .B1(new_n631), .B2(new_n423), .ZN(new_n632));
  INV_X1    g431(.A(new_n598), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n610), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(new_n576), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(new_n467), .A3(new_n401), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT45), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n632), .B2(new_n633), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n465), .A2(KEYINPUT44), .A3(new_n598), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n636), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n398), .A2(new_n400), .ZN(new_n645));
  OAI21_X1  g444(.A(G29gat), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n639), .A2(new_n646), .ZN(G1328gat));
  OAI21_X1  g446(.A(G36gat), .B1(new_n644), .B2(new_n455), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n637), .A2(new_n468), .A3(new_n301), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n651), .A2(KEYINPUT46), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT46), .B1(new_n651), .B2(new_n652), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n648), .B1(new_n653), .B2(new_n654), .ZN(G1329gat));
  INV_X1    g454(.A(new_n450), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n478), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n450), .B(KEYINPUT36), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n641), .A2(new_n658), .A3(new_n636), .A4(new_n642), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(G43gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(new_n660), .A3(KEYINPUT47), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n659), .A2(KEYINPUT105), .A3(G43gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n657), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT105), .B1(new_n659), .B2(G43gat), .ZN(new_n665));
  OAI211_X1 g464(.A(KEYINPUT106), .B(new_n662), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(new_n663), .A3(new_n657), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT106), .B1(new_n670), .B2(new_n662), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n661), .B1(new_n667), .B2(new_n671), .ZN(G1330gat));
  OAI21_X1  g471(.A(new_n483), .B1(new_n644), .B2(new_n417), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT48), .B1(new_n673), .B2(KEYINPUT107), .ZN(new_n674));
  INV_X1    g473(.A(new_n483), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n637), .A2(new_n424), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n673), .B(new_n676), .C1(KEYINPUT107), .C2(KEYINPUT48), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(G1331gat));
  AOI22_X1  g479(.A1(new_n523), .A2(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n635), .A2(new_n633), .A3(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n632), .A2(new_n575), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n401), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n301), .ZN(new_n686));
  NOR2_X1   g485(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n687));
  AND2_X1   g486(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n687), .B2(new_n686), .ZN(G1333gat));
  AOI21_X1  g489(.A(G71gat), .B1(new_n683), .B2(new_n656), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n658), .A2(G71gat), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n683), .B2(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g493(.A1(new_n683), .A2(new_n424), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g495(.A1(new_n635), .A2(new_n529), .A3(new_n575), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n643), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT108), .B1(new_n698), .B2(new_n645), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G85gat), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n698), .A2(KEYINPUT108), .A3(new_n645), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n635), .A2(new_n529), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n634), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT51), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n634), .A2(KEYINPUT51), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n574), .A2(new_n401), .A3(new_n543), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT109), .ZN(new_n710));
  OAI22_X1  g509(.A1(new_n700), .A2(new_n701), .B1(new_n708), .B2(new_n710), .ZN(G1336gat));
  NAND3_X1  g510(.A1(new_n301), .A2(new_n544), .A3(new_n574), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT111), .Z(new_n713));
  INV_X1    g512(.A(new_n706), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT51), .B1(new_n634), .B2(new_n702), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT112), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n643), .A2(new_n301), .A3(new_n697), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(KEYINPUT110), .A3(G92gat), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n707), .A2(new_n720), .A3(new_n713), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n717), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n718), .A2(G92gat), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(KEYINPUT110), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n716), .B2(new_n723), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n726), .ZN(G1337gat));
  OAI21_X1  g526(.A(G99gat), .B1(new_n698), .B2(new_n452), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n450), .A2(G99gat), .A3(new_n575), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n708), .B2(new_n729), .ZN(G1338gat));
  NOR3_X1   g529(.A1(new_n575), .A2(G106gat), .A3(new_n417), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT113), .B1(new_n707), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G106gat), .B1(new_n698), .B2(new_n417), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g534(.A1(new_n557), .A2(new_n559), .A3(new_n564), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n562), .A2(KEYINPUT54), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT114), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n562), .A2(new_n739), .A3(KEYINPUT54), .A4(new_n736), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT54), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n569), .B1(new_n572), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n738), .A2(KEYINPUT55), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n570), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n740), .A2(new_n742), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT55), .B1(new_n746), .B2(new_n738), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n529), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n509), .A2(new_n510), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n502), .A2(new_n504), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n519), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n752), .A2(KEYINPUT115), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(KEYINPUT115), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n523), .A2(new_n524), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n574), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n598), .B1(new_n749), .B2(new_n756), .ZN(new_n757));
  AND4_X1   g556(.A1(new_n598), .A2(new_n755), .A3(new_n745), .A4(new_n748), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n681), .A2(new_n744), .A3(new_n747), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n755), .A2(new_n574), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n633), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n598), .A2(new_n755), .A3(new_n745), .A4(new_n748), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT116), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n610), .B1(new_n760), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n682), .A2(new_n574), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n301), .A2(new_n645), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n460), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n681), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n307), .ZN(G1340gat));
  NOR2_X1   g573(.A1(new_n772), .A2(new_n575), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(new_n315), .ZN(G1341gat));
  NOR2_X1   g575(.A1(new_n772), .A2(new_n610), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT117), .A2(G127gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1342gat));
  NAND2_X1  g578(.A1(new_n771), .A2(new_n598), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782));
  INV_X1    g581(.A(G134gat), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n781), .B(new_n460), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1343gat));
  NOR2_X1   g585(.A1(new_n658), .A2(new_n417), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n788), .A2(G141gat), .A3(new_n681), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n763), .A2(KEYINPUT119), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n757), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n792), .A3(new_n764), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n767), .B1(new_n793), .B2(new_n610), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT57), .B1(new_n794), .B2(new_n417), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n763), .A2(KEYINPUT116), .A3(new_n764), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n635), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n797), .B(new_n424), .C1(new_n800), .C2(new_n767), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n770), .A2(new_n452), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT118), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT120), .B1(new_n796), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n795), .A2(new_n806), .A3(new_n801), .A4(new_n803), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n807), .A3(new_n529), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n789), .B1(new_n808), .B2(G141gat), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n789), .A2(KEYINPUT58), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n804), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n331), .B1(new_n812), .B2(new_n529), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n813), .ZN(G1344gat));
  NOR3_X1   g613(.A1(new_n788), .A2(new_n335), .A3(new_n575), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n635), .B1(new_n763), .B2(new_n764), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n424), .B1(new_n767), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n797), .ZN(new_n818));
  OAI211_X1 g617(.A(KEYINPUT57), .B(new_n424), .C1(new_n800), .C2(new_n767), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n574), .A3(new_n803), .ZN(new_n824));
  AND2_X1   g623(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n815), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n805), .A2(new_n807), .A3(new_n574), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n335), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n828), .B2(KEYINPUT59), .ZN(G1345gat));
  AND3_X1   g628(.A1(new_n805), .A2(new_n635), .A3(new_n807), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n635), .A2(new_n326), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n830), .A2(new_n326), .B1(new_n788), .B2(new_n831), .ZN(G1346gat));
  NAND3_X1  g631(.A1(new_n805), .A2(new_n807), .A3(new_n598), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT122), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n805), .A2(new_n807), .A3(new_n835), .A4(new_n598), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(G162gat), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n781), .A2(new_n327), .A3(new_n787), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1347gat));
  NAND2_X1  g638(.A1(new_n301), .A2(new_n645), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT123), .Z(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n656), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n842), .A2(KEYINPUT124), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(KEYINPUT124), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n843), .A2(new_n417), .A3(new_n769), .A4(new_n844), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n517), .A3(new_n681), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n401), .B1(new_n766), .B2(new_n768), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n455), .A2(new_n456), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(G169gat), .B1(new_n850), .B2(new_n529), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n846), .A2(new_n851), .ZN(G1348gat));
  OAI21_X1  g651(.A(G176gat), .B1(new_n845), .B2(new_n575), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n575), .A2(G176gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n849), .B2(new_n854), .ZN(G1349gat));
  NOR2_X1   g654(.A1(new_n610), .A2(new_n233), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT125), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(G183gat), .B1(new_n845), .B2(new_n610), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g659(.A1(new_n849), .A2(G190gat), .A3(new_n633), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT126), .ZN(new_n862));
  OAI21_X1  g661(.A(G190gat), .B1(new_n845), .B2(new_n633), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(G1351gat));
  NAND4_X1  g666(.A1(new_n769), .A2(new_n645), .A3(new_n301), .A4(new_n787), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(G197gat), .B1(new_n869), .B2(new_n529), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n841), .A2(new_n452), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n769), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n424), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n819), .A2(new_n820), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n871), .B1(new_n874), .B2(new_n818), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n529), .A2(G197gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n870), .B1(new_n875), .B2(new_n876), .ZN(G1352gat));
  NOR3_X1   g676(.A1(new_n868), .A2(G204gat), .A3(new_n575), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT62), .ZN(new_n879));
  INV_X1    g678(.A(G204gat), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n575), .B(new_n871), .C1(new_n874), .C2(new_n818), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(G1353gat));
  NAND3_X1  g681(.A1(new_n869), .A2(new_n203), .A3(new_n635), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT63), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n884), .B(new_n203), .C1(new_n875), .C2(new_n635), .ZN(new_n885));
  INV_X1    g684(.A(new_n871), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n823), .A2(new_n635), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT63), .B1(new_n887), .B2(G211gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n883), .B1(new_n885), .B2(new_n888), .ZN(G1354gat));
  NAND3_X1  g688(.A1(new_n869), .A2(new_n204), .A3(new_n598), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n875), .A2(new_n598), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n204), .ZN(G1355gat));
endmodule


