//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT2), .B(G113), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT69), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT69), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n194), .A3(G116), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(KEYINPUT70), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT70), .B1(new_n195), .B2(new_n197), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n190), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(new_n197), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(new_n190), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  AOI21_X1  g027(.A(G146), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n206), .B(new_n209), .C1(new_n214), .C2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(G146), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(new_n213), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n207), .B(new_n219), .C1(new_n220), .C2(new_n215), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n216), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT64), .B(G143), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(G146), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n206), .B1(new_n225), .B2(new_n209), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G134), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G137), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(KEYINPUT11), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(G134), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT66), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(KEYINPUT66), .B(new_n234), .C1(new_n230), .C2(G137), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n232), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G131), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n230), .A2(G137), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n233), .B2(new_n234), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n231), .B2(KEYINPUT11), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n241), .B1(new_n243), .B2(new_n236), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT68), .B(G128), .Z(new_n248));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n218), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n225), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n218), .B1(new_n224), .B2(G146), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n245), .B1(new_n233), .B2(new_n240), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(new_n244), .B2(new_n245), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n227), .A2(new_n247), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT30), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n258), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n238), .A2(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n243), .A2(new_n236), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n245), .B1(new_n265), .B2(new_n232), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n216), .B1(new_n220), .B2(new_n215), .ZN(new_n268));
  INV_X1    g082(.A(new_n209), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT65), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n221), .A3(new_n217), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n263), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n227), .A2(KEYINPUT67), .A3(new_n247), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n262), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n205), .B(new_n260), .C1(new_n274), .C2(KEYINPUT30), .ZN(new_n275));
  INV_X1    g089(.A(new_n205), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n227), .A2(new_n247), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n276), .A2(new_n277), .A3(new_n261), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G237), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G210), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n282), .B(KEYINPUT27), .Z(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G101), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n283), .B(new_n284), .Z(new_n285));
  NAND3_X1  g099(.A1(new_n275), .A2(new_n279), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n275), .A2(KEYINPUT31), .A3(new_n279), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n276), .B1(new_n259), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n277), .A2(new_n292), .A3(new_n261), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n267), .A2(new_n271), .A3(new_n263), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT67), .B1(new_n227), .B2(new_n247), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n261), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n278), .B1(new_n299), .B2(new_n205), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n296), .B1(new_n300), .B2(new_n291), .ZN(new_n301));
  INV_X1    g115(.A(new_n285), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n189), .B1(new_n290), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT32), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT32), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n288), .A2(new_n289), .B1(new_n301), .B2(new_n302), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(new_n189), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n301), .A2(new_n285), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n275), .A2(new_n279), .A3(new_n302), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT29), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n259), .A2(new_n276), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT28), .B1(new_n278), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n285), .A2(KEYINPUT29), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n296), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n296), .A2(new_n313), .A3(KEYINPUT72), .A4(new_n314), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n188), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G472), .B1(new_n311), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n305), .A2(new_n308), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT90), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(G146), .B(new_n325), .C1(new_n329), .C2(new_n323), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(KEYINPUT19), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n280), .A2(new_n281), .A3(G214), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n224), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n280), .A2(new_n281), .A3(G143), .A4(G214), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G131), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n245), .B1(new_n333), .B2(new_n334), .ZN(new_n337));
  OAI221_X1 g151(.A(new_n330), .B1(new_n331), .B2(G146), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n326), .A2(new_n328), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n215), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n329), .A2(G146), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT18), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(new_n245), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n335), .A2(G131), .ZN(new_n345));
  OAI221_X1 g159(.A(new_n342), .B1(new_n335), .B2(new_n344), .C1(new_n345), .C2(new_n343), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n338), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT89), .ZN(new_n348));
  XNOR2_X1  g162(.A(G113), .B(G122), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n347), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n336), .A2(KEYINPUT17), .A3(new_n337), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n325), .B1(new_n329), .B2(new_n323), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n215), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT17), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n356), .B(new_n330), .C1(new_n345), .C2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n346), .B(new_n351), .C1(new_n354), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n348), .B1(new_n347), .B2(new_n352), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n322), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(G475), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n347), .A2(new_n352), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT89), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n365), .A2(KEYINPUT90), .A3(new_n359), .A4(new_n353), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(new_n359), .A3(new_n353), .ZN(new_n368));
  NOR3_X1   g182(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n367), .A2(KEYINPUT20), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n248), .A2(G143), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n224), .A2(G128), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G134), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n230), .A3(new_n372), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G107), .ZN(new_n377));
  INV_X1    g191(.A(G122), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G116), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n379), .B2(KEYINPUT14), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n196), .A2(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n382), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT9), .B(G234), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n388), .A2(new_n389), .A3(G953), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n372), .A2(new_n392), .B1(new_n248), .B2(G143), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n224), .A2(KEYINPUT13), .A3(G128), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n230), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n382), .B(G107), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n375), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n387), .B(new_n391), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n395), .A2(new_n397), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n385), .B1(new_n374), .B2(new_n375), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n390), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n188), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G478), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT15), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n402), .B(new_n404), .Z(new_n405));
  NAND2_X1  g219(.A1(G234), .A2(G237), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(G952), .A3(new_n281), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n407), .B(KEYINPUT91), .Z(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT21), .B(G898), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(G902), .A3(G953), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n408), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n354), .A2(new_n358), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n351), .B1(new_n414), .B2(new_n346), .ZN(new_n415));
  INV_X1    g229(.A(new_n359), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n188), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G475), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n370), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n389), .B1(G234), .B2(new_n188), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT75), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT23), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT69), .B(G119), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G128), .ZN(new_n425));
  OR2_X1    g239(.A1(KEYINPUT68), .A2(G128), .ZN(new_n426));
  NAND2_X1  g240(.A1(KEYINPUT68), .A2(G128), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(G119), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n423), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n192), .A2(new_n194), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT23), .B1(new_n430), .B2(new_n253), .ZN(new_n431));
  OAI21_X1  g245(.A(G110), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n356), .A2(new_n330), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n248), .A2(G119), .B1(new_n424), .B2(G128), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT24), .B(G110), .Z(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n330), .A2(new_n340), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n434), .A2(new_n435), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n431), .ZN(new_n442));
  INV_X1    g256(.A(G110), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n442), .B(new_n443), .C1(new_n434), .C2(new_n423), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n439), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n422), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n429), .A2(G110), .A3(new_n431), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n340), .B(new_n330), .C1(new_n447), .C2(new_n440), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT75), .A3(new_n437), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT22), .B(G137), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n446), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n448), .A2(KEYINPUT75), .A3(new_n437), .A4(new_n454), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT25), .B1(new_n458), .B2(new_n188), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT25), .ZN(new_n460));
  AOI211_X1 g274(.A(new_n460), .B(G902), .C1(new_n456), .C2(new_n457), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n421), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT76), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT76), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n464), .B(new_n421), .C1(new_n459), .C2(new_n461), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n421), .A2(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n463), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n321), .A2(new_n420), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(G221), .B1(new_n388), .B2(G902), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n471), .B(KEYINPUT77), .Z(new_n472));
  INV_X1    g286(.A(G469), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G140), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT78), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n281), .A2(G227), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g291(.A(KEYINPUT10), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n252), .A2(new_n254), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT83), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n214), .B2(new_n249), .ZN(new_n481));
  OAI211_X1 g295(.A(KEYINPUT83), .B(KEYINPUT1), .C1(new_n224), .C2(G146), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(G128), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n252), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n377), .A2(G104), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n350), .A2(G107), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT82), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n488), .B(G101), .C1(KEYINPUT82), .C2(new_n486), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT79), .B(G101), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT3), .B1(new_n350), .B2(G107), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT3), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n377), .A3(G104), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n490), .A2(new_n491), .A3(new_n493), .A4(new_n487), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n478), .B1(new_n485), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n478), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n256), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n493), .A3(new_n487), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n499), .A2(new_n500), .A3(G101), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n222), .A2(new_n226), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n499), .A2(G101), .ZN(new_n503));
  XOR2_X1   g317(.A(KEYINPUT79), .B(G101), .Z(new_n504));
  OAI21_X1  g318(.A(KEYINPUT4), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT80), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n499), .A2(G101), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT80), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n494), .A4(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT81), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n502), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n502), .B2(new_n510), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n496), .B(new_n498), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT84), .B1(new_n514), .B2(new_n247), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n491), .A2(new_n493), .A3(new_n487), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n500), .B1(new_n516), .B2(new_n490), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n508), .B1(new_n517), .B2(new_n507), .ZN(new_n518));
  INV_X1    g332(.A(new_n509), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n501), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n521), .A2(new_n270), .A3(new_n221), .A4(new_n217), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT81), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n502), .A2(new_n510), .A3(new_n511), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n496), .A2(new_n498), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT84), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n267), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n515), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n514), .A2(new_n247), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n477), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n495), .A2(new_n251), .A3(new_n255), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n485), .B2(new_n495), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n533), .A2(KEYINPUT12), .A3(new_n247), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT12), .B1(new_n533), .B2(new_n247), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n477), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n536), .B(new_n537), .C1(new_n515), .C2(new_n528), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n473), .B(new_n188), .C1(new_n531), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT86), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n482), .A2(G128), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n212), .A2(G143), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n215), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT83), .B1(new_n544), .B2(KEYINPUT1), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n484), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n495), .B1(new_n546), .B2(new_n255), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n498), .B1(new_n547), .B2(KEYINPUT10), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n523), .B2(new_n524), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n527), .B1(new_n549), .B2(new_n267), .ZN(new_n550));
  AND4_X1   g364(.A1(new_n527), .A2(new_n525), .A3(new_n526), .A4(new_n267), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n530), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n537), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n537), .B1(new_n515), .B2(new_n528), .ZN(new_n554));
  INV_X1    g368(.A(new_n536), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT86), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n557), .A2(new_n558), .A3(new_n473), .A4(new_n188), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n540), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n536), .B1(new_n515), .B2(new_n528), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(new_n477), .ZN(new_n562));
  INV_X1    g376(.A(new_n530), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n554), .B2(KEYINPUT85), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n477), .B1(new_n550), .B2(new_n551), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT85), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n562), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G469), .B1(new_n568), .B2(G902), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n472), .B1(new_n560), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G214), .B1(G237), .B2(G902), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n271), .A2(G125), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n251), .A2(new_n255), .A3(new_n327), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT87), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G224), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT7), .B1(new_n577), .B2(G953), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n578), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n572), .B(new_n573), .C1(new_n575), .C2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G110), .B(G122), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n501), .B1(new_n201), .B2(new_n204), .ZN(new_n584));
  INV_X1    g398(.A(new_n200), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(KEYINPUT5), .A3(new_n198), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT5), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n424), .A2(new_n587), .A3(G116), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n588), .A2(G113), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n495), .A2(new_n203), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n584), .A2(new_n510), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n589), .B1(new_n587), .B2(new_n202), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n203), .B1(new_n586), .B2(new_n589), .ZN(new_n595));
  INV_X1    g409(.A(new_n495), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n583), .B(KEYINPUT8), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n583), .A2(new_n592), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n582), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT6), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n592), .B2(new_n583), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n584), .A2(new_n510), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n590), .A2(new_n591), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n583), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n601), .A3(new_n606), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n577), .A2(G953), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n574), .B(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(G210), .B1(G237), .B2(G902), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n600), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n600), .B2(new_n612), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n571), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT88), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n600), .A2(new_n612), .ZN(new_n619));
  INV_X1    g433(.A(new_n613), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n600), .A2(new_n612), .A3(new_n613), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(KEYINPUT88), .A3(new_n571), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n470), .A2(new_n570), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(new_n504), .ZN(G3));
  INV_X1    g441(.A(new_n304), .ZN(new_n628));
  OAI21_X1  g442(.A(G472), .B1(new_n307), .B2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n468), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n570), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT92), .Z(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT95), .B(G478), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n402), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n402), .A2(KEYINPUT96), .A3(new_n634), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n398), .A2(new_n641), .A3(new_n401), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT93), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n398), .A2(KEYINPUT93), .A3(new_n401), .A4(new_n641), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n390), .A2(KEYINPUT94), .ZN(new_n646));
  OR3_X1    g460(.A1(new_n399), .A2(new_n400), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(new_n399), .B2(new_n400), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(KEYINPUT33), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n403), .A2(G902), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n644), .A2(new_n645), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n639), .A2(new_n640), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n640), .B1(new_n639), .B2(new_n651), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n370), .A2(new_n419), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n571), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n621), .B2(new_n622), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n412), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n633), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  INV_X1    g477(.A(KEYINPUT98), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n418), .B(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n405), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n367), .B(KEYINPUT20), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n659), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n633), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT99), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  AOI21_X1  g487(.A(G902), .B1(new_n553), .B2(new_n556), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n558), .B1(new_n674), .B2(new_n473), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n539), .A2(KEYINPUT86), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n569), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n448), .A2(new_n437), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT100), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n454), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n466), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n463), .A2(new_n465), .A3(new_n682), .ZN(new_n683));
  AND4_X1   g497(.A1(new_n420), .A2(new_n683), .A3(new_n628), .A4(new_n629), .ZN(new_n684));
  INV_X1    g498(.A(new_n472), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n677), .A2(new_n684), .A3(new_n685), .A4(new_n625), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  AND3_X1   g502(.A1(new_n321), .A2(new_n658), .A3(new_n683), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n406), .A2(new_n690), .A3(G902), .A4(G953), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT101), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n668), .B1(new_n408), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n689), .A2(new_n570), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  NAND2_X1  g509(.A1(new_n408), .A2(new_n692), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT39), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n570), .A2(KEYINPUT102), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT102), .B1(new_n570), .B2(new_n697), .ZN(new_n699));
  OR3_X1    g513(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT40), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT40), .B1(new_n698), .B2(new_n699), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n307), .A2(new_n306), .A3(new_n189), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n275), .A2(new_n279), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n285), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n278), .A2(new_n312), .ZN(new_n705));
  AOI21_X1  g519(.A(G902), .B1(new_n705), .B2(new_n302), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n187), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n683), .B1(new_n708), .B2(new_n308), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n623), .B(KEYINPUT38), .Z(new_n710));
  NOR2_X1   g524(.A1(new_n370), .A2(new_n419), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n710), .A2(new_n657), .A3(new_n711), .A4(new_n405), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n700), .A2(new_n701), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n220), .ZN(G45));
  NAND3_X1  g528(.A1(new_n654), .A2(new_n655), .A3(new_n696), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n689), .A2(new_n570), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  AOI21_X1  g532(.A(new_n473), .B1(new_n557), .B2(new_n188), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n560), .A2(new_n685), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n321), .A2(new_n469), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n719), .B1(new_n559), .B2(new_n540), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(KEYINPUT103), .A3(new_n685), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n723), .A2(new_n724), .A3(new_n660), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  AND3_X1   g543(.A1(new_n669), .A2(new_n321), .A3(new_n469), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n723), .A2(new_n726), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n723), .A2(new_n730), .A3(KEYINPUT104), .A4(new_n726), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  INV_X1    g550(.A(new_n721), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n321), .A2(new_n420), .A3(new_n683), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n658), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  OAI21_X1  g554(.A(KEYINPUT105), .B1(new_n711), .B2(new_n405), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  INV_X1    g556(.A(new_n405), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n742), .B(new_n743), .C1(new_n370), .C2(new_n419), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n741), .A2(new_n658), .A3(new_n412), .A4(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n285), .B1(new_n296), .B2(new_n313), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n288), .B2(new_n289), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n747), .A2(new_n189), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n469), .A2(new_n629), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n723), .A2(new_n726), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  NAND3_X1  g566(.A1(new_n683), .A2(new_n748), .A3(new_n629), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n715), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n685), .A3(new_n658), .A4(new_n725), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  AND4_X1   g570(.A1(KEYINPUT42), .A2(new_n654), .A3(new_n655), .A4(new_n696), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n623), .A2(new_n657), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n685), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n677), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT108), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n702), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n308), .B(new_n320), .C1(new_n702), .C2(new_n762), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n469), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT109), .B1(new_n761), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n320), .A2(new_n308), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n762), .B1(new_n304), .B2(KEYINPUT32), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n468), .B1(new_n770), .B2(new_n763), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n759), .B1(new_n560), .B2(new_n569), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n757), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n724), .A3(new_n716), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n776), .A2(KEYINPUT107), .A3(new_n777), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n775), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n245), .ZN(G33));
  NAND3_X1  g597(.A1(new_n773), .A2(new_n724), .A3(new_n693), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n654), .B2(new_n711), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n654), .A2(new_n787), .A3(new_n711), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n683), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n630), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n786), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n758), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n791), .A2(new_n786), .A3(new_n792), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(G469), .B1(new_n568), .B2(KEYINPUT45), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(KEYINPUT45), .B2(new_n568), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT46), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n473), .A2(new_n188), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n798), .B2(new_n800), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n560), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n796), .A2(new_n803), .A3(new_n685), .A4(new_n697), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n685), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n803), .A2(KEYINPUT47), .A3(new_n685), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n758), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n321), .A2(new_n715), .A3(new_n811), .A4(new_n469), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n324), .ZN(G42));
  INV_X1    g628(.A(new_n790), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n815), .A2(new_n408), .A3(new_n788), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n749), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n616), .A3(new_n721), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(KEYINPUT116), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n560), .A2(new_n720), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n408), .A3(new_n759), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n822), .A2(new_n789), .A3(new_n790), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT48), .B1(new_n823), .B2(new_n771), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(G952), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n826), .B(G953), .C1(new_n819), .C2(KEYINPUT116), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(KEYINPUT48), .A3(new_n771), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n708), .A2(new_n308), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n822), .A2(new_n469), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n655), .A3(new_n654), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n825), .A2(new_n827), .A3(new_n828), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n818), .A2(new_n811), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n821), .A2(new_n685), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n810), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n654), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n832), .A2(new_n711), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n817), .A2(new_n657), .A3(new_n710), .A4(new_n737), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n753), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n823), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n837), .A2(new_n839), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n834), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n842), .A2(new_n839), .A3(new_n844), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(new_n837), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n850), .B2(KEYINPUT51), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n845), .A2(KEYINPUT115), .A3(new_n846), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n727), .A2(new_n739), .A3(new_n751), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n735), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n782), .ZN(new_n856));
  INV_X1    g670(.A(new_n412), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n370), .A2(new_n419), .A3(new_n857), .A4(new_n405), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n858), .A2(new_n618), .A3(new_n624), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n677), .A2(new_n685), .A3(new_n631), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n686), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT110), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n686), .A2(new_n860), .A3(KEYINPUT110), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n656), .A2(new_n630), .A3(new_n857), .A4(new_n468), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n570), .B(new_n625), .C1(new_n865), .C2(new_n470), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n863), .A2(new_n866), .A3(KEYINPUT111), .A4(new_n864), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n667), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n405), .A2(new_n696), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n811), .A2(new_n872), .A3(new_n665), .A4(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n570), .A2(new_n874), .A3(new_n321), .A4(new_n683), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n773), .A2(new_n754), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n784), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n694), .A2(new_n755), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n741), .A2(new_n658), .A3(new_n744), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n570), .A2(new_n696), .A3(new_n709), .A4(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(KEYINPUT52), .A3(new_n717), .A4(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n694), .A2(new_n881), .A3(new_n717), .A4(new_n755), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n877), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n856), .A2(new_n871), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT53), .B1(new_n878), .B2(KEYINPUT52), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT53), .B1(new_n879), .B2(new_n884), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n869), .B2(new_n870), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT112), .B1(new_n855), .B2(new_n782), .ZN(new_n896));
  INV_X1    g710(.A(new_n781), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT107), .B1(new_n776), .B2(new_n777), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n767), .B(new_n774), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT112), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n735), .A4(new_n854), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n895), .A2(new_n896), .A3(new_n901), .A4(new_n886), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n889), .A2(new_n893), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n892), .A2(KEYINPUT113), .A3(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n903), .A2(KEYINPUT113), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n853), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(G952), .A2(G953), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT117), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n821), .A2(KEYINPUT49), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n821), .A2(KEYINPUT49), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n654), .A2(new_n685), .A3(new_n571), .A4(new_n711), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n468), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n829), .A3(new_n710), .A4(new_n912), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n906), .A2(new_n908), .B1(new_n909), .B2(new_n913), .ZN(G75));
  NAND2_X1  g728(.A1(new_n826), .A2(G953), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT118), .Z(new_n916));
  NAND2_X1  g730(.A1(new_n608), .A2(new_n609), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n611), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT55), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n188), .B1(new_n889), .B2(new_n902), .ZN(new_n920));
  AOI211_X1 g734(.A(KEYINPUT56), .B(new_n919), .C1(new_n920), .C2(G210), .ZN(new_n921));
  INV_X1    g735(.A(new_n919), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n889), .A2(new_n902), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(G210), .A3(G902), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT56), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n916), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(KEYINPUT119), .B(new_n916), .C1(new_n921), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(G51));
  XNOR2_X1  g745(.A(new_n798), .B(KEYINPUT121), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n920), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n800), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n889), .A2(new_n893), .A3(new_n902), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n893), .B1(new_n889), .B2(new_n902), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n933), .B1(new_n938), .B2(new_n557), .ZN(new_n939));
  INV_X1    g753(.A(new_n916), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT122), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  INV_X1    g756(.A(new_n557), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n923), .A2(KEYINPUT54), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n903), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n935), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n942), .B(new_n916), .C1(new_n946), .C2(new_n933), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n941), .A2(new_n947), .ZN(G54));
  AND3_X1   g762(.A1(new_n920), .A2(KEYINPUT58), .A3(G475), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n362), .A2(new_n366), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n916), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n950), .B2(new_n949), .ZN(G60));
  INV_X1    g766(.A(new_n945), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT59), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n644), .A2(new_n645), .A3(new_n649), .A4(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n916), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n904), .A2(new_n905), .A3(new_n955), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n644), .A2(new_n645), .A3(new_n649), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(G63));
  NAND2_X1  g774(.A1(G217), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT60), .Z(new_n962));
  AOI21_X1  g776(.A(new_n458), .B1(new_n923), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(new_n940), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT61), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n923), .A2(new_n681), .A3(new_n962), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n964), .B(new_n967), .C1(new_n965), .C2(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(G66));
  AOI21_X1  g785(.A(new_n281), .B1(new_n410), .B2(G224), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n871), .A2(new_n735), .A3(new_n854), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(KEYINPUT124), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(KEYINPUT124), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n972), .B1(new_n976), .B2(new_n281), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n917), .B1(G898), .B2(new_n281), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n977), .B(new_n978), .Z(G69));
  OAI21_X1  g793(.A(new_n260), .B1(new_n274), .B2(KEYINPUT30), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT125), .Z(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(new_n331), .ZN(new_n982));
  INV_X1    g796(.A(new_n806), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n771), .A2(new_n880), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n983), .B(new_n697), .C1(new_n796), .C2(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n879), .A2(new_n717), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n899), .A3(new_n784), .A4(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n281), .B1(new_n987), .B2(new_n813), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n690), .A2(G953), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n698), .A2(new_n699), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n711), .A2(new_n743), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n811), .B1(new_n656), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(new_n724), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n804), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n810), .B2(new_n812), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n713), .A2(new_n986), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(KEYINPUT62), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n281), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n990), .B1(new_n1001), .B2(new_n982), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n281), .B1(G227), .B2(G900), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1002), .B(new_n1003), .Z(G72));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n976), .B2(new_n1000), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n285), .A3(new_n703), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n704), .A2(new_n310), .A3(new_n1006), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n891), .A2(KEYINPUT127), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT127), .B1(new_n891), .B2(new_n1009), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1008), .B(new_n916), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n987), .A2(new_n813), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1013), .A2(new_n974), .A3(new_n975), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n1014), .A2(KEYINPUT126), .A3(new_n1006), .ZN(new_n1015));
  AOI21_X1  g829(.A(KEYINPUT126), .B1(new_n1014), .B2(new_n1006), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1015), .A2(new_n1016), .A3(new_n310), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1012), .A2(new_n1017), .ZN(G57));
endmodule


