

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(n395), .B(n394), .ZN(n542) );
  NOR2_X1 U325 ( .A1(n422), .A2(n529), .ZN(n572) );
  INV_X1 U326 ( .A(n542), .ZN(n544) );
  XNOR2_X1 U327 ( .A(n345), .B(n344), .ZN(n579) );
  XNOR2_X1 U328 ( .A(n579), .B(KEYINPUT41), .ZN(n551) );
  XOR2_X1 U329 ( .A(n484), .B(KEYINPUT28), .Z(n548) );
  XNOR2_X1 U330 ( .A(n461), .B(KEYINPUT58), .ZN(n462) );
  XNOR2_X1 U331 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(G50GAT), .B(G162GAT), .Z(n435) );
  XOR2_X1 U333 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n293) );
  XNOR2_X1 U334 ( .A(G134GAT), .B(KEYINPUT73), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U336 ( .A(n435), .B(n294), .Z(n296) );
  NAND2_X1 U337 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n313) );
  XOR2_X1 U339 ( .A(KEYINPUT72), .B(KEYINPUT74), .Z(n298) );
  XNOR2_X1 U340 ( .A(KEYINPUT75), .B(KEYINPUT11), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n300) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n299), .B(G218GAT), .ZN(n316) );
  XOR2_X1 U344 ( .A(n300), .B(n316), .Z(n311) );
  INV_X1 U345 ( .A(KEYINPUT67), .ZN(n301) );
  NAND2_X1 U346 ( .A1(KEYINPUT7), .A2(n301), .ZN(n304) );
  INV_X1 U347 ( .A(KEYINPUT7), .ZN(n302) );
  NAND2_X1 U348 ( .A1(n302), .A2(KEYINPUT67), .ZN(n303) );
  NAND2_X1 U349 ( .A1(n304), .A2(n303), .ZN(n306) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G29GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U352 ( .A(KEYINPUT8), .B(n307), .Z(n349) );
  XOR2_X1 U353 ( .A(G85GAT), .B(G92GAT), .Z(n309) );
  XNOR2_X1 U354 ( .A(G99GAT), .B(G106GAT), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n336) );
  XNOR2_X1 U356 ( .A(n349), .B(n336), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n570) );
  INV_X1 U359 ( .A(n570), .ZN(n384) );
  XOR2_X1 U360 ( .A(KEYINPUT76), .B(n384), .Z(n490) );
  XOR2_X1 U361 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n397) );
  XOR2_X1 U362 ( .A(G92GAT), .B(KEYINPUT99), .Z(n315) );
  NAND2_X1 U363 ( .A1(G226GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n317) );
  XOR2_X1 U365 ( .A(n317), .B(n316), .Z(n321) );
  XOR2_X1 U366 ( .A(G211GAT), .B(KEYINPUT90), .Z(n319) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n428) );
  XNOR2_X1 U369 ( .A(n428), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U371 ( .A(G176GAT), .B(G64GAT), .Z(n343) );
  XOR2_X1 U372 ( .A(n322), .B(n343), .Z(n327) );
  XOR2_X1 U373 ( .A(G169GAT), .B(G8GAT), .Z(n352) );
  XOR2_X1 U374 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n324) );
  XNOR2_X1 U375 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U377 ( .A(KEYINPUT89), .B(n325), .Z(n457) );
  XNOR2_X1 U378 ( .A(n352), .B(n457), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n533) );
  XNOR2_X1 U380 ( .A(G78GAT), .B(G204GAT), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n328), .B(G148GAT), .ZN(n433) );
  XOR2_X1 U382 ( .A(G120GAT), .B(G71GAT), .Z(n448) );
  XNOR2_X1 U383 ( .A(n433), .B(n448), .ZN(n329) );
  AND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  NAND2_X1 U385 ( .A1(n329), .A2(n330), .ZN(n334) );
  INV_X1 U386 ( .A(n329), .ZN(n332) );
  INV_X1 U387 ( .A(n330), .ZN(n331) );
  NAND2_X1 U388 ( .A1(n332), .A2(n331), .ZN(n333) );
  NAND2_X1 U389 ( .A1(n334), .A2(n333), .ZN(n335) );
  XOR2_X1 U390 ( .A(n335), .B(KEYINPUT32), .Z(n338) );
  XNOR2_X1 U391 ( .A(n336), .B(KEYINPUT31), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U393 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n340) );
  XNOR2_X1 U394 ( .A(KEYINPUT33), .B(KEYINPUT68), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U396 ( .A(n342), .B(n341), .Z(n345) );
  XOR2_X1 U397 ( .A(KEYINPUT13), .B(G57GAT), .Z(n374) );
  XNOR2_X1 U398 ( .A(n343), .B(n374), .ZN(n344) );
  XOR2_X1 U399 ( .A(G15GAT), .B(G22GAT), .Z(n347) );
  XNOR2_X1 U400 ( .A(G141GAT), .B(G197GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n360) );
  XOR2_X1 U403 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n351) );
  XNOR2_X1 U404 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n356) );
  XOR2_X1 U406 ( .A(G36GAT), .B(G50GAT), .Z(n354) );
  XOR2_X1 U407 ( .A(G113GAT), .B(G1GAT), .Z(n411) );
  XNOR2_X1 U408 ( .A(n352), .B(n411), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U410 ( .A(n356), .B(n355), .Z(n358) );
  NAND2_X1 U411 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U413 ( .A(n360), .B(n359), .Z(n549) );
  NAND2_X1 U414 ( .A1(n551), .A2(n549), .ZN(n362) );
  XNOR2_X1 U415 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n386) );
  XOR2_X1 U417 ( .A(G64GAT), .B(G71GAT), .Z(n364) );
  XNOR2_X1 U418 ( .A(G8GAT), .B(G183GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U420 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n366) );
  XNOR2_X1 U421 ( .A(G1GAT), .B(KEYINPUT82), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U423 ( .A(n368), .B(n367), .Z(n373) );
  XOR2_X1 U424 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n370) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U427 ( .A(KEYINPUT78), .B(n371), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U429 ( .A(n374), .B(G78GAT), .Z(n376) );
  XOR2_X1 U430 ( .A(G22GAT), .B(G155GAT), .Z(n434) );
  XNOR2_X1 U431 ( .A(G211GAT), .B(n434), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U433 ( .A(n378), .B(n377), .Z(n383) );
  XOR2_X1 U434 ( .A(G15GAT), .B(G127GAT), .Z(n445) );
  XOR2_X1 U435 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n380) );
  XNOR2_X1 U436 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n445), .B(n381), .ZN(n382) );
  XOR2_X1 U439 ( .A(n383), .B(n382), .Z(n554) );
  NOR2_X1 U440 ( .A1(n384), .A2(n554), .ZN(n385) );
  AND2_X1 U441 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n387), .B(KEYINPUT47), .ZN(n393) );
  INV_X1 U443 ( .A(n554), .ZN(n584) );
  INV_X1 U444 ( .A(n490), .ZN(n557) );
  XOR2_X1 U445 ( .A(KEYINPUT36), .B(n557), .Z(n588) );
  NOR2_X1 U446 ( .A1(n584), .A2(n588), .ZN(n389) );
  XNOR2_X1 U447 ( .A(KEYINPUT45), .B(KEYINPUT115), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n391) );
  INV_X1 U449 ( .A(n549), .ZN(n574) );
  NAND2_X1 U450 ( .A1(n574), .A2(n579), .ZN(n390) );
  OR2_X1 U451 ( .A1(n391), .A2(n390), .ZN(n392) );
  NAND2_X1 U452 ( .A1(n393), .A2(n392), .ZN(n395) );
  XNOR2_X1 U453 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n394) );
  NAND2_X1 U454 ( .A1(n533), .A2(n542), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n422) );
  XOR2_X1 U456 ( .A(G57GAT), .B(G148GAT), .Z(n399) );
  XNOR2_X1 U457 ( .A(G120GAT), .B(G127GAT), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U459 ( .A(G85GAT), .B(G155GAT), .Z(n401) );
  XNOR2_X1 U460 ( .A(G29GAT), .B(G162GAT), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n421) );
  XOR2_X1 U463 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n405) );
  XNOR2_X1 U464 ( .A(KEYINPUT93), .B(KEYINPUT97), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U466 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n407) );
  XNOR2_X1 U467 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n419) );
  XNOR2_X1 U470 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n410), .B(KEYINPUT86), .ZN(n449) );
  XOR2_X1 U472 ( .A(n449), .B(n411), .Z(n413) );
  NAND2_X1 U473 ( .A1(G225GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U475 ( .A(n414), .B(KEYINPUT98), .Z(n417) );
  XNOR2_X1 U476 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n415) );
  XNOR2_X1 U477 ( .A(n415), .B(KEYINPUT2), .ZN(n429) );
  XNOR2_X1 U478 ( .A(n429), .B(KEYINPUT1), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n529) );
  XOR2_X1 U482 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n424) );
  XNOR2_X1 U483 ( .A(G218GAT), .B(G106GAT), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n439) );
  XOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n426) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U488 ( .A(n427), .B(KEYINPUT24), .Z(n431) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U491 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n484) );
  NAND2_X1 U495 ( .A1(n572), .A2(n484), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n440), .B(KEYINPUT120), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n441), .B(KEYINPUT55), .ZN(n460) );
  XOR2_X1 U498 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n443) );
  XNOR2_X1 U499 ( .A(G190GAT), .B(KEYINPUT88), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U501 ( .A(n444), .B(G99GAT), .Z(n447) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n453) );
  XOR2_X1 U504 ( .A(n449), .B(n448), .Z(n451) );
  NAND2_X1 U505 ( .A1(G227GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U507 ( .A(n453), .B(n452), .Z(n459) );
  XOR2_X1 U508 ( .A(G176GAT), .B(KEYINPUT64), .Z(n455) );
  XNOR2_X1 U509 ( .A(G169GAT), .B(G113GAT), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U511 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(n545) );
  NAND2_X1 U513 ( .A1(n460), .A2(n545), .ZN(n469) );
  NOR2_X1 U514 ( .A1(n490), .A2(n469), .ZN(n463) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n574), .A2(n469), .ZN(n465) );
  XNOR2_X1 U517 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n465), .B(n464), .ZN(G1348GAT) );
  INV_X1 U519 ( .A(n551), .ZN(n565) );
  NOR2_X1 U520 ( .A1(n565), .A2(n469), .ZN(n468) );
  XNOR2_X1 U521 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n466) );
  XNOR2_X1 U522 ( .A(n466), .B(G176GAT), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n468), .B(n467), .ZN(G1349GAT) );
  NOR2_X1 U524 ( .A1(n584), .A2(n469), .ZN(n472) );
  XNOR2_X1 U525 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(G183GAT), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n472), .B(n471), .ZN(G1350GAT) );
  XOR2_X1 U528 ( .A(KEYINPUT104), .B(KEYINPUT34), .Z(n496) );
  NAND2_X1 U529 ( .A1(n549), .A2(n579), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT71), .ZN(n507) );
  NAND2_X1 U531 ( .A1(n545), .A2(n533), .ZN(n474) );
  XOR2_X1 U532 ( .A(KEYINPUT101), .B(n474), .Z(n475) );
  NAND2_X1 U533 ( .A1(n475), .A2(n484), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(KEYINPUT25), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(KEYINPUT102), .ZN(n480) );
  NOR2_X1 U536 ( .A1(n545), .A2(n484), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT26), .B(n478), .ZN(n573) );
  XNOR2_X1 U538 ( .A(n533), .B(KEYINPUT27), .ZN(n483) );
  AND2_X1 U539 ( .A1(n573), .A2(n483), .ZN(n479) );
  NOR2_X1 U540 ( .A1(n480), .A2(n479), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT103), .B(n481), .Z(n482) );
  NOR2_X1 U542 ( .A1(n529), .A2(n482), .ZN(n489) );
  NAND2_X1 U543 ( .A1(n529), .A2(n483), .ZN(n543) );
  NOR2_X1 U544 ( .A1(n545), .A2(n543), .ZN(n486) );
  INV_X1 U545 ( .A(n548), .ZN(n485) );
  NAND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT100), .B(n487), .Z(n488) );
  NOR2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n504) );
  XOR2_X1 U549 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n492) );
  NAND2_X1 U550 ( .A1(n490), .A2(n554), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(KEYINPUT16), .ZN(n494) );
  NOR2_X1 U553 ( .A1(n504), .A2(n494), .ZN(n518) );
  AND2_X1 U554 ( .A1(n507), .A2(n518), .ZN(n502) );
  NAND2_X1 U555 ( .A1(n502), .A2(n529), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U557 ( .A(G1GAT), .B(n497), .Z(G1324GAT) );
  NAND2_X1 U558 ( .A1(n502), .A2(n533), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n498), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n500) );
  NAND2_X1 U561 ( .A1(n502), .A2(n545), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U563 ( .A(G15GAT), .B(n501), .Z(G1326GAT) );
  NAND2_X1 U564 ( .A1(n502), .A2(n548), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n510) );
  NOR2_X1 U567 ( .A1(n588), .A2(n504), .ZN(n505) );
  NAND2_X1 U568 ( .A1(n584), .A2(n505), .ZN(n506) );
  XNOR2_X1 U569 ( .A(KEYINPUT37), .B(n506), .ZN(n528) );
  NAND2_X1 U570 ( .A1(n528), .A2(n507), .ZN(n508) );
  XOR2_X1 U571 ( .A(KEYINPUT38), .B(n508), .Z(n515) );
  NAND2_X1 U572 ( .A1(n529), .A2(n515), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G29GAT), .B(n511), .ZN(G1328GAT) );
  NAND2_X1 U575 ( .A1(n515), .A2(n533), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U577 ( .A1(n515), .A2(n545), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT40), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G43GAT), .B(n514), .ZN(G1330GAT) );
  XOR2_X1 U580 ( .A(G50GAT), .B(KEYINPUT107), .Z(n517) );
  NAND2_X1 U581 ( .A1(n548), .A2(n515), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1331GAT) );
  NOR2_X1 U583 ( .A1(n565), .A2(n549), .ZN(n527) );
  AND2_X1 U584 ( .A1(n527), .A2(n518), .ZN(n524) );
  NAND2_X1 U585 ( .A1(n524), .A2(n529), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n519), .B(KEYINPUT42), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1332GAT) );
  NAND2_X1 U589 ( .A1(n524), .A2(n533), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U591 ( .A1(n524), .A2(n545), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n523), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U593 ( .A(G78GAT), .B(KEYINPUT43), .Z(n526) );
  NAND2_X1 U594 ( .A1(n524), .A2(n548), .ZN(n525) );
  XNOR2_X1 U595 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n531) );
  AND2_X1 U597 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n537), .A2(n529), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U600 ( .A(G85GAT), .B(n532), .ZN(G1336GAT) );
  XOR2_X1 U601 ( .A(G92GAT), .B(KEYINPUT111), .Z(n535) );
  NAND2_X1 U602 ( .A1(n537), .A2(n533), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(G1337GAT) );
  NAND2_X1 U604 ( .A1(n537), .A2(n545), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U606 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n539) );
  NAND2_X1 U608 ( .A1(n537), .A2(n548), .ZN(n538) );
  XNOR2_X1 U609 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(G1339GAT) );
  NOR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n561) );
  NAND2_X1 U612 ( .A1(n545), .A2(n561), .ZN(n546) );
  XOR2_X1 U613 ( .A(KEYINPUT117), .B(n546), .Z(n547) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n549), .A2(n558), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U617 ( .A(G120GAT), .B(KEYINPUT49), .Z(n553) );
  NAND2_X1 U618 ( .A1(n558), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1341GAT) );
  NAND2_X1 U620 ( .A1(n554), .A2(n558), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT50), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G127GAT), .B(n556), .ZN(G1342GAT) );
  XOR2_X1 U623 ( .A(G134GAT), .B(KEYINPUT51), .Z(n560) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1343GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n573), .ZN(n569) );
  NOR2_X1 U627 ( .A1(n574), .A2(n569), .ZN(n562) );
  XOR2_X1 U628 ( .A(G141GAT), .B(n562), .Z(G1344GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n564) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n567) );
  NOR2_X1 U632 ( .A1(n565), .A2(n569), .ZN(n566) );
  XOR2_X1 U633 ( .A(n567), .B(n566), .Z(G1345GAT) );
  NOR2_X1 U634 ( .A1(n584), .A2(n569), .ZN(n568) );
  XOR2_X1 U635 ( .A(G155GAT), .B(n568), .Z(G1346GAT) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(G162GAT), .B(n571), .Z(G1347GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n573), .ZN(n587) );
  NOR2_X1 U639 ( .A1(n574), .A2(n587), .ZN(n578) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT124), .ZN(n576) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n587), .A2(n579), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n587), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

