

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U546 ( .A1(n517), .A2(G2104), .ZN(n852) );
  NOR2_X1 U547 ( .A1(n670), .A2(n717), .ZN(n510) );
  NAND2_X1 U548 ( .A1(n652), .A2(G1341), .ZN(n511) );
  INV_X1 U549 ( .A(n652), .ZN(n632) );
  XNOR2_X1 U550 ( .A(n640), .B(KEYINPUT101), .ZN(n641) );
  XNOR2_X1 U551 ( .A(n642), .B(n641), .ZN(n643) );
  INV_X1 U552 ( .A(KEYINPUT102), .ZN(n650) );
  NAND2_X1 U553 ( .A1(n678), .A2(n590), .ZN(n652) );
  NOR2_X1 U554 ( .A1(G651), .A2(n570), .ZN(n774) );
  AND2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n856) );
  NAND2_X1 U556 ( .A1(n856), .A2(G113), .ZN(n514) );
  INV_X1 U557 ( .A(G2105), .ZN(n517) );
  NAND2_X1 U558 ( .A1(G101), .A2(n852), .ZN(n512) );
  XOR2_X1 U559 ( .A(KEYINPUT23), .B(n512), .Z(n513) );
  NAND2_X1 U560 ( .A1(n514), .A2(n513), .ZN(n521) );
  XNOR2_X1 U561 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n516) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  XNOR2_X2 U563 ( .A(n516), .B(n515), .ZN(n853) );
  NAND2_X1 U564 ( .A1(G137), .A2(n853), .ZN(n519) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n517), .ZN(n858) );
  NAND2_X1 U566 ( .A1(G125), .A2(n858), .ZN(n518) );
  NAND2_X1 U567 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U568 ( .A1(n521), .A2(n520), .ZN(G160) );
  NAND2_X1 U569 ( .A1(G102), .A2(n852), .ZN(n523) );
  NAND2_X1 U570 ( .A1(G138), .A2(n853), .ZN(n522) );
  NAND2_X1 U571 ( .A1(n523), .A2(n522), .ZN(n527) );
  NAND2_X1 U572 ( .A1(G114), .A2(n856), .ZN(n525) );
  NAND2_X1 U573 ( .A1(G126), .A2(n858), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U575 ( .A1(n527), .A2(n526), .ZN(G164) );
  NOR2_X1 U576 ( .A1(G543), .A2(G651), .ZN(n528) );
  XNOR2_X1 U577 ( .A(n528), .B(KEYINPUT64), .ZN(n767) );
  NAND2_X1 U578 ( .A1(G91), .A2(n767), .ZN(n529) );
  XOR2_X1 U579 ( .A(KEYINPUT69), .B(n529), .Z(n531) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n570) );
  INV_X1 U581 ( .A(G651), .ZN(n533) );
  NOR2_X1 U582 ( .A1(n570), .A2(n533), .ZN(n770) );
  NAND2_X1 U583 ( .A1(n770), .A2(G78), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U585 ( .A(KEYINPUT70), .B(n532), .Z(n538) );
  NOR2_X1 U586 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n534), .Z(n766) );
  NAND2_X1 U588 ( .A1(G65), .A2(n766), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G53), .A2(n774), .ZN(n535) );
  AND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n538), .A2(n537), .ZN(G299) );
  NAND2_X1 U592 ( .A1(G64), .A2(n766), .ZN(n540) );
  NAND2_X1 U593 ( .A1(G52), .A2(n774), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U595 ( .A(KEYINPUT68), .B(n541), .ZN(n546) );
  NAND2_X1 U596 ( .A1(n770), .A2(G77), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G90), .A2(n767), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U599 ( .A(KEYINPUT9), .B(n544), .Z(n545) );
  NOR2_X1 U600 ( .A1(n546), .A2(n545), .ZN(G171) );
  INV_X1 U601 ( .A(G171), .ZN(G301) );
  NAND2_X1 U602 ( .A1(n774), .A2(G51), .ZN(n547) );
  XOR2_X1 U603 ( .A(KEYINPUT77), .B(n547), .Z(n549) );
  NAND2_X1 U604 ( .A1(n766), .A2(G63), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U606 ( .A(KEYINPUT6), .B(n550), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G89), .A2(n767), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G76), .A2(n770), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U611 ( .A(KEYINPUT5), .B(n554), .Z(n555) );
  NOR2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n559) );
  XNOR2_X1 U613 ( .A(KEYINPUT79), .B(KEYINPUT7), .ZN(n557) );
  XNOR2_X1 U614 ( .A(n557), .B(KEYINPUT78), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n559), .B(n558), .ZN(G168) );
  XOR2_X1 U616 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U617 ( .A1(n770), .A2(G75), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G88), .A2(n767), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G62), .A2(n766), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G50), .A2(n774), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U623 ( .A1(n565), .A2(n564), .ZN(G166) );
  XNOR2_X1 U624 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  NAND2_X1 U625 ( .A1(G49), .A2(n774), .ZN(n567) );
  NAND2_X1 U626 ( .A1(G74), .A2(G651), .ZN(n566) );
  NAND2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U628 ( .A(KEYINPUT86), .B(n568), .ZN(n569) );
  NOR2_X1 U629 ( .A1(n766), .A2(n569), .ZN(n572) );
  NAND2_X1 U630 ( .A1(n570), .A2(G87), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U632 ( .A1(n766), .A2(G61), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G86), .A2(n767), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U635 ( .A1(G73), .A2(n770), .ZN(n575) );
  XNOR2_X1 U636 ( .A(n575), .B(KEYINPUT2), .ZN(n576) );
  XNOR2_X1 U637 ( .A(n576), .B(KEYINPUT87), .ZN(n577) );
  NOR2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U639 ( .A(n579), .B(KEYINPUT88), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G48), .A2(n774), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n581), .A2(n580), .ZN(G305) );
  NAND2_X1 U642 ( .A1(n770), .A2(G72), .ZN(n583) );
  NAND2_X1 U643 ( .A1(G85), .A2(n767), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U645 ( .A(KEYINPUT66), .B(n584), .ZN(n587) );
  NAND2_X1 U646 ( .A1(G60), .A2(n766), .ZN(n585) );
  XNOR2_X1 U647 ( .A(KEYINPUT67), .B(n585), .ZN(n586) );
  NOR2_X1 U648 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n774), .A2(G47), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n589), .A2(n588), .ZN(G290) );
  NOR2_X1 U651 ( .A1(G164), .A2(G1384), .ZN(n678) );
  NAND2_X1 U652 ( .A1(G160), .A2(G40), .ZN(n677) );
  XOR2_X1 U653 ( .A(KEYINPUT96), .B(n677), .Z(n590) );
  NAND2_X1 U654 ( .A1(n632), .A2(G2072), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT27), .ZN(n593) );
  INV_X1 U656 ( .A(G1956), .ZN(n982) );
  NOR2_X1 U657 ( .A1(n982), .A2(n632), .ZN(n592) );
  NOR2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n595) );
  INV_X1 U659 ( .A(G299), .ZN(n596) );
  NOR2_X1 U660 ( .A1(n595), .A2(n596), .ZN(n594) );
  XOR2_X1 U661 ( .A(n594), .B(KEYINPUT28), .Z(n630) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(n628) );
  XOR2_X1 U663 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n598) );
  NAND2_X1 U664 ( .A1(G56), .A2(n766), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n598), .B(n597), .ZN(n604) );
  NAND2_X1 U666 ( .A1(G81), .A2(n767), .ZN(n599) );
  XNOR2_X1 U667 ( .A(n599), .B(KEYINPUT12), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G68), .A2(n770), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U670 ( .A(KEYINPUT13), .B(n602), .Z(n603) );
  NOR2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U672 ( .A1(n774), .A2(G43), .ZN(n605) );
  NAND2_X1 U673 ( .A1(n606), .A2(n605), .ZN(n952) );
  XOR2_X1 U674 ( .A(G1996), .B(KEYINPUT99), .Z(n906) );
  NAND2_X1 U675 ( .A1(n632), .A2(n906), .ZN(n607) );
  XNOR2_X1 U676 ( .A(KEYINPUT26), .B(n607), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n608), .A2(n511), .ZN(n609) );
  NOR2_X1 U678 ( .A1(n952), .A2(n609), .ZN(n623) );
  NAND2_X1 U679 ( .A1(G92), .A2(n767), .ZN(n610) );
  XNOR2_X1 U680 ( .A(n610), .B(KEYINPUT74), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G66), .A2(n766), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT75), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G54), .A2(n774), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n770), .A2(G79), .ZN(n616) );
  XOR2_X1 U687 ( .A(KEYINPUT76), .B(n616), .Z(n617) );
  NOR2_X1 U688 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U689 ( .A(KEYINPUT15), .B(n619), .ZN(n968) );
  NAND2_X1 U690 ( .A1(G1348), .A2(n652), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n632), .A2(G2067), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n624) );
  NOR2_X1 U693 ( .A1(n968), .A2(n624), .ZN(n622) );
  OR2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n968), .A2(n624), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n631), .B(KEYINPUT29), .ZN(n638) );
  NOR2_X1 U700 ( .A1(n632), .A2(G1961), .ZN(n633) );
  XOR2_X1 U701 ( .A(KEYINPUT97), .B(n633), .Z(n635) );
  XOR2_X1 U702 ( .A(G2078), .B(KEYINPUT25), .Z(n907) );
  NOR2_X1 U703 ( .A1(n907), .A2(n652), .ZN(n634) );
  NOR2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n644) );
  NOR2_X1 U705 ( .A1(n644), .A2(G301), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n636), .B(KEYINPUT98), .ZN(n637) );
  NOR2_X1 U707 ( .A1(n638), .A2(n637), .ZN(n649) );
  NAND2_X1 U708 ( .A1(G8), .A2(n652), .ZN(n717) );
  NOR2_X1 U709 ( .A1(G1966), .A2(n717), .ZN(n663) );
  NOR2_X1 U710 ( .A1(G2084), .A2(n652), .ZN(n664) );
  NOR2_X1 U711 ( .A1(n663), .A2(n664), .ZN(n639) );
  NAND2_X1 U712 ( .A1(G8), .A2(n639), .ZN(n642) );
  XOR2_X1 U713 ( .A(KEYINPUT30), .B(KEYINPUT100), .Z(n640) );
  NOR2_X1 U714 ( .A1(G168), .A2(n643), .ZN(n646) );
  AND2_X1 U715 ( .A1(G301), .A2(n644), .ZN(n645) );
  NOR2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U717 ( .A(n647), .B(KEYINPUT31), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n651) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(n661) );
  NAND2_X1 U720 ( .A1(n661), .A2(G286), .ZN(n657) );
  NOR2_X1 U721 ( .A1(G1971), .A2(n717), .ZN(n654) );
  NOR2_X1 U722 ( .A1(G2090), .A2(n652), .ZN(n653) );
  NOR2_X1 U723 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n655), .A2(G303), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U726 ( .A(KEYINPUT103), .B(n658), .Z(n659) );
  NAND2_X1 U727 ( .A1(G8), .A2(n659), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(KEYINPUT32), .ZN(n668) );
  INV_X1 U729 ( .A(n661), .ZN(n662) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U731 ( .A1(G8), .A2(n664), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n712) );
  NOR2_X1 U734 ( .A1(G1976), .A2(G288), .ZN(n673) );
  NOR2_X1 U735 ( .A1(G1971), .A2(G303), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n673), .A2(n669), .ZN(n960) );
  NAND2_X1 U737 ( .A1(n712), .A2(n960), .ZN(n671) );
  NAND2_X1 U738 ( .A1(G1976), .A2(G288), .ZN(n956) );
  INV_X1 U739 ( .A(n956), .ZN(n670) );
  AND2_X1 U740 ( .A1(n671), .A2(n510), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n672), .A2(KEYINPUT33), .ZN(n676) );
  NAND2_X1 U742 ( .A1(n673), .A2(KEYINPUT33), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n674), .A2(n717), .ZN(n675) );
  NOR2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n709) );
  XOR2_X1 U745 ( .A(G1981), .B(G305), .Z(n949) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n736) );
  XNOR2_X1 U747 ( .A(KEYINPUT37), .B(G2067), .ZN(n733) );
  NAND2_X1 U748 ( .A1(G116), .A2(n856), .ZN(n680) );
  NAND2_X1 U749 ( .A1(G128), .A2(n858), .ZN(n679) );
  NAND2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U751 ( .A(n681), .B(KEYINPUT35), .ZN(n686) );
  NAND2_X1 U752 ( .A1(G104), .A2(n852), .ZN(n683) );
  NAND2_X1 U753 ( .A1(G140), .A2(n853), .ZN(n682) );
  NAND2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U755 ( .A(KEYINPUT34), .B(n684), .Z(n685) );
  NAND2_X1 U756 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U757 ( .A(n687), .B(KEYINPUT36), .Z(n869) );
  NOR2_X1 U758 ( .A1(n733), .A2(n869), .ZN(n935) );
  NAND2_X1 U759 ( .A1(n736), .A2(n935), .ZN(n731) );
  NAND2_X1 U760 ( .A1(G117), .A2(n856), .ZN(n689) );
  NAND2_X1 U761 ( .A1(G129), .A2(n858), .ZN(n688) );
  NAND2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U763 ( .A1(G105), .A2(n852), .ZN(n690) );
  XNOR2_X1 U764 ( .A(n690), .B(KEYINPUT38), .ZN(n691) );
  XNOR2_X1 U765 ( .A(n691), .B(KEYINPUT93), .ZN(n692) );
  NOR2_X1 U766 ( .A1(n693), .A2(n692), .ZN(n695) );
  NAND2_X1 U767 ( .A1(n853), .A2(G141), .ZN(n694) );
  NAND2_X1 U768 ( .A1(n695), .A2(n694), .ZN(n864) );
  NAND2_X1 U769 ( .A1(G1996), .A2(n864), .ZN(n696) );
  XNOR2_X1 U770 ( .A(n696), .B(KEYINPUT94), .ZN(n705) );
  NAND2_X1 U771 ( .A1(G107), .A2(n856), .ZN(n698) );
  NAND2_X1 U772 ( .A1(G119), .A2(n858), .ZN(n697) );
  NAND2_X1 U773 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U774 ( .A1(n852), .A2(G95), .ZN(n699) );
  XOR2_X1 U775 ( .A(KEYINPUT92), .B(n699), .Z(n700) );
  NOR2_X1 U776 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U777 ( .A1(n853), .A2(G131), .ZN(n702) );
  NAND2_X1 U778 ( .A1(n703), .A2(n702), .ZN(n865) );
  NAND2_X1 U779 ( .A1(G1991), .A2(n865), .ZN(n704) );
  NAND2_X1 U780 ( .A1(n705), .A2(n704), .ZN(n932) );
  NAND2_X1 U781 ( .A1(n736), .A2(n932), .ZN(n706) );
  XNOR2_X1 U782 ( .A(KEYINPUT95), .B(n706), .ZN(n728) );
  INV_X1 U783 ( .A(n728), .ZN(n707) );
  AND2_X1 U784 ( .A1(n731), .A2(n707), .ZN(n719) );
  AND2_X1 U785 ( .A1(n949), .A2(n719), .ZN(n708) );
  NAND2_X1 U786 ( .A1(n709), .A2(n708), .ZN(n723) );
  NOR2_X1 U787 ( .A1(G2090), .A2(G303), .ZN(n710) );
  NAND2_X1 U788 ( .A1(G8), .A2(n710), .ZN(n711) );
  NAND2_X1 U789 ( .A1(n712), .A2(n711), .ZN(n714) );
  AND2_X1 U790 ( .A1(n717), .A2(n719), .ZN(n713) );
  AND2_X1 U791 ( .A1(n714), .A2(n713), .ZN(n721) );
  NOR2_X1 U792 ( .A1(G1981), .A2(G305), .ZN(n715) );
  XOR2_X1 U793 ( .A(n715), .B(KEYINPUT24), .Z(n716) );
  NOR2_X1 U794 ( .A1(n717), .A2(n716), .ZN(n718) );
  AND2_X1 U795 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U796 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U797 ( .A1(n723), .A2(n722), .ZN(n725) );
  XNOR2_X1 U798 ( .A(G1986), .B(G290), .ZN(n962) );
  NAND2_X1 U799 ( .A1(n962), .A2(n736), .ZN(n724) );
  NAND2_X1 U800 ( .A1(n725), .A2(n724), .ZN(n739) );
  NOR2_X1 U801 ( .A1(G1996), .A2(n864), .ZN(n927) );
  NOR2_X1 U802 ( .A1(G1986), .A2(G290), .ZN(n726) );
  NOR2_X1 U803 ( .A1(G1991), .A2(n865), .ZN(n930) );
  NOR2_X1 U804 ( .A1(n726), .A2(n930), .ZN(n727) );
  NOR2_X1 U805 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U806 ( .A1(n927), .A2(n729), .ZN(n730) );
  XNOR2_X1 U807 ( .A(KEYINPUT39), .B(n730), .ZN(n732) );
  NAND2_X1 U808 ( .A1(n732), .A2(n731), .ZN(n735) );
  AND2_X1 U809 ( .A1(n733), .A2(n869), .ZN(n734) );
  XOR2_X1 U810 ( .A(KEYINPUT104), .B(n734), .Z(n942) );
  NAND2_X1 U811 ( .A1(n735), .A2(n942), .ZN(n737) );
  NAND2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U814 ( .A(n740), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U815 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U816 ( .A(G57), .ZN(G237) );
  INV_X1 U817 ( .A(G132), .ZN(G219) );
  NAND2_X1 U818 ( .A1(G7), .A2(G661), .ZN(n741) );
  XNOR2_X1 U819 ( .A(n741), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U820 ( .A(G223), .ZN(n808) );
  NAND2_X1 U821 ( .A1(n808), .A2(G567), .ZN(n742) );
  XOR2_X1 U822 ( .A(KEYINPUT11), .B(n742), .Z(G234) );
  INV_X1 U823 ( .A(G860), .ZN(n748) );
  NOR2_X1 U824 ( .A1(n748), .A2(n952), .ZN(n743) );
  XNOR2_X1 U825 ( .A(n743), .B(KEYINPUT73), .ZN(G153) );
  NAND2_X1 U826 ( .A1(G868), .A2(G301), .ZN(n745) );
  INV_X1 U827 ( .A(G868), .ZN(n790) );
  NAND2_X1 U828 ( .A1(n968), .A2(n790), .ZN(n744) );
  NAND2_X1 U829 ( .A1(n745), .A2(n744), .ZN(G284) );
  NAND2_X1 U830 ( .A1(G868), .A2(G286), .ZN(n747) );
  NAND2_X1 U831 ( .A1(G299), .A2(n790), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n747), .A2(n746), .ZN(G297) );
  NAND2_X1 U833 ( .A1(n748), .A2(G559), .ZN(n749) );
  INV_X1 U834 ( .A(n968), .ZN(n777) );
  NAND2_X1 U835 ( .A1(n749), .A2(n777), .ZN(n750) );
  XNOR2_X1 U836 ( .A(n750), .B(KEYINPUT80), .ZN(n751) );
  XNOR2_X1 U837 ( .A(KEYINPUT16), .B(n751), .ZN(G148) );
  NOR2_X1 U838 ( .A1(G868), .A2(n952), .ZN(n754) );
  NAND2_X1 U839 ( .A1(G868), .A2(n777), .ZN(n752) );
  NOR2_X1 U840 ( .A1(G559), .A2(n752), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n754), .A2(n753), .ZN(G282) );
  XNOR2_X1 U842 ( .A(G2100), .B(KEYINPUT83), .ZN(n765) );
  NAND2_X1 U843 ( .A1(G111), .A2(n856), .ZN(n755) );
  XNOR2_X1 U844 ( .A(n755), .B(KEYINPUT82), .ZN(n759) );
  XOR2_X1 U845 ( .A(KEYINPUT81), .B(KEYINPUT18), .Z(n757) );
  NAND2_X1 U846 ( .A1(G123), .A2(n858), .ZN(n756) );
  XNOR2_X1 U847 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n763) );
  NAND2_X1 U849 ( .A1(G99), .A2(n852), .ZN(n761) );
  NAND2_X1 U850 ( .A1(G135), .A2(n853), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n929) );
  XNOR2_X1 U853 ( .A(n929), .B(G2096), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(G156) );
  NAND2_X1 U855 ( .A1(n766), .A2(G67), .ZN(n769) );
  NAND2_X1 U856 ( .A1(G93), .A2(n767), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n770), .A2(G80), .ZN(n771) );
  XOR2_X1 U859 ( .A(KEYINPUT84), .B(n771), .Z(n772) );
  NOR2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n776) );
  NAND2_X1 U861 ( .A1(n774), .A2(G55), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n789) );
  NAND2_X1 U863 ( .A1(n777), .A2(G559), .ZN(n787) );
  XNOR2_X1 U864 ( .A(n952), .B(n787), .ZN(n778) );
  NOR2_X1 U865 ( .A1(n778), .A2(G860), .ZN(n779) );
  XNOR2_X1 U866 ( .A(n779), .B(KEYINPUT85), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n789), .B(n780), .ZN(G145) );
  XNOR2_X1 U868 ( .A(KEYINPUT19), .B(G305), .ZN(n781) );
  XNOR2_X1 U869 ( .A(n781), .B(n789), .ZN(n782) );
  XNOR2_X1 U870 ( .A(G166), .B(n782), .ZN(n785) );
  XNOR2_X1 U871 ( .A(G290), .B(G299), .ZN(n783) );
  XNOR2_X1 U872 ( .A(n783), .B(G288), .ZN(n784) );
  XNOR2_X1 U873 ( .A(n785), .B(n784), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n952), .B(n786), .ZN(n878) );
  XNOR2_X1 U875 ( .A(n787), .B(n878), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n788), .A2(G868), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(G295) );
  NAND2_X1 U879 ( .A1(G2078), .A2(G2084), .ZN(n793) );
  XOR2_X1 U880 ( .A(KEYINPUT20), .B(n793), .Z(n794) );
  NAND2_X1 U881 ( .A1(G2090), .A2(n794), .ZN(n795) );
  XNOR2_X1 U882 ( .A(KEYINPUT21), .B(n795), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n796), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U884 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U885 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U886 ( .A1(G219), .A2(G220), .ZN(n797) );
  XOR2_X1 U887 ( .A(KEYINPUT22), .B(n797), .Z(n798) );
  NOR2_X1 U888 ( .A1(G218), .A2(n798), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G96), .A2(n799), .ZN(n813) );
  NAND2_X1 U890 ( .A1(G2106), .A2(n813), .ZN(n803) );
  NAND2_X1 U891 ( .A1(G69), .A2(G120), .ZN(n800) );
  NOR2_X1 U892 ( .A1(G237), .A2(n800), .ZN(n801) );
  NAND2_X1 U893 ( .A1(G108), .A2(n801), .ZN(n814) );
  NAND2_X1 U894 ( .A1(G567), .A2(n814), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U896 ( .A(KEYINPUT89), .B(n804), .ZN(G319) );
  INV_X1 U897 ( .A(G319), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G661), .A2(G483), .ZN(n805) );
  XNOR2_X1 U899 ( .A(KEYINPUT90), .B(n805), .ZN(n806) );
  NOR2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n812), .A2(G36), .ZN(G176) );
  NAND2_X1 U902 ( .A1(G2106), .A2(n808), .ZN(G217) );
  NAND2_X1 U903 ( .A1(G15), .A2(G2), .ZN(n809) );
  XNOR2_X1 U904 ( .A(KEYINPUT107), .B(n809), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n810), .A2(G661), .ZN(G259) );
  NAND2_X1 U906 ( .A1(G3), .A2(G1), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(G188) );
  XOR2_X1 U908 ( .A(G96), .B(KEYINPUT108), .Z(G221) );
  INV_X1 U910 ( .A(G120), .ZN(G236) );
  INV_X1 U911 ( .A(G69), .ZN(G235) );
  NOR2_X1 U912 ( .A1(n814), .A2(n813), .ZN(G325) );
  INV_X1 U913 ( .A(G325), .ZN(G261) );
  XOR2_X1 U914 ( .A(KEYINPUT109), .B(G2090), .Z(n816) );
  XNOR2_X1 U915 ( .A(G2072), .B(G2078), .ZN(n815) );
  XNOR2_X1 U916 ( .A(n816), .B(n815), .ZN(n817) );
  XOR2_X1 U917 ( .A(n817), .B(G2096), .Z(n819) );
  XNOR2_X1 U918 ( .A(G2067), .B(G2084), .ZN(n818) );
  XNOR2_X1 U919 ( .A(n819), .B(n818), .ZN(n823) );
  XOR2_X1 U920 ( .A(G2100), .B(KEYINPUT43), .Z(n821) );
  XNOR2_X1 U921 ( .A(KEYINPUT42), .B(G2678), .ZN(n820) );
  XNOR2_X1 U922 ( .A(n821), .B(n820), .ZN(n822) );
  XOR2_X1 U923 ( .A(n823), .B(n822), .Z(G227) );
  XNOR2_X1 U924 ( .A(G1996), .B(KEYINPUT110), .ZN(n833) );
  XOR2_X1 U925 ( .A(G1981), .B(G1961), .Z(n825) );
  XNOR2_X1 U926 ( .A(G1991), .B(G1966), .ZN(n824) );
  XNOR2_X1 U927 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U928 ( .A(G1976), .B(G1971), .Z(n827) );
  XNOR2_X1 U929 ( .A(G1986), .B(G1956), .ZN(n826) );
  XNOR2_X1 U930 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U931 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U932 ( .A(G2474), .B(KEYINPUT41), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(G229) );
  NAND2_X1 U935 ( .A1(G124), .A2(n858), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n834), .B(KEYINPUT44), .ZN(n837) );
  NAND2_X1 U937 ( .A1(G112), .A2(n856), .ZN(n835) );
  XOR2_X1 U938 ( .A(KEYINPUT111), .B(n835), .Z(n836) );
  NAND2_X1 U939 ( .A1(n837), .A2(n836), .ZN(n841) );
  NAND2_X1 U940 ( .A1(G100), .A2(n852), .ZN(n839) );
  NAND2_X1 U941 ( .A1(G136), .A2(n853), .ZN(n838) );
  NAND2_X1 U942 ( .A1(n839), .A2(n838), .ZN(n840) );
  NOR2_X1 U943 ( .A1(n841), .A2(n840), .ZN(G162) );
  NAND2_X1 U944 ( .A1(G118), .A2(n856), .ZN(n850) );
  XNOR2_X1 U945 ( .A(KEYINPUT113), .B(KEYINPUT45), .ZN(n845) );
  NAND2_X1 U946 ( .A1(G106), .A2(n852), .ZN(n843) );
  NAND2_X1 U947 ( .A1(G142), .A2(n853), .ZN(n842) );
  NAND2_X1 U948 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U949 ( .A(n845), .B(n844), .ZN(n848) );
  NAND2_X1 U950 ( .A1(n858), .A2(G130), .ZN(n846) );
  XOR2_X1 U951 ( .A(KEYINPUT112), .B(n846), .Z(n847) );
  NOR2_X1 U952 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U953 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n851), .B(n929), .ZN(n868) );
  NAND2_X1 U955 ( .A1(G103), .A2(n852), .ZN(n855) );
  NAND2_X1 U956 ( .A1(G139), .A2(n853), .ZN(n854) );
  NAND2_X1 U957 ( .A1(n855), .A2(n854), .ZN(n863) );
  NAND2_X1 U958 ( .A1(n856), .A2(G115), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n857), .B(KEYINPUT114), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G127), .A2(n858), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(KEYINPUT47), .B(n861), .Z(n862) );
  NOR2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n921) );
  XNOR2_X1 U964 ( .A(n921), .B(n864), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U966 ( .A(n868), .B(n867), .Z(n871) );
  XOR2_X1 U967 ( .A(G160), .B(n869), .Z(n870) );
  XNOR2_X1 U968 ( .A(n871), .B(n870), .ZN(n876) );
  XOR2_X1 U969 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n873) );
  XNOR2_X1 U970 ( .A(G162), .B(KEYINPUT115), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U972 ( .A(G164), .B(n874), .Z(n875) );
  XNOR2_X1 U973 ( .A(n876), .B(n875), .ZN(n877) );
  NOR2_X1 U974 ( .A1(G37), .A2(n877), .ZN(G395) );
  XNOR2_X1 U975 ( .A(G171), .B(G286), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n880), .B(n968), .ZN(n881) );
  NOR2_X1 U978 ( .A1(G37), .A2(n881), .ZN(G397) );
  XNOR2_X1 U979 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n883) );
  NOR2_X1 U980 ( .A1(G227), .A2(G229), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n883), .B(n882), .ZN(n896) );
  XNOR2_X1 U982 ( .A(G2435), .B(G2443), .ZN(n893) );
  XOR2_X1 U983 ( .A(G2454), .B(G2430), .Z(n885) );
  XNOR2_X1 U984 ( .A(G2446), .B(KEYINPUT105), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U986 ( .A(G2451), .B(G2427), .Z(n887) );
  XNOR2_X1 U987 ( .A(G1341), .B(G1348), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U989 ( .A(n889), .B(n888), .Z(n891) );
  XNOR2_X1 U990 ( .A(KEYINPUT106), .B(G2438), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  NAND2_X1 U993 ( .A1(n894), .A2(G14), .ZN(n899) );
  NAND2_X1 U994 ( .A1(G319), .A2(n899), .ZN(n895) );
  NOR2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n898) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n897) );
  NAND2_X1 U997 ( .A1(n898), .A2(n897), .ZN(G225) );
  INV_X1 U998 ( .A(G225), .ZN(G308) );
  INV_X1 U999 ( .A(G108), .ZN(G238) );
  INV_X1 U1000 ( .A(n899), .ZN(G401) );
  XNOR2_X1 U1001 ( .A(G2067), .B(G26), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(G2072), .B(G33), .ZN(n900) );
  NOR2_X1 U1003 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U1004 ( .A1(G28), .A2(n902), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(G25), .B(G1991), .ZN(n903) );
  XNOR2_X1 U1006 ( .A(KEYINPUT120), .B(n903), .ZN(n904) );
  NOR2_X1 U1007 ( .A1(n905), .A2(n904), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n906), .B(G32), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(G27), .B(n907), .ZN(n908) );
  NOR2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n912), .B(KEYINPUT53), .ZN(n915) );
  XOR2_X1 U1013 ( .A(G2084), .B(G34), .Z(n913) );
  XNOR2_X1 U1014 ( .A(KEYINPUT54), .B(n913), .ZN(n914) );
  NAND2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(G35), .B(G2090), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1018 ( .A(KEYINPUT121), .B(n918), .Z(n919) );
  NOR2_X1 U1019 ( .A1(G29), .A2(n919), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n920), .B(KEYINPUT55), .ZN(n948) );
  XOR2_X1 U1021 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n945) );
  XNOR2_X1 U1022 ( .A(G2072), .B(n921), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(G164), .B(G2078), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(n922), .B(KEYINPUT118), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1026 ( .A(n925), .B(KEYINPUT50), .ZN(n941) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1029 ( .A(KEYINPUT51), .B(n928), .Z(n939) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n934) );
  XOR2_X1 U1031 ( .A(G160), .B(G2084), .Z(n931) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1035 ( .A(KEYINPUT117), .B(n937), .Z(n938) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(n945), .B(n944), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(G29), .A2(n946), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n1003) );
  XNOR2_X1 U1042 ( .A(G1966), .B(G168), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(KEYINPUT57), .B(n951), .ZN(n967) );
  XOR2_X1 U1045 ( .A(n952), .B(G1341), .Z(n954) );
  XNOR2_X1 U1046 ( .A(G171), .B(G1961), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n965) );
  NAND2_X1 U1048 ( .A1(G1971), .A2(G303), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(G1956), .B(G299), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1054 ( .A(KEYINPUT122), .B(n963), .Z(n964) );
  NOR2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n970) );
  XNOR2_X1 U1057 ( .A(G1348), .B(n968), .ZN(n969) );
  NOR2_X1 U1058 ( .A1(n970), .A2(n969), .ZN(n972) );
  XOR2_X1 U1059 ( .A(KEYINPUT56), .B(G16), .Z(n971) );
  NOR2_X1 U1060 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1061 ( .A(KEYINPUT123), .B(n973), .Z(n1000) );
  XOR2_X1 U1062 ( .A(G1986), .B(G24), .Z(n975) );
  XOR2_X1 U1063 ( .A(G1971), .B(G22), .Z(n974) );
  NAND2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(G23), .B(G1976), .ZN(n976) );
  NOR2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1067 ( .A(KEYINPUT58), .B(n978), .Z(n995) );
  XOR2_X1 U1068 ( .A(G1961), .B(G5), .Z(n990) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(G1981), .B(G6), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(KEYINPUT124), .B(n981), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(n982), .B(G20), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1075 ( .A(KEYINPUT59), .B(G1348), .Z(n985) );
  XNOR2_X1 U1076 ( .A(G4), .B(n985), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(KEYINPUT60), .B(n988), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G21), .B(G1966), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(KEYINPUT125), .B(n993), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1084 ( .A(KEYINPUT61), .B(n996), .Z(n997) );
  NOR2_X1 U1085 ( .A1(G16), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(KEYINPUT126), .B(n998), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1001), .B(KEYINPUT127), .ZN(n1002) );
  NOR2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(G11), .ZN(n1005) );
  XOR2_X1 U1091 ( .A(KEYINPUT62), .B(n1005), .Z(G311) );
  INV_X1 U1092 ( .A(G311), .ZN(G150) );
endmodule

