//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n202), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n210), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n213), .B1(new_n216), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT64), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G68), .Z(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND2_X1  g0043(.A1(new_n209), .A2(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n214), .ZN(new_n245));
  INV_X1    g0045(.A(G13), .ZN(new_n246));
  NOR3_X1   g0046(.A1(new_n246), .A2(new_n208), .A3(G1), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n249), .B1(new_n207), .B2(G20), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n248), .A2(new_n250), .B1(new_n249), .B2(new_n247), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n208), .A2(new_n252), .A3(KEYINPUT69), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G20), .B2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G150), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n252), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n257), .B(new_n258), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n245), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n251), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT9), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(KEYINPUT71), .A3(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n266), .A2(KEYINPUT71), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(KEYINPUT71), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n214), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n252), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n279), .A2(G223), .B1(new_n282), .B2(G77), .ZN(new_n283));
  INV_X1    g0083(.A(G222), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT68), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n274), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n288), .B1(new_n287), .B2(new_n286), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT67), .B1(new_n272), .B2(new_n214), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT67), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n291), .A2(new_n292), .A3(G1), .A4(G13), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(G274), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(KEYINPUT65), .A2(G45), .ZN(new_n295));
  NOR2_X1   g0095(.A1(KEYINPUT65), .A2(G45), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n295), .A2(new_n296), .A3(G41), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT66), .B1(new_n297), .B2(G1), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT65), .ZN(new_n299));
  INV_X1    g0099(.A(G45), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G41), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT65), .A2(G45), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT66), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(new_n207), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n294), .B1(new_n298), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n290), .A2(new_n293), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(G226), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n289), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  INV_X1    g0112(.A(G200), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n289), .B2(new_n310), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT72), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n271), .B1(new_n311), .B2(new_n312), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT10), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n311), .A2(new_n312), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n270), .B2(new_n267), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n314), .A2(new_n315), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n317), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n265), .B1(new_n311), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n289), .A2(new_n328), .A3(new_n310), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  AND4_X1   g0131(.A1(G232), .A2(new_n290), .A3(new_n293), .A4(new_n308), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT77), .B1(new_n307), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n290), .A2(G274), .A3(new_n293), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n304), .A2(new_n305), .A3(new_n207), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n305), .B1(new_n304), .B2(new_n207), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT77), .ZN(new_n338));
  INV_X1    g0138(.A(new_n332), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n277), .A2(new_n278), .ZN(new_n341));
  INV_X1    g0141(.A(G226), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G1698), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n341), .B(new_n343), .C1(G223), .C2(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G87), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n274), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n333), .A2(new_n340), .A3(new_n328), .A4(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n215), .B1(new_n209), .B2(G33), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n341), .A2(new_n350), .A3(G20), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT7), .B1(new_n282), .B2(new_n208), .ZN(new_n352));
  OAI21_X1  g0152(.A(G68), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n256), .A2(G159), .ZN(new_n354));
  INV_X1    g0154(.A(G58), .ZN(new_n355));
  INV_X1    g0155(.A(G68), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n357), .B2(new_n201), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n353), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n350), .B1(new_n341), .B2(G20), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n356), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT16), .B1(new_n365), .B2(new_n359), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n349), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n261), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n207), .A2(G20), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n248), .A2(new_n371), .B1(new_n247), .B2(new_n261), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n348), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n337), .A2(new_n339), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n346), .B1(new_n375), .B2(KEYINPUT77), .ZN(new_n376));
  AOI21_X1  g0176(.A(G169), .B1(new_n376), .B2(new_n340), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT18), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT17), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n333), .A2(new_n340), .A3(G190), .A4(new_n347), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n361), .B1(new_n353), .B2(new_n360), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n365), .A2(KEYINPUT16), .A3(new_n359), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n245), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n383), .A3(new_n372), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n313), .B1(new_n376), .B2(new_n340), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n379), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(new_n372), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n333), .A2(new_n340), .A3(new_n347), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n326), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n387), .A2(new_n389), .A3(new_n390), .A4(new_n348), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n367), .A2(new_n373), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(G200), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT17), .A4(new_n380), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n378), .A2(new_n386), .A3(new_n391), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n309), .A2(G244), .ZN(new_n396));
  NOR2_X1   g0196(.A1(G232), .A2(G1698), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n275), .A2(G238), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n341), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(new_n273), .C1(G107), .C2(new_n341), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n337), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n312), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n248), .A2(G77), .A3(new_n369), .ZN(new_n403));
  INV_X1    g0203(.A(new_n247), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT15), .B(G87), .ZN(new_n405));
  INV_X1    g0205(.A(G77), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n405), .A2(new_n260), .B1(new_n208), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n256), .B2(new_n368), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n403), .B1(G77), .B2(new_n404), .C1(new_n408), .C2(new_n349), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(G200), .B2(new_n401), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n402), .B1(new_n410), .B2(KEYINPUT70), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(KEYINPUT70), .B2(new_n410), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n401), .A2(new_n326), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n409), .B(new_n413), .C1(G179), .C2(new_n401), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n331), .A2(new_n395), .A3(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n290), .A2(G238), .A3(new_n293), .A4(new_n308), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G226), .A2(G1698), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n228), .B2(G1698), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n419), .B1(new_n421), .B2(new_n341), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n417), .B1(new_n422), .B2(new_n274), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n307), .A2(new_n423), .A3(KEYINPUT13), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n342), .A2(new_n275), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n228), .A2(G1698), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n426), .B(new_n427), .C1(new_n280), .C2(new_n281), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n418), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n309), .A2(G238), .B1(new_n429), .B2(new_n273), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n425), .B1(new_n430), .B2(new_n337), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G190), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT13), .B1(new_n307), .B2(new_n423), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n337), .A3(new_n425), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G200), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n248), .A2(G68), .A3(new_n369), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n247), .A2(new_n356), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT12), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n256), .A2(G50), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n259), .A2(G77), .B1(G20), .B2(new_n356), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n245), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT11), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n438), .B(new_n440), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n445), .B2(new_n444), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n433), .A2(new_n437), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT73), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n433), .A2(KEYINPUT73), .A3(new_n437), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(G169), .B1(new_n424), .B2(new_n431), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n454), .A2(KEYINPUT14), .B1(new_n432), .B2(G179), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n326), .B1(new_n434), .B2(new_n435), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT74), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT14), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n457), .B1(new_n456), .B2(new_n458), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT75), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n436), .A2(new_n458), .A3(G169), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT74), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(KEYINPUT75), .A3(new_n455), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n447), .B(KEYINPUT76), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n453), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n416), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT21), .ZN(new_n474));
  OAI211_X1 g0274(.A(G264), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(new_n275), .C1(new_n280), .C2(new_n281), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n277), .A2(G303), .A3(new_n278), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n273), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(KEYINPUT82), .A3(new_n273), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n207), .A2(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(G274), .A3(new_n290), .A4(new_n293), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n300), .A2(G1), .ZN(new_n490));
  INV_X1    g0290(.A(new_n487), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n485), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(new_n290), .A3(G270), .A4(new_n293), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n483), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(G20), .B1(G33), .B2(G283), .ZN(new_n496));
  INV_X1    g0296(.A(G97), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(G33), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G116), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G20), .ZN(new_n500));
  AND4_X1   g0300(.A1(KEYINPUT20), .A2(new_n245), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n244), .A2(new_n214), .B1(G20), .B2(new_n499), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT20), .B1(new_n502), .B2(new_n498), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n247), .A2(new_n499), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n207), .A2(G33), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n349), .A2(new_n404), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n507), .B2(new_n499), .ZN(new_n508));
  OAI21_X1  g0308(.A(G169), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n474), .B1(new_n495), .B2(new_n509), .ZN(new_n510));
  OAI221_X1 g0310(.A(new_n505), .B1(new_n499), .B2(new_n507), .C1(new_n501), .C2(new_n503), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n489), .A2(G179), .A3(new_n493), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n483), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n483), .A2(new_n494), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n511), .A2(new_n514), .A3(KEYINPUT21), .A4(G169), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n510), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n511), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n483), .A2(G190), .A3(new_n494), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n517), .B(new_n518), .C1(new_n495), .C2(new_n313), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n252), .A2(new_n499), .ZN(new_n522));
  AOI21_X1  g0322(.A(G1698), .B1(new_n277), .B2(new_n278), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(G238), .ZN(new_n524));
  OAI211_X1 g0324(.A(G244), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n274), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT81), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n290), .A2(G274), .A3(new_n490), .A4(new_n293), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n290), .A2(G250), .A3(new_n484), .A4(new_n293), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n528), .A2(new_n529), .ZN(new_n532));
  INV_X1    g0332(.A(new_n522), .ZN(new_n533));
  INV_X1    g0333(.A(G238), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n525), .B(new_n533), .C1(new_n285), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n273), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT81), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n326), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n527), .B1(new_n526), .B2(new_n530), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n532), .A2(new_n536), .A3(KEYINPUT81), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n328), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(G20), .B1(new_n277), .B2(new_n278), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G68), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT19), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n260), .B2(new_n497), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n208), .B1(new_n418), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G87), .B2(new_n205), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(new_n245), .B1(new_n247), .B2(new_n405), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n507), .B2(new_n405), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n538), .A2(new_n541), .A3(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n542), .A2(new_n552), .A3(G87), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n208), .B(G87), .C1(new_n280), .C2(new_n281), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT22), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT24), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n208), .B2(G107), .ZN(new_n559));
  INV_X1    g0359(.A(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(KEYINPUT23), .A3(G20), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n559), .A2(new_n561), .B1(new_n522), .B2(new_n208), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n556), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n557), .B1(new_n556), .B2(new_n562), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n245), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n507), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT25), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n404), .B2(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n560), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n567), .A2(G107), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n341), .A2(G257), .A3(G1698), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G294), .ZN(new_n573));
  OAI211_X1 g0373(.A(G250), .B(new_n275), .C1(new_n280), .C2(new_n281), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n492), .A2(new_n290), .A3(new_n293), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n273), .A2(new_n575), .B1(new_n576), .B2(G264), .ZN(new_n577));
  AOI21_X1  g0377(.A(G200), .B1(new_n577), .B2(new_n489), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n273), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(G264), .ZN(new_n580));
  AND4_X1   g0380(.A1(new_n312), .A2(new_n579), .A3(new_n580), .A4(new_n489), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n566), .B(new_n571), .C1(new_n578), .C2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(G200), .B1(new_n531), .B2(new_n537), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n539), .A2(G190), .A3(new_n540), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n567), .A2(G87), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n549), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n577), .A2(new_n328), .A3(new_n489), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n579), .A2(new_n580), .A3(new_n489), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n326), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n552), .B1(new_n542), .B2(G87), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n554), .A2(KEYINPUT22), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n562), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT24), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n349), .B1(new_n594), .B2(new_n563), .ZN(new_n595));
  INV_X1    g0395(.A(new_n571), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n588), .B(new_n590), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n551), .A2(new_n582), .A3(new_n587), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(G244), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT79), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT79), .ZN(new_n601));
  OAI211_X1 g0401(.A(KEYINPUT4), .B(new_n600), .C1(new_n523), .C2(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n279), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT4), .ZN(new_n604));
  OAI211_X1 g0404(.A(KEYINPUT79), .B(new_n604), .C1(new_n285), .C2(new_n599), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n273), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n492), .A2(new_n290), .A3(G257), .A4(new_n293), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n489), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n326), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT6), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n497), .A2(new_n560), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n204), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n560), .A2(KEYINPUT6), .A3(G97), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n618));
  OAI21_X1  g0418(.A(G107), .B1(new_n351), .B2(new_n352), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n245), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n247), .A2(new_n497), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT78), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(G97), .B2(new_n567), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n609), .B1(new_n606), .B2(new_n273), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n328), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n612), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n611), .A2(KEYINPUT80), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT80), .ZN(new_n630));
  OAI21_X1  g0430(.A(G200), .B1(new_n626), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n621), .B(new_n624), .C1(new_n611), .C2(new_n312), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n598), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n473), .A2(new_n521), .A3(new_n635), .ZN(G372));
  AND3_X1   g0436(.A1(new_n612), .A2(new_n625), .A3(new_n627), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n551), .A3(new_n587), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n526), .A2(new_n530), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n541), .B(new_n550), .C1(G169), .C2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n584), .B(new_n586), .C1(new_n313), .C2(new_n640), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n637), .A2(new_n642), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n639), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT83), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n639), .A2(KEYINPUT83), .A3(new_n644), .A4(new_n641), .ZN(new_n648));
  INV_X1    g0448(.A(new_n516), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n597), .ZN(new_n650));
  INV_X1    g0450(.A(new_n634), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n641), .A2(new_n643), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n650), .A2(new_n651), .A3(new_n582), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n473), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT84), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n467), .A2(KEYINPUT75), .A3(new_n455), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT75), .B1(new_n467), .B2(new_n455), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n470), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n453), .B2(new_n414), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n386), .A3(new_n394), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n378), .A2(new_n391), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n663), .A2(new_n325), .B1(new_n329), .B2(new_n327), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n656), .A2(new_n664), .ZN(G369));
  NAND2_X1  g0465(.A1(new_n582), .A2(new_n597), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n246), .A2(G1), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n208), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(G213), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n595), .B2(new_n596), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n597), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n676), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n676), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n521), .B1(new_n517), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n516), .A2(new_n511), .A3(new_n676), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(KEYINPUT86), .B(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT87), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT87), .ZN(new_n690));
  AOI211_X1 g0490(.A(new_n690), .B(new_n687), .C1(new_n684), .C2(new_n685), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n682), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n516), .A2(new_n683), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n694), .A2(new_n666), .B1(new_n597), .B2(new_n676), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n693), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n211), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G1), .A3(new_n700), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n701), .A2(KEYINPUT88), .B1(new_n217), .B2(new_n699), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(KEYINPUT88), .B2(new_n701), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT28), .Z(new_n704));
  NAND3_X1  g0504(.A1(new_n635), .A2(new_n521), .A3(new_n683), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT91), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n539), .A2(new_n540), .A3(new_n577), .ZN(new_n708));
  INV_X1    g0508(.A(new_n482), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT82), .B1(new_n478), .B2(new_n273), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n512), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT89), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n483), .A2(KEYINPUT89), .A3(new_n512), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n708), .A2(new_n626), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n716), .B(new_n609), .C1(new_n606), .C2(new_n273), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n708), .A2(new_n714), .A3(new_n713), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT90), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n589), .B(new_n328), .C1(new_n526), .C2(new_n530), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n495), .A2(new_n721), .A3(new_n626), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT89), .B1(new_n483), .B2(new_n512), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n539), .A2(new_n540), .A3(new_n577), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT90), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n714), .A4(new_n718), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n717), .A2(new_n720), .A3(new_n723), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n635), .A2(KEYINPUT91), .A3(new_n521), .A4(new_n683), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n707), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n720), .A2(new_n728), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n722), .B1(new_n716), .B2(new_n715), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n683), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(KEYINPUT31), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n688), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n652), .A2(new_n637), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT26), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n653), .A2(new_n739), .A3(new_n741), .A4(new_n641), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n683), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n654), .A2(new_n683), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n745), .A2(KEYINPUT29), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n738), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n704), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR2_X1   g0549(.A1(new_n246), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n207), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n698), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT92), .Z(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n214), .B1(G20), .B2(new_n326), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n208), .B1(new_n758), .B2(G190), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n497), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n312), .A2(new_n313), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n208), .A2(G179), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G87), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n282), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT95), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n208), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n758), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n208), .A2(new_n328), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n313), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n767), .B(new_n772), .C1(new_n356), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n328), .A2(G200), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(G20), .A3(G190), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n768), .A2(new_n781), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n355), .B1(new_n783), .B2(new_n406), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n773), .A2(new_n761), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n774), .A2(new_n762), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n249), .B1(new_n786), .B2(new_n560), .ZN(new_n787));
  OR4_X1    g0587(.A1(new_n760), .A2(new_n780), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n782), .A2(new_n789), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n785), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n341), .B(new_n791), .C1(G326), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n779), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT33), .B(G317), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n759), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G294), .ZN(new_n798));
  INV_X1    g0598(.A(G303), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n763), .A2(new_n799), .B1(new_n783), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n769), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G329), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n793), .A2(new_n796), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n757), .B1(new_n788), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT94), .Z(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n756), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n697), .A2(new_n341), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n301), .A2(new_n303), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n217), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT93), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT93), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n300), .C2(new_n242), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n697), .A2(new_n282), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n816), .A2(G355), .B1(new_n499), .B2(new_n697), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n755), .B(new_n805), .C1(new_n809), .C2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT97), .Z(new_n820));
  INV_X1    g0620(.A(new_n808), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n686), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT98), .ZN(new_n823));
  INV_X1    g0623(.A(new_n689), .ZN(new_n824));
  INV_X1    g0624(.A(new_n691), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n686), .A2(new_n688), .B1(new_n698), .B2(new_n752), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(G396));
  NOR2_X1   g0628(.A1(new_n676), .A2(new_n414), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n676), .A2(new_n409), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n412), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n829), .B1(new_n831), .B2(new_n414), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n654), .A2(new_n683), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n414), .ZN(new_n834));
  INV_X1    g0634(.A(new_n829), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT101), .ZN(new_n837));
  INV_X1    g0637(.A(new_n745), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n753), .B1(new_n839), .B2(new_n738), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n738), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n756), .A2(new_n806), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT99), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n754), .B1(G77), .B2(new_n843), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n764), .A2(new_n786), .B1(new_n783), .B2(new_n499), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G303), .B2(new_n792), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n782), .A2(new_n847), .B1(new_n769), .B2(new_n800), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n282), .B1(new_n763), .B2(new_n560), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n848), .A2(new_n849), .A3(new_n760), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n779), .B(KEYINPUT100), .Z(new_n851));
  OAI211_X1 g0651(.A(new_n846), .B(new_n850), .C1(new_n851), .C2(new_n790), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n341), .B1(new_n786), .B2(new_n356), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n763), .A2(new_n249), .B1(new_n769), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(G58), .C2(new_n797), .ZN(new_n856));
  INV_X1    g0656(.A(new_n782), .ZN(new_n857));
  INV_X1    g0657(.A(new_n783), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n857), .A2(G143), .B1(new_n858), .B2(G159), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  INV_X1    g0660(.A(G150), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n859), .B1(new_n860), .B2(new_n785), .C1(new_n779), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT34), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n856), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n862), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(KEYINPUT34), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n852), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n844), .B1(new_n867), .B2(new_n756), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n832), .B2(new_n807), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n841), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G384));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n673), .B1(new_n367), .B2(new_n373), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n374), .B2(new_n377), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n384), .A2(new_n385), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n387), .A2(new_n389), .A3(new_n348), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n392), .A2(new_n393), .A3(new_n380), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n873), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(KEYINPUT103), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n873), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n395), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT103), .B1(new_n876), .B2(new_n880), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n872), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n876), .A2(new_n880), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT103), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n883), .A4(new_n881), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n886), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n659), .A2(new_n676), .ZN(new_n892));
  INV_X1    g0692(.A(new_n890), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT104), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n876), .B2(new_n880), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n877), .A2(new_n878), .A3(new_n873), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT104), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n895), .A2(KEYINPUT105), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT105), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n883), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n893), .B1(new_n900), .B2(new_n872), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n891), .B(new_n892), .C1(new_n901), .C2(KEYINPUT39), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n662), .A2(new_n673), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n470), .A2(new_n676), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n659), .A2(new_n452), .A3(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n470), .B(new_n676), .C1(new_n469), .C2(new_n453), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n835), .B2(new_n833), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n886), .A2(new_n890), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n902), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n746), .A2(new_n744), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n473), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n664), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n911), .B(new_n914), .Z(new_n915));
  NAND2_X1  g0715(.A1(new_n899), .A2(new_n883), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n895), .A2(KEYINPUT105), .A3(new_n897), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n872), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n890), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n731), .A2(new_n730), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT106), .B1(new_n735), .B2(KEYINPUT31), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n729), .A2(new_n676), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT106), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT31), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n920), .A2(new_n921), .A3(new_n707), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n836), .B1(new_n905), .B2(new_n906), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT40), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n909), .A2(new_n926), .A3(new_n927), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n919), .A2(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n473), .A2(new_n926), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n688), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n931), .B2(new_n932), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n915), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n915), .A2(new_n934), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n935), .B(new_n936), .C1(new_n207), .C2(new_n750), .ZN(new_n937));
  OAI21_X1  g0737(.A(G77), .B1(new_n355), .B2(new_n356), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n217), .A2(new_n938), .B1(G50), .B2(new_n356), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(G1), .A3(new_n246), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT102), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n499), .B(new_n216), .C1(new_n617), .C2(KEYINPUT35), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(KEYINPUT35), .B2(new_n617), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT36), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n944), .B2(new_n943), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n937), .A2(new_n946), .ZN(G367));
  NAND2_X1  g0747(.A1(new_n676), .A2(new_n625), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n651), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n637), .A2(new_n676), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n694), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(new_n667), .A3(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n679), .B1(new_n632), .B2(new_n633), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n676), .B1(new_n955), .B2(new_n628), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n953), .B2(KEYINPUT42), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n683), .A2(new_n586), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n652), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n641), .B2(new_n958), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n954), .A2(new_n957), .B1(KEYINPUT43), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n693), .A2(new_n951), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n698), .B(KEYINPUT41), .Z(new_n966));
  INV_X1    g0766(.A(new_n951), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n967), .A2(new_n968), .A3(new_n695), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n967), .B2(new_n695), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n967), .A2(new_n695), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n967), .A2(KEYINPUT44), .A3(new_n695), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n692), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(KEYINPUT107), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n971), .A2(new_n976), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n693), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n681), .A2(new_n694), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n952), .A2(new_n667), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n824), .A2(new_n825), .A3(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n983), .B(new_n982), .C1(new_n689), .C2(new_n691), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n979), .A2(KEYINPUT107), .A3(new_n693), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n981), .A2(new_n748), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n966), .B1(new_n990), .B2(new_n748), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n965), .B1(new_n991), .B2(new_n752), .ZN(new_n992));
  INV_X1    g0792(.A(new_n810), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n809), .B1(new_n211), .B2(new_n405), .C1(new_n993), .C2(new_n234), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n763), .A2(new_n499), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT46), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n759), .A2(new_n560), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n786), .A2(new_n497), .ZN(new_n998));
  NOR4_X1   g0798(.A1(new_n996), .A2(new_n341), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n782), .A2(new_n799), .B1(new_n783), .B2(new_n790), .ZN(new_n1000));
  INV_X1    g0800(.A(G317), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n785), .A2(new_n800), .B1(new_n769), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n999), .B(new_n1003), .C1(new_n851), .C2(new_n847), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n858), .A2(G50), .B1(new_n802), .B2(G137), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n861), .B2(new_n782), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n759), .A2(new_n356), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n341), .B1(new_n786), .B2(new_n406), .ZN(new_n1008));
  INV_X1    g0808(.A(G143), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n785), .A2(new_n1009), .B1(new_n763), .B2(new_n355), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n851), .B2(new_n770), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1004), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT47), .Z(new_n1014));
  OAI211_X1 g0814(.A(new_n754), .B(new_n994), .C1(new_n1014), .C2(new_n757), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT108), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n821), .B2(new_n960), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n992), .A2(new_n1017), .ZN(G387));
  INV_X1    g0818(.A(new_n231), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n993), .B1(new_n1019), .B2(new_n811), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n700), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n816), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n700), .B(new_n300), .C1(new_n356), .C2(new_n406), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT50), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n261), .B2(G50), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n368), .A2(KEYINPUT50), .A3(new_n249), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1022), .A2(new_n1027), .B1(G107), .B2(new_n211), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n755), .B1(new_n1028), .B2(new_n809), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n682), .B2(new_n821), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n802), .A2(G326), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n786), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n341), .B1(new_n1032), .B2(G116), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n763), .A2(new_n847), .B1(new_n759), .B2(new_n790), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G322), .A2(new_n792), .B1(new_n858), .B2(G303), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n1001), .B2(new_n782), .C1(new_n851), .C2(new_n800), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n1037), .B2(new_n1036), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT49), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1031), .B(new_n1033), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n779), .A2(new_n261), .B1(new_n356), .B2(new_n783), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT109), .Z(new_n1044));
  AOI22_X1  g0844(.A1(new_n792), .A2(G159), .B1(new_n802), .B2(G150), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n249), .B2(new_n782), .C1(new_n406), .C2(new_n763), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n759), .A2(new_n405), .ZN(new_n1047));
  OR4_X1    g0847(.A1(new_n282), .A2(new_n1046), .A3(new_n998), .A4(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1041), .A2(new_n1042), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1030), .B1(new_n1049), .B2(new_n756), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n988), .B2(new_n752), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n988), .A2(new_n738), .A3(new_n744), .A4(new_n746), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n698), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n748), .A2(new_n988), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(G393));
  NAND2_X1  g0855(.A1(new_n980), .A2(new_n977), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(new_n751), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n967), .A2(new_n808), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n809), .B1(new_n497), .B2(new_n211), .C1(new_n993), .C2(new_n238), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n754), .A2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n783), .A2(new_n261), .B1(new_n769), .B2(new_n1009), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n341), .B1(new_n759), .B2(new_n406), .C1(new_n764), .C2(new_n786), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n763), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1061), .B(new_n1062), .C1(G68), .C2(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n861), .A2(new_n785), .B1(new_n782), .B2(new_n770), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1065), .B(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1064), .B(new_n1067), .C1(new_n851), .C2(new_n249), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT111), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n783), .A2(new_n847), .B1(new_n769), .B2(new_n789), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n282), .B1(new_n759), .B2(new_n499), .C1(new_n560), .C2(new_n786), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(G283), .C2(new_n1063), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1001), .A2(new_n785), .B1(new_n782), .B2(new_n800), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1072), .B(new_n1075), .C1(new_n851), .C2(new_n799), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1068), .A2(KEYINPUT111), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1069), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1060), .B1(new_n1078), .B2(new_n756), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1057), .B1(new_n1058), .B2(new_n1079), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1052), .A2(new_n1056), .A3(KEYINPUT113), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT113), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n990), .A2(new_n698), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(G390));
  OAI21_X1  g0885(.A(new_n891), .B1(new_n901), .B2(KEYINPUT39), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT114), .B1(new_n908), .B2(new_n892), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT114), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n892), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n833), .A2(new_n835), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1088), .B(new_n1089), .C1(new_n1090), .C2(new_n907), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1086), .A2(new_n1087), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n742), .A2(new_n683), .A3(new_n834), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(new_n835), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n919), .B(new_n1089), .C1(new_n907), .C2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n688), .B(new_n832), .C1(new_n732), .C2(new_n736), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1096), .A2(new_n907), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1092), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n926), .A2(G330), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n927), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n473), .A2(new_n1100), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n913), .A2(new_n664), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1097), .A2(new_n1094), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1100), .A2(new_n837), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1106), .B1(new_n907), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1096), .A2(new_n907), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1090), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1105), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1103), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n698), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1063), .A2(G150), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G128), .A2(new_n792), .B1(new_n857), .B2(G132), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n769), .C1(new_n783), .C2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1117), .B(new_n1121), .C1(G159), .C2(new_n797), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n341), .B1(new_n786), .B2(new_n249), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT115), .Z(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(new_n860), .C2(new_n851), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n782), .A2(new_n499), .B1(new_n759), .B2(new_n406), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT116), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n785), .A2(new_n790), .B1(new_n786), .B2(new_n356), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n783), .A2(new_n497), .B1(new_n769), .B2(new_n847), .ZN(new_n1129));
  NOR4_X1   g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n341), .A4(new_n765), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n851), .B2(new_n560), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1132), .A2(new_n756), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n754), .B1(new_n368), .B2(new_n843), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n807), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1133), .B(new_n1134), .C1(new_n1086), .C2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1103), .B2(new_n752), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1115), .A2(new_n1137), .ZN(G378));
  NAND2_X1  g0938(.A1(new_n1113), .A2(new_n1105), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n919), .A2(new_n928), .ZN(new_n1140));
  INV_X1    g0940(.A(G330), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n930), .B2(new_n929), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n674), .A2(new_n265), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n331), .A2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n319), .A2(new_n324), .B1(new_n329), .B2(new_n327), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1145), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1144), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n331), .A2(new_n1145), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n1143), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1140), .A2(new_n1142), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n902), .B(new_n910), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1154), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1140), .A2(new_n1142), .A3(new_n1154), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n911), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT57), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n699), .B1(new_n1139), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1105), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1108), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1110), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1167), .B1(new_n1103), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1162), .A2(KEYINPUT120), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT120), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1160), .A2(new_n911), .A3(new_n1173), .A4(new_n1161), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1172), .A2(KEYINPUT119), .A3(new_n1157), .A4(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1157), .A2(KEYINPUT119), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1173), .B1(new_n1177), .B2(new_n911), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1174), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1171), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1166), .B1(new_n1181), .B2(KEYINPUT57), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n752), .B(new_n698), .C1(new_n249), .C2(new_n842), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT118), .Z(new_n1185));
  NOR2_X1   g0985(.A1(new_n341), .A2(G41), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(G33), .A2(G41), .ZN(new_n1187));
  OR3_X1    g0987(.A1(new_n1186), .A2(G50), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1032), .A2(G58), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n560), .B2(new_n782), .C1(new_n405), .C2(new_n783), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1186), .B1(new_n790), .B2(new_n769), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n785), .A2(new_n499), .B1(new_n763), .B2(new_n406), .ZN(new_n1192));
  OR3_X1    g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n1007), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1190), .B(new_n1193), .C1(G97), .C2(new_n794), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1188), .B1(new_n1194), .B2(KEYINPUT58), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT117), .Z(new_n1196));
  NOR2_X1   g0996(.A1(new_n763), .A2(new_n1120), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n785), .A2(new_n1119), .B1(new_n783), .B2(new_n860), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(G128), .C2(new_n857), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n854), .B2(new_n779), .C1(new_n861), .C2(new_n759), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  INV_X1    g1001(.A(G124), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1187), .B1(new_n769), .B2(new_n1202), .C1(new_n770), .C2(new_n786), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1200), .B2(KEYINPUT59), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1201), .A2(new_n1204), .B1(new_n1194), .B2(KEYINPUT58), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1196), .A2(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1185), .B1(new_n757), .B2(new_n1206), .C1(new_n1159), .C2(new_n807), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1180), .A2(new_n1175), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n1209), .B2(new_n752), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1183), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(G375));
  NAND2_X1  g1013(.A1(new_n907), .A2(new_n806), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n754), .B1(G68), .B2(new_n843), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n858), .A2(G107), .B1(new_n802), .B2(G303), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n497), .B2(new_n763), .C1(new_n847), .C2(new_n785), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n341), .B(new_n1217), .C1(G77), .C2(new_n1032), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1047), .B1(G283), .B2(new_n857), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT121), .Z(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n499), .C2(new_n851), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n858), .A2(G150), .B1(new_n802), .B2(G128), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n770), .B2(new_n763), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G132), .A2(new_n792), .B1(new_n857), .B2(G137), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n341), .A3(new_n1189), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G50), .C2(new_n797), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n851), .B2(new_n1120), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1221), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1215), .B1(new_n1228), .B2(new_n756), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT122), .Z(new_n1230));
  AOI22_X1  g1030(.A1(new_n1170), .A2(new_n752), .B1(new_n1214), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n966), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1111), .A2(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1170), .A2(new_n1105), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1231), .B1(new_n1233), .B2(new_n1234), .ZN(G381));
  OR2_X1    g1035(.A1(new_n1212), .A2(KEYINPUT123), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1212), .A2(KEYINPUT123), .ZN(new_n1237));
  OR4_X1    g1037(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1238), .A2(G387), .A3(G378), .A4(G381), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .ZN(G407));
  INV_X1    g1040(.A(G378), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n675), .A2(G213), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1236), .A2(new_n1241), .A3(new_n1237), .A4(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1045(.A1(new_n1181), .A2(new_n1232), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1208), .B1(new_n1163), .B2(new_n752), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G378), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1139), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n698), .B1(new_n1171), .B2(new_n1164), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G378), .B(new_n1210), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT124), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1182), .A2(new_n1253), .A3(G378), .A4(new_n1210), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1248), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1111), .A2(KEYINPUT60), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n699), .B1(new_n1256), .B2(new_n1234), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1234), .B2(new_n1256), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1231), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n870), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(G384), .A3(new_n1231), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1255), .A2(new_n1262), .A3(new_n1243), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT125), .B1(new_n1263), .B2(KEYINPUT63), .ZN(new_n1264));
  AND3_X1   g1064(.A1(G390), .A2(new_n992), .A3(new_n1017), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G390), .B1(new_n992), .B2(new_n1017), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT126), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(G396), .B(G393), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1268), .B(KEYINPUT126), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT127), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1248), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1242), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1243), .A2(G2897), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1260), .A2(new_n1261), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1274), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1262), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1277), .A2(new_n1242), .A3(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1263), .A2(KEYINPUT63), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1264), .A2(new_n1283), .A3(new_n1288), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1277), .A2(new_n1292), .A3(new_n1242), .A4(new_n1284), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1282), .B1(new_n1255), .B2(new_n1243), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1271), .A3(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1263), .A2(new_n1292), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1291), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1290), .A2(new_n1297), .ZN(G405));
  AOI21_X1  g1098(.A(G378), .B1(new_n1182), .B2(new_n1210), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1275), .A2(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1291), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1284), .ZN(G402));
endmodule


