

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n388) );
  XNOR2_X1 U325 ( .A(KEYINPUT109), .B(KEYINPUT47), .ZN(n408) );
  XNOR2_X1 U326 ( .A(n409), .B(n408), .ZN(n416) );
  INV_X1 U327 ( .A(KEYINPUT48), .ZN(n417) );
  XNOR2_X1 U328 ( .A(n418), .B(n417), .ZN(n527) );
  INV_X1 U329 ( .A(G183GAT), .ZN(n453) );
  XNOR2_X1 U330 ( .A(n453), .B(KEYINPUT120), .ZN(n454) );
  XNOR2_X1 U331 ( .A(n455), .B(n454), .ZN(G1350GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n293) );
  XNOR2_X1 U333 ( .A(KEYINPUT80), .B(KEYINPUT12), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n311) );
  XOR2_X1 U335 ( .A(G22GAT), .B(G155GAT), .Z(n316) );
  XOR2_X1 U336 ( .A(n316), .B(G71GAT), .Z(n295) );
  XOR2_X1 U337 ( .A(G15GAT), .B(G127GAT), .Z(n442) );
  XNOR2_X1 U338 ( .A(G183GAT), .B(n442), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n307) );
  XOR2_X1 U340 ( .A(G64GAT), .B(G78GAT), .Z(n297) );
  XNOR2_X1 U341 ( .A(G8GAT), .B(G211GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U343 ( .A(KEYINPUT84), .B(KEYINPUT82), .Z(n299) );
  XNOR2_X1 U344 ( .A(KEYINPUT15), .B(KEYINPUT83), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U346 ( .A(n301), .B(n300), .Z(n305) );
  XNOR2_X1 U347 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n302), .B(KEYINPUT68), .ZN(n381) );
  XNOR2_X1 U349 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n303), .B(KEYINPUT70), .ZN(n391) );
  XNOR2_X1 U351 ( .A(n381), .B(n391), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(n307), .B(n306), .Z(n309) );
  NAND2_X1 U354 ( .A1(G231GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n582) );
  INV_X1 U357 ( .A(n582), .ZN(n482) );
  XOR2_X1 U358 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n313) );
  XNOR2_X1 U359 ( .A(G197GAT), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n315) );
  XOR2_X1 U361 ( .A(G218GAT), .B(KEYINPUT89), .Z(n314) );
  XOR2_X1 U362 ( .A(n315), .B(n314), .Z(n432) );
  XOR2_X1 U363 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n318) );
  XOR2_X1 U364 ( .A(G50GAT), .B(G162GAT), .Z(n365) );
  XNOR2_X1 U365 ( .A(n365), .B(n316), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n328) );
  XOR2_X1 U367 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n326) );
  XOR2_X1 U368 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n320) );
  XNOR2_X1 U369 ( .A(G78GAT), .B(G148GAT), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n322) );
  XOR2_X1 U371 ( .A(G106GAT), .B(G204GAT), .Z(n321) );
  XOR2_X1 U372 ( .A(n322), .B(n321), .Z(n401) );
  XOR2_X1 U373 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n324) );
  XNOR2_X1 U374 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n345) );
  XNOR2_X1 U376 ( .A(n401), .B(n345), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U378 ( .A(n328), .B(n327), .Z(n330) );
  NAND2_X1 U379 ( .A1(G228GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n432), .B(n331), .ZN(n462) );
  XOR2_X1 U382 ( .A(G162GAT), .B(G127GAT), .Z(n333) );
  XNOR2_X1 U383 ( .A(G29GAT), .B(G134GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U385 ( .A(G57GAT), .B(G155GAT), .Z(n335) );
  XNOR2_X1 U386 ( .A(G120GAT), .B(G148GAT), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U388 ( .A(n337), .B(n336), .Z(n342) );
  XOR2_X1 U389 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n339) );
  NAND2_X1 U390 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U392 ( .A(KEYINPUT93), .B(n340), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n342), .B(n341), .ZN(n351) );
  XOR2_X1 U394 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n344) );
  XNOR2_X1 U395 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n349) );
  XOR2_X1 U397 ( .A(KEYINPUT78), .B(G85GAT), .Z(n347) );
  XOR2_X1 U398 ( .A(G113GAT), .B(KEYINPUT0), .Z(n446) );
  XNOR2_X1 U399 ( .A(n446), .B(n345), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U401 ( .A(n349), .B(n348), .Z(n350) );
  XOR2_X1 U402 ( .A(n351), .B(n350), .Z(n516) );
  INV_X1 U403 ( .A(n516), .ZN(n489) );
  INV_X1 U404 ( .A(KEYINPUT54), .ZN(n435) );
  XOR2_X1 U405 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n353) );
  XNOR2_X1 U406 ( .A(G190GAT), .B(KEYINPUT77), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U408 ( .A(KEYINPUT78), .B(G106GAT), .Z(n355) );
  XNOR2_X1 U409 ( .A(G36GAT), .B(G99GAT), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n369) );
  XOR2_X1 U412 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n359) );
  XNOR2_X1 U413 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n358) );
  XOR2_X1 U414 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U415 ( .A(G85GAT), .B(G92GAT), .Z(n394) );
  XNOR2_X1 U416 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n360), .B(KEYINPUT7), .ZN(n382) );
  XOR2_X1 U418 ( .A(n394), .B(n382), .Z(n362) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n367) );
  XOR2_X1 U422 ( .A(G43GAT), .B(G134GAT), .Z(n447) );
  XNOR2_X1 U423 ( .A(n447), .B(n365), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U425 ( .A(n369), .B(n368), .Z(n565) );
  INV_X1 U426 ( .A(n565), .ZN(n553) );
  XNOR2_X1 U427 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n405) );
  XOR2_X1 U428 ( .A(G22GAT), .B(G141GAT), .Z(n371) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(G197GAT), .ZN(n370) );
  XOR2_X1 U430 ( .A(n371), .B(n370), .Z(n386) );
  XOR2_X1 U431 ( .A(G36GAT), .B(G8GAT), .Z(n428) );
  XOR2_X1 U432 ( .A(G15GAT), .B(G113GAT), .Z(n373) );
  XNOR2_X1 U433 ( .A(G43GAT), .B(G50GAT), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U435 ( .A(n428), .B(n374), .Z(n376) );
  NAND2_X1 U436 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U438 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n378) );
  XNOR2_X1 U439 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U441 ( .A(n380), .B(n379), .Z(n384) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n575) );
  INV_X1 U445 ( .A(KEYINPUT41), .ZN(n403) );
  AND2_X1 U446 ( .A1(G230GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U448 ( .A(n389), .B(KEYINPUT31), .Z(n393) );
  XNOR2_X1 U449 ( .A(G99GAT), .B(G71GAT), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n390), .B(G120GAT), .ZN(n439) );
  XNOR2_X1 U451 ( .A(n439), .B(n391), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n396) );
  XOR2_X1 U454 ( .A(KEYINPUT76), .B(G64GAT), .Z(n426) );
  XNOR2_X1 U455 ( .A(n394), .B(n426), .ZN(n395) );
  XOR2_X1 U456 ( .A(n396), .B(n395), .Z(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n400) );
  XNOR2_X1 U458 ( .A(G176GAT), .B(KEYINPUT32), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n578) );
  XNOR2_X1 U461 ( .A(n403), .B(n578), .ZN(n548) );
  AND2_X1 U462 ( .A1(n575), .A2(n548), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n406) );
  NOR2_X1 U464 ( .A1(n553), .A2(n406), .ZN(n407) );
  NAND2_X1 U465 ( .A1(n482), .A2(n407), .ZN(n409) );
  XNOR2_X1 U466 ( .A(KEYINPUT45), .B(KEYINPUT110), .ZN(n411) );
  XOR2_X1 U467 ( .A(KEYINPUT36), .B(n553), .Z(n587) );
  NOR2_X1 U468 ( .A1(n482), .A2(n587), .ZN(n410) );
  XOR2_X1 U469 ( .A(n411), .B(n410), .Z(n412) );
  NOR2_X1 U470 ( .A1(n575), .A2(n412), .ZN(n414) );
  INV_X1 U471 ( .A(n578), .ZN(n413) );
  NAND2_X1 U472 ( .A1(n414), .A2(n413), .ZN(n415) );
  NAND2_X1 U473 ( .A1(n416), .A2(n415), .ZN(n418) );
  XOR2_X1 U474 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n420) );
  XNOR2_X1 U475 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U477 ( .A(n421), .B(G183GAT), .Z(n423) );
  XNOR2_X1 U478 ( .A(G169GAT), .B(G176GAT), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n451) );
  XOR2_X1 U480 ( .A(KEYINPUT80), .B(G92GAT), .Z(n425) );
  NAND2_X1 U481 ( .A1(G226GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U483 ( .A(n427), .B(n426), .Z(n430) );
  XNOR2_X1 U484 ( .A(n428), .B(G204GAT), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n451), .B(n431), .ZN(n433) );
  XOR2_X1 U487 ( .A(n433), .B(n432), .Z(n518) );
  NOR2_X1 U488 ( .A1(n527), .A2(n518), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n436) );
  NOR2_X1 U490 ( .A1(n489), .A2(n436), .ZN(n573) );
  NAND2_X1 U491 ( .A1(n462), .A2(n573), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n437), .B(KEYINPUT116), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n438), .B(KEYINPUT55), .ZN(n452) );
  XOR2_X1 U494 ( .A(KEYINPUT85), .B(n439), .Z(n441) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n445) );
  XNOR2_X1 U497 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U499 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n521) );
  INV_X1 U503 ( .A(n521), .ZN(n531) );
  NAND2_X1 U504 ( .A1(n452), .A2(n531), .ZN(n566) );
  NOR2_X1 U505 ( .A1(n482), .A2(n566), .ZN(n455) );
  NOR2_X1 U506 ( .A1(n553), .A2(n482), .ZN(n456) );
  XNOR2_X1 U507 ( .A(KEYINPUT16), .B(n456), .ZN(n471) );
  XOR2_X1 U508 ( .A(KEYINPUT28), .B(KEYINPUT65), .Z(n457) );
  XOR2_X1 U509 ( .A(n462), .B(n457), .Z(n498) );
  INV_X1 U510 ( .A(n498), .ZN(n530) );
  INV_X1 U511 ( .A(n518), .ZN(n492) );
  XNOR2_X1 U512 ( .A(KEYINPUT27), .B(n492), .ZN(n461) );
  NAND2_X1 U513 ( .A1(n489), .A2(n461), .ZN(n528) );
  XNOR2_X1 U514 ( .A(n521), .B(KEYINPUT87), .ZN(n458) );
  NOR2_X1 U515 ( .A1(n528), .A2(n458), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n530), .A2(n459), .ZN(n470) );
  NOR2_X1 U517 ( .A1(n462), .A2(n531), .ZN(n460) );
  XOR2_X1 U518 ( .A(n460), .B(KEYINPUT26), .Z(n546) );
  INV_X1 U519 ( .A(n546), .ZN(n572) );
  NAND2_X1 U520 ( .A1(n461), .A2(n572), .ZN(n467) );
  NAND2_X1 U521 ( .A1(n492), .A2(n531), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n464), .B(KEYINPUT25), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT94), .B(n465), .Z(n466) );
  NAND2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n468), .A2(n516), .ZN(n469) );
  NAND2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n481) );
  NAND2_X1 U528 ( .A1(n471), .A2(n481), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(KEYINPUT95), .ZN(n500) );
  INV_X1 U530 ( .A(n575), .ZN(n556) );
  NOR2_X1 U531 ( .A1(n556), .A2(n578), .ZN(n486) );
  NAND2_X1 U532 ( .A1(n500), .A2(n486), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT96), .B(n473), .Z(n479) );
  NAND2_X1 U534 ( .A1(n479), .A2(n489), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n479), .A2(n492), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U540 ( .A1(n531), .A2(n479), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NAND2_X1 U542 ( .A1(n498), .A2(n479), .ZN(n480) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(n480), .ZN(G1327GAT) );
  XOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT39), .Z(n491) );
  XOR2_X1 U545 ( .A(KEYINPUT98), .B(KEYINPUT38), .Z(n488) );
  NAND2_X1 U546 ( .A1(n482), .A2(n481), .ZN(n483) );
  NOR2_X1 U547 ( .A1(n587), .A2(n483), .ZN(n485) );
  XNOR2_X1 U548 ( .A(KEYINPUT97), .B(KEYINPUT37), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n485), .B(n484), .ZN(n515) );
  NAND2_X1 U550 ( .A1(n515), .A2(n486), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(n497) );
  NAND2_X1 U552 ( .A1(n497), .A2(n489), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n497), .A2(n492), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT99), .Z(n495) );
  NAND2_X1 U557 ( .A1(n497), .A2(n531), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U562 ( .A(n548), .ZN(n559) );
  NOR2_X1 U563 ( .A1(n575), .A2(n559), .ZN(n514) );
  NAND2_X1 U564 ( .A1(n514), .A2(n500), .ZN(n501) );
  XOR2_X1 U565 ( .A(KEYINPUT101), .B(n501), .Z(n510) );
  NOR2_X1 U566 ( .A1(n510), .A2(n516), .ZN(n505) );
  XOR2_X1 U567 ( .A(KEYINPUT100), .B(KEYINPUT102), .Z(n503) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U571 ( .A1(n518), .A2(n510), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT103), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n521), .A2(n510), .ZN(n508) );
  XOR2_X1 U575 ( .A(n508), .B(KEYINPUT104), .Z(n509) );
  XNOR2_X1 U576 ( .A(G71GAT), .B(n509), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n530), .A2(n510), .ZN(n512) );
  XNOR2_X1 U578 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U580 ( .A(G78GAT), .B(n513), .Z(G1335GAT) );
  NAND2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n516), .A2(n523), .ZN(n517) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n518), .A2(n523), .ZN(n519) );
  XOR2_X1 U585 ( .A(KEYINPUT106), .B(n519), .Z(n520) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n523), .ZN(n522) );
  XOR2_X1 U588 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  NOR2_X1 U589 ( .A1(n530), .A2(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT107), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(KEYINPUT111), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U596 ( .A1(n545), .A2(n532), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n575), .A2(n541), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n535) );
  NAND2_X1 U600 ( .A1(n541), .A2(n548), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT112), .Z(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n539) );
  NAND2_X1 U605 ( .A1(n541), .A2(n582), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U609 ( .A1(n541), .A2(n553), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n544), .Z(G1343GAT) );
  NOR2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n575), .A2(n554), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U616 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n582), .A2(n554), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n566), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(KEYINPUT117), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n566), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n561) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(KEYINPUT56), .B(n562), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT58), .B(n567), .Z(n568) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n568), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT122), .B(n571), .Z(n577) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT121), .B(n574), .Z(n586) );
  INV_X1 U641 ( .A(n586), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n585) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n589) );
  NOR2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U653 ( .A(n589), .B(n588), .Z(n590) );
  XNOR2_X1 U654 ( .A(KEYINPUT124), .B(n590), .ZN(G1355GAT) );
endmodule

