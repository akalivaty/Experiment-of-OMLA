//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G210), .A3(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n187), .B(KEYINPUT69), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(G210), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G101), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(new_n196), .A3(new_n194), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT2), .A2(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT2), .A3(G113), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n207));
  INV_X1    g021(.A(G113), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G116), .B(G119), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n210), .B1(new_n206), .B2(new_n209), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G134), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(G137), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT11), .A3(G134), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(G137), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n216), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n215), .A2(G137), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n217), .A2(G134), .ZN(new_n223));
  OAI21_X1  g037(.A(G131), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT1), .B1(new_n228), .B2(G146), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G128), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G143), .B(G146), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(KEYINPUT1), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n221), .A2(new_n224), .A3(KEYINPUT66), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n227), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n216), .A2(new_n218), .A3(new_n220), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n221), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n236), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  OR2_X1    g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n234), .A2(KEYINPUT65), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n236), .A2(KEYINPUT0), .A3(G128), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n245), .A2(new_n248), .A3(new_n251), .A4(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n213), .B1(new_n242), .B2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n229), .A2(G128), .B1(new_n232), .B2(new_n233), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n238), .A2(new_n232), .A3(new_n233), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n221), .B(new_n224), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n244), .A2(new_n221), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n213), .B(new_n257), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT28), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(KEYINPUT70), .B(KEYINPUT28), .C1(new_n254), .C2(new_n261), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n213), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n253), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n225), .A2(new_n226), .B1(new_n235), .B2(new_n239), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n241), .A2(new_n271), .B1(new_n272), .B2(new_n245), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n274));
  OAI211_X1 g088(.A(new_n269), .B(new_n270), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n200), .A3(new_n260), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n275), .A2(new_n200), .A3(KEYINPUT31), .A4(new_n260), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n201), .A2(new_n268), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT71), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n268), .A2(new_n201), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n278), .A2(new_n279), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n281), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n264), .A2(new_n200), .A3(new_n265), .A4(new_n267), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n275), .A2(new_n260), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT29), .B1(new_n292), .B2(new_n201), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n213), .B1(new_n253), .B2(new_n257), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT28), .B1(new_n261), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n267), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n200), .A2(KEYINPUT29), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G472), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n281), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT72), .A3(KEYINPUT32), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n290), .A2(new_n303), .A3(new_n306), .A4(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n310));
  INV_X1    g124(.A(G953), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(G221), .A3(G234), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT77), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT22), .B(G137), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n237), .A2(G119), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT73), .ZN(new_n318));
  INV_X1    g132(.A(G119), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G128), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n320), .B(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT24), .B(G110), .ZN(new_n324));
  INV_X1    g138(.A(G110), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n326));
  AND2_X1   g140(.A1(KEYINPUT23), .A2(G119), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n326), .A2(new_n317), .B1(new_n237), .B2(new_n327), .ZN(new_n328));
  OAI22_X1  g142(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n330), .A2(KEYINPUT16), .A3(G140), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G146), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(new_n331), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(G146), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n334), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(KEYINPUT75), .A3(G146), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n329), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G125), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n330), .A2(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT76), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n332), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n348), .A3(new_n231), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n328), .A2(new_n325), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n324), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n318), .B2(new_n322), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n338), .B(new_n349), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n316), .B1(new_n341), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n338), .A2(new_n335), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n336), .A2(new_n337), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n231), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n340), .A3(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n328), .A2(new_n325), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n361), .B(new_n362), .C1(new_n324), .C2(new_n323), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n354), .A3(new_n315), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n356), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n356), .A2(new_n364), .A3(KEYINPUT25), .A4(new_n357), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G217), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(G234), .B2(new_n357), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n356), .A2(new_n364), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n371), .A2(G902), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n310), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n371), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n367), .B2(new_n368), .ZN(new_n378));
  INV_X1    g192(.A(new_n375), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT78), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n309), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT9), .B(G234), .ZN(new_n383));
  OAI21_X1  g197(.A(G221), .B1(new_n383), .B2(G902), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G469), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(new_n357), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n229), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT79), .B(KEYINPUT1), .C1(new_n228), .C2(G146), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(G128), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n256), .B1(new_n392), .B2(new_n234), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G104), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(G107), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n395), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n394), .A2(G107), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n397), .A2(G104), .ZN(new_n403));
  OAI21_X1  g217(.A(G101), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n388), .B1(new_n393), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n391), .A2(G128), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT79), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n234), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n239), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n401), .A2(new_n404), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(KEYINPUT80), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT10), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n240), .A3(KEYINPUT10), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n395), .A2(new_n398), .A3(new_n400), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(G101), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n417), .A2(G101), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n416), .B1(new_n422), .B2(new_n259), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n415), .A2(new_n424), .A3(KEYINPUT83), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT83), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT10), .B1(new_n406), .B2(new_n412), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(new_n423), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n428), .A3(new_n245), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n423), .B1(new_n413), .B2(new_n414), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n258), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G140), .ZN(new_n433));
  INV_X1    g247(.A(G227), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(G953), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n433), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n405), .A2(new_n235), .A3(new_n239), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n393), .A2(new_n388), .A3(new_n405), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT80), .B1(new_n410), .B2(new_n411), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT12), .A3(new_n245), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT81), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n441), .A2(KEYINPUT81), .A3(KEYINPUT12), .A4(new_n245), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n245), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n436), .B1(new_n430), .B2(new_n258), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n437), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n387), .B1(new_n452), .B2(new_n386), .ZN(new_n453));
  INV_X1    g267(.A(new_n436), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n431), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT82), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n450), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n458), .A3(new_n429), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT12), .B1(new_n441), .B2(new_n245), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(new_n443), .B2(new_n442), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n461), .A2(new_n445), .B1(new_n258), .B2(new_n430), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n459), .B(G469), .C1(new_n462), .C2(new_n454), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n385), .B1(new_n453), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n240), .A2(new_n330), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n248), .A2(new_n251), .A3(G125), .A4(new_n252), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT85), .B(G224), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(G953), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n469), .B(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n210), .A2(KEYINPUT5), .ZN(new_n474));
  INV_X1    g288(.A(G116), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n475), .A2(KEYINPUT5), .A3(G119), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n208), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n411), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(G110), .B(G122), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n479), .B(new_n480), .C1(new_n422), .C2(new_n213), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT6), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n479), .B1(new_n422), .B2(new_n213), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n480), .A2(KEYINPUT84), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(KEYINPUT6), .A3(new_n484), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n472), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n480), .B(KEYINPUT8), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n478), .A2(new_n473), .B1(new_n401), .B2(new_n404), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n479), .B2(KEYINPUT86), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n411), .A2(new_n493), .A3(new_n473), .A4(new_n478), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n471), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT7), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n469), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n467), .A2(new_n468), .A3(new_n497), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n481), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n357), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n466), .B1(new_n488), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n501), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n492), .A2(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n489), .ZN(new_n506));
  AOI21_X1  g320(.A(G902), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n469), .B(new_n496), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n481), .A2(KEYINPUT6), .B1(new_n483), .B2(new_n484), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n483), .A2(KEYINPUT6), .A3(new_n484), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n511), .A3(new_n465), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n503), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G214), .B1(G237), .B2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n345), .A2(G146), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n349), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G237), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n311), .A3(G214), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n228), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n522));
  NAND2_X1  g336(.A1(KEYINPUT18), .A2(G131), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n522), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT18), .A3(G131), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n518), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G113), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n394), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n525), .A2(G131), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n521), .A2(new_n219), .A3(new_n522), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n525), .A2(KEYINPUT17), .A3(G131), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n527), .B(new_n529), .C1(new_n535), .C2(new_n361), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n526), .A2(new_n524), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n530), .A2(new_n532), .B1(G146), .B2(new_n333), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n345), .A2(KEYINPUT19), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n346), .A2(new_n348), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n231), .B(new_n539), .C1(new_n540), .C2(KEYINPUT19), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n518), .A2(new_n537), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n536), .B1(new_n542), .B2(new_n529), .ZN(new_n543));
  NOR2_X1   g357(.A1(G475), .A2(G902), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT20), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT20), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n543), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n339), .A2(new_n533), .A3(new_n340), .A4(new_n534), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n529), .B1(new_n550), .B2(new_n527), .ZN(new_n551));
  INV_X1    g365(.A(new_n536), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n357), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G475), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n228), .A2(G128), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n237), .A2(G143), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT90), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT90), .ZN(new_n560));
  AOI21_X1  g374(.A(G134), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n560), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n562), .A2(new_n215), .A3(new_n558), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT91), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G122), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n565), .A2(KEYINPUT87), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(KEYINPUT87), .ZN(new_n567));
  OAI21_X1  g381(.A(G116), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT88), .B1(new_n565), .B2(G116), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT88), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n475), .A3(G122), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT14), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n569), .A2(new_n571), .A3(KEYINPUT92), .A4(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n569), .A2(new_n571), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n568), .B(new_n573), .C1(new_n574), .C2(new_n572), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT92), .B1(new_n574), .B2(new_n572), .ZN(new_n576));
  OAI21_X1  g390(.A(G107), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n569), .A2(new_n571), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n568), .A2(new_n397), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n559), .A2(G134), .A3(new_n560), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n215), .B1(new_n562), .B2(new_n558), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT91), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n564), .A2(new_n577), .A3(new_n580), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n556), .A2(KEYINPUT89), .A3(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n587), .B(new_n557), .C1(new_n586), .C2(new_n556), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT89), .B1(new_n556), .B2(new_n586), .ZN(new_n589));
  OAI21_X1  g403(.A(G134), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n568), .A2(new_n578), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n397), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n590), .B(new_n582), .C1(new_n592), .C2(new_n579), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n383), .A2(new_n370), .A3(G953), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n585), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n585), .B2(new_n593), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n357), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(G478), .ZN(new_n599));
  NOR2_X1   g413(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n585), .A2(new_n593), .ZN(new_n605));
  INV_X1    g419(.A(new_n594), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n595), .ZN(new_n608));
  INV_X1    g422(.A(new_n603), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n357), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n555), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(G234), .A2(G237), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(G952), .A3(new_n311), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT21), .B(G898), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(G902), .A3(G953), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT94), .Z(new_n619));
  AND2_X1   g433(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n464), .A2(new_n516), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n382), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n280), .B2(G902), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(KEYINPUT95), .B(G472), .C1(new_n280), .C2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n283), .A2(new_n288), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n455), .B1(new_n461), .B2(new_n445), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n454), .B1(new_n429), .B2(new_n431), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n386), .B(new_n357), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n387), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n463), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n381), .A2(new_n637), .A3(new_n384), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n624), .B1(new_n632), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n630), .B1(new_n627), .B2(new_n628), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(new_n464), .A3(KEYINPUT96), .A4(new_n381), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n503), .A2(KEYINPUT97), .A3(new_n512), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n507), .A2(new_n511), .A3(new_n644), .A4(new_n465), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n643), .A2(new_n514), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n619), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n608), .A2(KEYINPUT33), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n607), .A2(new_n649), .A3(new_n595), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n648), .A2(G478), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n599), .A2(new_n357), .ZN(new_n652));
  AOI21_X1  g466(.A(G902), .B1(new_n607), .B2(new_n595), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n652), .B1(new_n653), .B2(new_n599), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n555), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n642), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT98), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  NAND3_X1  g474(.A1(new_n546), .A2(KEYINPUT99), .A3(new_n548), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n547), .B1(new_n543), .B2(new_n544), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n662), .A2(new_n663), .B1(new_n553), .B2(G475), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n611), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n646), .A2(new_n619), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n642), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT100), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT35), .B(G107), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  NAND2_X1  g485(.A1(new_n363), .A2(new_n354), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n316), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n374), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n372), .A2(new_n675), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n629), .A2(new_n631), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n621), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  OAI21_X1  g494(.A(new_n614), .B1(new_n617), .B2(G900), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n665), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n643), .A2(new_n514), .A3(new_n645), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n309), .A2(new_n464), .A3(new_n676), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XOR2_X1   g500(.A(new_n513), .B(KEYINPUT38), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n555), .A2(new_n611), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n676), .A2(new_n688), .A3(new_n515), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n637), .A2(new_n384), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n681), .B(KEYINPUT39), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT40), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n276), .ZN(new_n695));
  INV_X1    g509(.A(new_n295), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n200), .B1(new_n260), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n357), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G472), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n290), .A2(new_n306), .A3(new_n308), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n690), .A2(new_n694), .A3(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n691), .A2(KEYINPUT40), .A3(new_n693), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n228), .ZN(G45));
  NAND4_X1  g518(.A1(new_n555), .A2(new_n651), .A3(new_n654), .A4(new_n681), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n683), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n309), .A2(new_n464), .A3(new_n676), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  AOI22_X1  g522(.A1(new_n432), .A2(new_n436), .B1(new_n449), .B2(new_n450), .ZN(new_n709));
  OAI21_X1  g523(.A(G469), .B1(new_n709), .B2(G902), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n384), .A3(new_n635), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n710), .A2(KEYINPUT101), .A3(new_n384), .A4(new_n635), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n382), .A2(new_n715), .A3(new_n656), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT102), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n716), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n309), .A2(new_n713), .A3(new_n381), .A4(new_n714), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n666), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n475), .ZN(G18));
  AND4_X1   g536(.A1(new_n384), .A2(new_n646), .A3(new_n635), .A4(new_n710), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n309), .A2(new_n723), .A3(new_n620), .A4(new_n676), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NOR2_X1   g539(.A1(new_n647), .A2(new_n688), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n200), .B1(new_n296), .B2(new_n267), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n285), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n281), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n727), .B1(new_n278), .B2(new_n279), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT103), .B1(new_n732), .B2(new_n282), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n378), .A2(new_n379), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n625), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n726), .A2(new_n737), .A3(new_n713), .A4(new_n714), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  AOI21_X1  g553(.A(new_n730), .B1(new_n729), .B2(new_n281), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n732), .A2(KEYINPUT103), .A3(new_n282), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n625), .B(new_n676), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n705), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n723), .A3(new_n744), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n555), .A2(new_n651), .A3(new_n654), .A4(new_n681), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n734), .A3(new_n625), .A4(new_n676), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n646), .A2(new_n710), .A3(new_n384), .A4(new_n635), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT104), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  NAND4_X1  g565(.A1(new_n286), .A2(KEYINPUT105), .A3(KEYINPUT32), .A4(new_n281), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n289), .B1(new_n280), .B2(new_n282), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n303), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT105), .B1(new_n307), .B2(KEYINPUT32), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n735), .B(new_n746), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n503), .A2(new_n514), .A3(new_n512), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n637), .A2(new_n384), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT42), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n637), .A2(new_n384), .A3(new_n758), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n705), .A2(KEYINPUT42), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n309), .A3(new_n381), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n219), .ZN(G33));
  INV_X1    g579(.A(new_n682), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n761), .A2(new_n309), .A3(new_n381), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  INV_X1    g583(.A(new_n459), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n454), .B1(new_n449), .B2(new_n431), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n459), .B(KEYINPUT45), .C1(new_n462), .C2(new_n454), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(G469), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n636), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n775), .A2(new_n776), .B1(new_n386), .B2(new_n452), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n636), .ZN(new_n778));
  AOI211_X1 g592(.A(new_n385), .B(new_n693), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n651), .A2(new_n654), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n555), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT43), .B1(new_n780), .B2(new_n555), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n676), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n640), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(KEYINPUT44), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(KEYINPUT44), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n788), .A2(KEYINPUT106), .A3(new_n758), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT106), .B1(new_n788), .B2(new_n758), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n779), .B(new_n787), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  XOR2_X1   g605(.A(KEYINPUT107), .B(G137), .Z(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(G39));
  AOI21_X1  g607(.A(new_n385), .B1(new_n777), .B2(new_n778), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n309), .A2(new_n381), .A3(new_n705), .A4(new_n757), .ZN(new_n797));
  NOR2_X1   g611(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n796), .B(new_n797), .C1(new_n794), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n801));
  INV_X1    g615(.A(new_n711), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n758), .ZN(new_n803));
  INV_X1    g617(.A(new_n381), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n803), .A2(new_n700), .A3(new_n804), .A4(new_n614), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n549), .A3(new_n554), .A4(new_n780), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n783), .A2(new_n784), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n803), .A2(new_n614), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n806), .B1(new_n742), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n807), .A2(new_n736), .A3(new_n614), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n687), .A2(new_n514), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n802), .A3(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n812), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT50), .B1(new_n812), .B2(KEYINPUT114), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n813), .B2(new_n814), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n809), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n794), .A2(new_n798), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n794), .B2(new_n795), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n710), .A2(new_n635), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT109), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n824), .A2(new_n385), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n758), .B(new_n810), .C1(new_n822), .C2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n818), .B2(new_n819), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n801), .B1(new_n820), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n735), .B1(new_n754), .B2(new_n755), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n808), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n830), .A2(KEYINPUT48), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n311), .A2(G952), .ZN(new_n832));
  INV_X1    g646(.A(new_n655), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n832), .B1(new_n805), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n830), .A2(KEYINPUT48), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n810), .A2(new_n646), .A3(new_n802), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT117), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n831), .A2(new_n834), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n809), .A2(new_n801), .A3(new_n813), .A4(new_n814), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n838), .B1(new_n826), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n828), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n661), .A2(new_n664), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n604), .A2(new_n610), .A3(new_n681), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT110), .B1(new_n844), .B2(new_n758), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT110), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n842), .A2(new_n757), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n309), .A3(new_n464), .A4(new_n676), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n761), .A2(new_n743), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n767), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT111), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n849), .A2(new_n767), .A3(new_n853), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n621), .B1(new_n382), .B2(new_n677), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n612), .B1(new_n780), .B2(new_n555), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n857), .A2(new_n516), .A3(new_n619), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n639), .A2(new_n641), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n760), .A2(new_n763), .ZN(new_n862));
  INV_X1    g676(.A(new_n656), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n724), .B(new_n738), .C1(new_n720), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n721), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n855), .A2(new_n861), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n744), .B1(new_n743), .B2(new_n723), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT104), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n685), .B(new_n707), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n683), .A2(new_n688), .ZN(new_n873));
  INV_X1    g687(.A(new_n681), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n873), .A2(new_n676), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n700), .A3(new_n464), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n869), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT52), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n750), .A2(new_n685), .A3(new_n707), .A4(new_n876), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n869), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n867), .A2(new_n868), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n880), .B(KEYINPUT52), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT53), .B1(new_n866), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(KEYINPUT54), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n868), .B1(new_n866), .B2(new_n885), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n862), .A2(KEYINPUT53), .A3(new_n856), .A4(new_n859), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n854), .B2(new_n852), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  OR3_X1    g705(.A1(new_n864), .A2(new_n891), .A3(new_n721), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n864), .B2(new_n721), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n883), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n887), .B1(KEYINPUT54), .B2(new_n896), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n841), .A2(new_n897), .B1(G952), .B2(G953), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n781), .A2(new_n735), .A3(new_n384), .A4(new_n514), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n700), .A2(new_n687), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n824), .B(KEYINPUT49), .Z(new_n901));
  OAI21_X1  g715(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(G75));
  NAND3_X1  g716(.A1(new_n896), .A2(G210), .A3(G902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n509), .A2(new_n510), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n508), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  AOI22_X1  g723(.A1(new_n905), .A2(new_n908), .B1(new_n909), .B2(new_n903), .ZN(new_n910));
  AND4_X1   g724(.A1(KEYINPUT118), .A2(new_n903), .A3(new_n909), .A4(new_n908), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n311), .A2(G952), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(G51));
  XNOR2_X1  g727(.A(new_n387), .B(KEYINPUT57), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n888), .A2(new_n895), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n915), .B1(new_n888), .B2(new_n895), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT119), .ZN(new_n919));
  INV_X1    g733(.A(new_n709), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n921), .B(new_n914), .C1(new_n916), .C2(new_n917), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n896), .A2(G902), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n924), .A2(new_n774), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n912), .B1(new_n923), .B2(new_n925), .ZN(G54));
  INV_X1    g740(.A(new_n543), .ZN(new_n927));
  NAND2_X1  g741(.A1(KEYINPUT58), .A2(G475), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n912), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(G60));
  NAND2_X1  g747(.A1(new_n648), .A2(new_n650), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n652), .B(KEYINPUT59), .Z(new_n935));
  OAI211_X1 g749(.A(new_n934), .B(new_n935), .C1(new_n916), .C2(new_n917), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n930), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n934), .B1(new_n897), .B2(new_n935), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G63));
  XNOR2_X1  g753(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT60), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n888), .B2(new_n895), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n930), .B1(new_n943), .B2(new_n373), .ZN(new_n944));
  INV_X1    g758(.A(new_n942), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n896), .A2(new_n674), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(KEYINPUT120), .B(new_n940), .C1(new_n944), .C2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n946), .B(new_n930), .C1(new_n373), .C2(new_n943), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n940), .B1(new_n950), .B2(KEYINPUT120), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(G66));
  OAI21_X1  g766(.A(G953), .B1(new_n470), .B2(new_n615), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n860), .A2(new_n721), .A3(new_n864), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n906), .B1(G898), .B2(new_n311), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  OR2_X1    g771(.A1(new_n273), .A2(new_n274), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(new_n270), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n539), .B1(new_n540), .B2(KEYINPUT19), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n959), .B(new_n960), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n791), .A2(new_n799), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n703), .A2(new_n872), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n691), .A2(new_n693), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n382), .A2(new_n966), .A3(new_n758), .A4(new_n857), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n963), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n962), .B1(new_n968), .B2(G953), .ZN(new_n969));
  INV_X1    g783(.A(G900), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(G953), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT123), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n829), .A2(new_n873), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n779), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n767), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n872), .A2(new_n764), .A3(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n791), .A2(new_n799), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n972), .B1(new_n978), .B2(new_n311), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT124), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n961), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n969), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n434), .B2(new_n970), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT122), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT125), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n985), .A2(KEYINPUT125), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n983), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n983), .B2(new_n987), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n292), .A2(new_n201), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(new_n276), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n884), .A2(new_n886), .A3(new_n995), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n292), .B(KEYINPUT126), .Z(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(new_n201), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n912), .B1(new_n998), .B2(new_n993), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n201), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n978), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n997), .A2(new_n201), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n968), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n861), .A2(new_n865), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n996), .B(new_n999), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(G57));
endmodule


