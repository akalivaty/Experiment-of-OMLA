//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(G110), .B(G122), .Z(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT85), .ZN(new_n191));
  XNOR2_X1  g005(.A(G116), .B(G119), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(KEYINPUT70), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(KEYINPUT70), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT5), .ZN(new_n195));
  NOR3_X1   g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G116), .ZN(new_n198));
  OAI21_X1  g012(.A(G113), .B1(new_n198), .B2(KEYINPUT5), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n191), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT79), .B1(new_n201), .B2(G104), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(G104), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n207), .A2(G101), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n204), .B2(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n201), .A2(KEYINPUT3), .A3(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n201), .A2(G104), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT77), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n214), .B1(new_n210), .B2(new_n211), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT77), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(new_n213), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n208), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n222));
  OR3_X1    g036(.A1(new_n222), .A2(KEYINPUT2), .A3(G113), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(KEYINPUT2), .B2(G113), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n223), .A2(new_n224), .B1(KEYINPUT2), .B2(G113), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n192), .ZN(new_n226));
  INV_X1    g040(.A(new_n199), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n192), .B(KEYINPUT70), .ZN(new_n228));
  OAI211_X1 g042(.A(KEYINPUT85), .B(new_n227), .C1(new_n228), .C2(new_n195), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n200), .A2(new_n221), .A3(new_n226), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n212), .A2(new_n215), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT78), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n231), .A2(new_n235), .A3(new_n232), .A4(G101), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n231), .A2(G101), .ZN(new_n238));
  AND4_X1   g052(.A1(new_n219), .A2(new_n212), .A3(new_n213), .A4(new_n215), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n219), .B1(new_n218), .B2(new_n213), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT4), .B(new_n238), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n193), .A2(new_n194), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n226), .B1(new_n242), .B2(new_n225), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n237), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n190), .B1(new_n230), .B2(new_n244), .ZN(new_n245));
  OR2_X1    g059(.A1(new_n245), .A2(KEYINPUT86), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n230), .A2(new_n190), .A3(new_n244), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(KEYINPUT86), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n246), .A2(KEYINPUT6), .A3(new_n247), .A4(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n245), .A2(KEYINPUT87), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT87), .B1(new_n245), .B2(new_n250), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  OR2_X1    g068(.A1(KEYINPUT65), .A2(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT65), .A2(G146), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n258));
  OAI21_X1  g072(.A(G128), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n254), .A2(G146), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n256), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(G143), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G128), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT65), .A2(G146), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT65), .A2(G146), .ZN(new_n268));
  OAI21_X1  g082(.A(G143), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n270));
  NOR2_X1   g084(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n266), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n267), .A2(new_n268), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n261), .B1(new_n274), .B2(new_n254), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT68), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G146), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G143), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n269), .A2(G128), .A3(new_n279), .A4(new_n258), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n265), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G125), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT0), .B(G128), .Z(new_n284));
  NAND2_X1  g098(.A1(new_n264), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n269), .A2(KEYINPUT0), .A3(G128), .A4(new_n279), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G125), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G224), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(G953), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n291), .B(KEYINPUT88), .Z(new_n292));
  XNOR2_X1  g106(.A(new_n289), .B(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n249), .A2(new_n253), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT7), .B1(new_n290), .B2(G953), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n283), .A2(new_n288), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT89), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n289), .A2(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n207), .A2(G101), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n239), .B2(new_n240), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n200), .A2(new_n301), .A3(new_n226), .A4(new_n229), .ZN(new_n302));
  XOR2_X1   g116(.A(new_n189), .B(KEYINPUT8), .Z(new_n303));
  AOI21_X1  g117(.A(new_n199), .B1(KEYINPUT5), .B2(new_n192), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n225), .B2(new_n192), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n302), .B(new_n303), .C1(new_n301), .C2(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n299), .A2(new_n247), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n298), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n294), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G210), .B1(G237), .B2(G902), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n294), .A2(new_n310), .A3(new_n308), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n188), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G952), .ZN(new_n315));
  AOI211_X1 g129(.A(G953), .B(new_n315), .C1(G234), .C2(G237), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G902), .ZN(new_n318));
  INV_X1    g132(.A(G953), .ZN(new_n319));
  AOI211_X1 g133(.A(new_n318), .B(new_n319), .C1(G234), .C2(G237), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT21), .B(G898), .Z(new_n322));
  OAI21_X1  g136(.A(new_n317), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT100), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(G475), .A2(G902), .ZN(new_n326));
  AND2_X1   g140(.A1(G125), .A2(G140), .ZN(new_n327));
  NOR2_X1   g141(.A1(G125), .A2(G140), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT16), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n282), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(G146), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT75), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(new_n330), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n277), .ZN(new_n334));
  NOR2_X1   g148(.A1(G237), .A2(G953), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G214), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n254), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(G143), .A3(G214), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G131), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT17), .ZN(new_n341));
  INV_X1    g155(.A(G131), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n342), .A3(new_n338), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n339), .A2(KEYINPUT17), .A3(G131), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n332), .A2(new_n334), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G113), .B(G122), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT93), .B(G104), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT94), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n337), .A2(KEYINPUT90), .A3(new_n338), .ZN(new_n352));
  NAND2_X1  g166(.A1(KEYINPUT18), .A2(G131), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n337), .A2(KEYINPUT90), .A3(new_n338), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT91), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n327), .A2(new_n328), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n263), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n277), .B2(new_n359), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n357), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n358), .B1(new_n357), .B2(new_n361), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n346), .B(new_n351), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT95), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n357), .A2(new_n361), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT91), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n357), .A2(new_n358), .A3(new_n361), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT95), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n346), .A4(new_n351), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n340), .A2(new_n343), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n359), .A2(KEYINPUT92), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT19), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n331), .B(new_n373), .C1(new_n375), .C2(new_n274), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n349), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n372), .A2(KEYINPUT96), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT96), .B1(new_n372), .B2(new_n379), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT20), .B(new_n326), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n372), .A2(new_n379), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n326), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n349), .B1(new_n369), .B2(new_n346), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n365), .B2(new_n371), .ZN(new_n388));
  OAI21_X1  g202(.A(G475), .B1(new_n388), .B2(G902), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n382), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT97), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n382), .A2(new_n389), .A3(KEYINPUT97), .A4(new_n386), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G116), .B(G122), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n201), .ZN(new_n396));
  XOR2_X1   g210(.A(G128), .B(G143), .Z(new_n397));
  OR2_X1    g211(.A1(new_n397), .A2(G134), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT13), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n254), .A3(G128), .ZN(new_n400));
  OAI211_X1 g214(.A(G134), .B(new_n400), .C1(new_n397), .C2(new_n399), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT98), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n397), .A2(G134), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G116), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT14), .A3(G122), .ZN(new_n408));
  INV_X1    g222(.A(new_n395), .ZN(new_n409));
  OAI211_X1 g223(.A(G107), .B(new_n408), .C1(new_n409), .C2(KEYINPUT14), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n406), .B(new_n410), .C1(G107), .C2(new_n409), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT9), .B(G234), .Z(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(G217), .A3(new_n319), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n412), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n318), .ZN(new_n416));
  INV_X1    g230(.A(G478), .ZN(new_n417));
  NOR2_X1   g231(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT99), .A2(KEYINPUT15), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n416), .B(new_n421), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n325), .A2(new_n394), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(G472), .A2(G902), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n265), .A2(new_n276), .A3(new_n280), .ZN(new_n425));
  INV_X1    g239(.A(G137), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G134), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT11), .ZN(new_n429));
  INV_X1    g243(.A(G134), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n426), .A2(KEYINPUT11), .A3(G134), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n428), .A2(new_n342), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n430), .A2(G137), .ZN(new_n434));
  OAI21_X1  g248(.A(G131), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n425), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n243), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n285), .A2(new_n286), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n431), .A2(new_n432), .ZN(new_n440));
  OAI21_X1  g254(.A(G131), .B1(new_n440), .B2(new_n427), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n433), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n335), .A2(G210), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(G101), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT72), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT72), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n451), .A3(new_n448), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n442), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT66), .B1(new_n454), .B2(new_n287), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT66), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n439), .A2(new_n456), .A3(new_n442), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n437), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND4_X1   g274(.A1(KEYINPUT71), .A2(new_n437), .A3(KEYINPUT30), .A4(new_n443), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n425), .A2(new_n436), .B1(new_n442), .B2(new_n439), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT71), .B1(new_n462), .B2(KEYINPUT30), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n243), .B(new_n460), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT31), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n453), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT28), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n444), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n458), .A2(new_n243), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n462), .A2(KEYINPUT28), .A3(new_n438), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n448), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n465), .B1(new_n453), .B2(new_n464), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n424), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT32), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT74), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n453), .A2(new_n464), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT31), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n466), .A3(new_n473), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(KEYINPUT32), .A3(new_n424), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n478), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n482), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n424), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n464), .A2(new_n444), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n472), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n468), .A2(new_n470), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n448), .A3(new_n469), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n462), .A2(new_n438), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n490), .A2(KEYINPUT29), .A3(new_n495), .A4(new_n448), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n488), .A2(KEYINPUT73), .A3(new_n489), .A4(new_n491), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n494), .A2(new_n318), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G472), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n486), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n197), .A2(G128), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n501), .A2(KEYINPUT23), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n266), .A2(G119), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(KEYINPUT23), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n501), .A2(new_n503), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  OAI22_X1  g322(.A1(new_n506), .A2(G110), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n331), .A3(new_n360), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT76), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n332), .A2(new_n334), .B1(G110), .B2(new_n506), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n508), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  XOR2_X1   g329(.A(KEYINPUT22), .B(G137), .Z(new_n516));
  AND3_X1   g330(.A1(new_n319), .A2(G221), .A3(G234), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n515), .B(new_n519), .ZN(new_n520));
  OR3_X1    g334(.A1(new_n520), .A2(KEYINPUT25), .A3(G902), .ZN(new_n521));
  INV_X1    g335(.A(G217), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(G234), .B2(new_n318), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT25), .B1(new_n520), .B2(G902), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OR3_X1    g339(.A1(new_n520), .A2(G902), .A3(new_n523), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G221), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n413), .B2(new_n318), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT84), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT80), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT1), .ZN(new_n534));
  OAI21_X1  g348(.A(G128), .B1(new_n261), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n257), .B2(new_n278), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n280), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n301), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n221), .A2(KEYINPUT80), .A3(new_n537), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n539), .A2(new_n540), .B1(new_n281), .B2(new_n301), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n532), .B1(new_n541), .B2(new_n454), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n301), .A2(new_n280), .A3(new_n276), .A4(new_n265), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n301), .A2(new_n538), .A3(new_n533), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT80), .B1(new_n221), .B2(new_n537), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT12), .A3(new_n442), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n542), .A2(new_n547), .A3(KEYINPUT83), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT83), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n532), .C1(new_n541), .C2(new_n454), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n539), .B2(new_n540), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n425), .A2(KEYINPUT10), .A3(new_n221), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n237), .A2(new_n439), .A3(new_n241), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT82), .B1(new_n557), .B2(new_n454), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT82), .ZN(new_n559));
  NOR4_X1   g373(.A1(new_n553), .A2(new_n556), .A3(new_n559), .A4(new_n442), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n548), .B(new_n550), .C1(new_n558), .C2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G140), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n319), .A2(G227), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n531), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n551), .B1(new_n544), .B2(new_n545), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n567), .A2(new_n454), .A3(new_n555), .A4(new_n554), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n559), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n557), .A2(KEYINPUT82), .A3(new_n454), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n539), .A2(new_n540), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n454), .B1(new_n571), .B2(new_n543), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n549), .B1(new_n572), .B2(KEYINPUT12), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n569), .A2(new_n570), .B1(new_n573), .B2(new_n542), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n574), .A2(KEYINPUT84), .A3(new_n564), .A4(new_n550), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n558), .A2(new_n560), .B1(new_n454), .B2(new_n557), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n565), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n566), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G469), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(new_n318), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n318), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n564), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n564), .B2(new_n561), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n581), .B1(new_n583), .B2(G469), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n530), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n423), .A2(new_n500), .A3(new_n528), .A4(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  AND2_X1   g401(.A1(new_n585), .A2(new_n528), .ZN(new_n588));
  INV_X1    g402(.A(G472), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n482), .B2(new_n318), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT101), .ZN(new_n591));
  INV_X1    g405(.A(new_n590), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n476), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n591), .B1(new_n593), .B2(KEYINPUT101), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n416), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(G478), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n415), .A2(KEYINPUT33), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n414), .B(KEYINPUT102), .Z(new_n600));
  NAND3_X1  g414(.A1(new_n412), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n412), .B2(new_n414), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(new_n412), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT33), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n598), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n597), .B1(new_n605), .B2(G478), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n394), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n325), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n595), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  OAI21_X1  g426(.A(new_n326), .B1(new_n380), .B2(new_n381), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n385), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n614), .A2(new_n389), .A3(new_n382), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n422), .A4(new_n324), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n614), .A2(new_n422), .A3(new_n389), .A4(new_n382), .ZN(new_n618));
  INV_X1    g432(.A(new_n324), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT104), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n595), .A2(new_n314), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NAND2_X1  g438(.A1(new_n580), .A2(new_n584), .ZN(new_n625));
  INV_X1    g439(.A(new_n530), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n515), .B(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n629), .B(new_n318), .C1(new_n522), .C2(G234), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n525), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n423), .A3(new_n594), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  OR2_X1    g450(.A1(new_n321), .A2(G900), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n317), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n618), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n314), .A2(new_n631), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n500), .A2(new_n585), .A3(new_n640), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  XNOR2_X1  g458(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n638), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n585), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT40), .Z(new_n648));
  AND3_X1   g462(.A1(new_n294), .A2(new_n310), .A3(new_n308), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n310), .B1(new_n294), .B2(new_n308), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT38), .ZN(new_n652));
  INV_X1    g466(.A(new_n394), .ZN(new_n653));
  INV_X1    g467(.A(new_n422), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n480), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n448), .B1(new_n495), .B2(new_n444), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n318), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(G472), .ZN(new_n659));
  AOI211_X1 g473(.A(new_n188), .B(new_n631), .C1(new_n486), .C2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n648), .A2(new_n655), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT106), .B(G143), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G45));
  NAND3_X1  g477(.A1(new_n394), .A2(new_n607), .A3(new_n638), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(new_n500), .A3(new_n642), .A4(new_n585), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  AOI22_X1  g481(.A1(new_n484), .A2(new_n485), .B1(new_n498), .B2(G472), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n527), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n578), .A2(new_n318), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G469), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n671), .A2(new_n626), .A3(new_n580), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n669), .A2(new_n609), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT41), .B(G113), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G15));
  NAND4_X1  g489(.A1(new_n671), .A2(new_n626), .A3(new_n580), .A4(new_n314), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n669), .A2(new_n677), .A3(new_n621), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  NAND4_X1  g493(.A1(new_n672), .A2(new_n423), .A3(new_n500), .A4(new_n631), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G119), .ZN(G21));
  AND3_X1   g495(.A1(new_n394), .A2(new_n314), .A3(new_n422), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n448), .B1(new_n490), .B2(new_n495), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n656), .B2(new_n465), .ZN(new_n684));
  AOI211_X1 g498(.A(G472), .B(G902), .C1(new_n684), .C2(new_n481), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n527), .A2(new_n685), .A3(new_n590), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n672), .A2(new_n682), .A3(new_n324), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G122), .ZN(G24));
  NOR3_X1   g502(.A1(new_n632), .A2(new_n590), .A3(new_n685), .ZN(new_n689));
  AND4_X1   g503(.A1(KEYINPUT107), .A2(new_n394), .A3(new_n607), .A4(new_n638), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n606), .B1(new_n392), .B2(new_n393), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT107), .B1(new_n691), .B2(new_n638), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n677), .B(new_n689), .C1(new_n690), .C2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  NAND2_X1  g508(.A1(new_n312), .A2(new_n313), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT108), .B1(new_n695), .B2(new_n188), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n651), .A2(new_n697), .A3(new_n187), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n585), .B(new_n700), .C1(new_n690), .C2(new_n692), .ZN(new_n701));
  INV_X1    g515(.A(new_n669), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT109), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT107), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n664), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n691), .A2(KEYINPUT107), .A3(new_n638), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n627), .A2(new_n699), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n669), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n703), .A2(new_n704), .A3(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n499), .A2(new_n483), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n527), .B1(new_n713), .B2(new_n478), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n708), .A3(new_n709), .A4(KEYINPUT42), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  OAI21_X1  g531(.A(KEYINPUT110), .B1(new_n618), .B2(new_n639), .ZN(new_n718));
  OR3_X1    g532(.A1(new_n618), .A2(KEYINPUT110), .A3(new_n639), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n709), .A2(new_n669), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G134), .ZN(G36));
  NAND2_X1  g535(.A1(new_n653), .A2(new_n607), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n653), .A2(KEYINPUT43), .A3(new_n607), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n594), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n726), .A2(new_n727), .A3(new_n631), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n727), .B1(new_n726), .B2(new_n631), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n583), .A2(KEYINPUT45), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n583), .A2(KEYINPUT45), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n732), .A2(new_n733), .A3(new_n579), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n731), .B1(new_n734), .B2(new_n581), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT111), .ZN(new_n736));
  OR3_X1    g550(.A1(new_n734), .A2(new_n731), .A3(new_n581), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(new_n731), .C1(new_n734), .C2(new_n581), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n580), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n626), .A3(new_n646), .A4(new_n700), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n730), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n426), .ZN(G39));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n626), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n699), .A2(new_n664), .ZN(new_n749));
  AOI22_X1  g563(.A1(new_n740), .A2(new_n626), .B1(new_n745), .B2(new_n746), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n748), .B(new_n749), .C1(new_n747), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n500), .A2(new_n528), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT113), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n747), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n740), .B2(new_n626), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n745), .A2(new_n746), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n744), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n756), .B1(new_n758), .B2(new_n755), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n752), .A4(new_n749), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G140), .ZN(G42));
  INV_X1    g577(.A(new_n722), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n671), .A2(new_n580), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n764), .B(new_n652), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n486), .A2(new_n659), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n527), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n768), .A2(new_n626), .A3(new_n187), .A4(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n693), .A2(new_n643), .A3(new_n666), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n625), .A2(new_n626), .A3(new_n632), .A4(new_n638), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT114), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n585), .A2(new_n776), .A3(new_n632), .A4(new_n638), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n769), .A2(new_n775), .A3(new_n682), .A4(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT115), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n696), .A2(new_n615), .A3(new_n698), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n422), .A2(new_n639), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n633), .A2(new_n782), .A3(new_n500), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n689), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n720), .B(new_n784), .C1(new_n701), .C2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n678), .A2(new_n673), .A3(new_n680), .A4(new_n687), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n608), .B1(new_n394), .B2(new_n654), .ZN(new_n788));
  INV_X1    g602(.A(new_n325), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n588), .A2(new_n788), .A3(new_n789), .A4(new_n594), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n634), .A3(new_n586), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n786), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT115), .B(KEYINPUT52), .C1(new_n773), .C2(new_n778), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n781), .A2(new_n716), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT52), .B1(new_n773), .B2(new_n778), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n676), .B1(new_n706), .B2(new_n707), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n627), .A2(new_n668), .A3(new_n641), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n798), .A2(new_n689), .B1(new_n799), .B2(new_n640), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n775), .A2(new_n769), .A3(new_n682), .A4(new_n777), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n780), .A3(new_n666), .A4(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(KEYINPUT53), .A3(new_n716), .A4(new_n792), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n772), .B1(new_n796), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n806));
  NAND2_X1  g620(.A1(new_n794), .A2(KEYINPUT53), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n803), .A2(new_n795), .A3(new_n716), .A4(new_n792), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n724), .A2(new_n725), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n316), .A3(new_n686), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n766), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n626), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n700), .B(new_n813), .C1(new_n759), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n672), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n317), .A3(new_n699), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n770), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n394), .A3(new_n607), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n652), .A2(new_n188), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n812), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n822), .A2(KEYINPUT50), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(KEYINPUT50), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n818), .A2(new_n811), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n689), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT117), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n816), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n816), .A2(new_n825), .A3(KEYINPUT51), .A4(new_n828), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n826), .A2(new_n714), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT48), .Z(new_n834));
  OAI211_X1 g648(.A(G952), .B(new_n319), .C1(new_n819), .C2(new_n608), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n831), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n812), .A2(new_n676), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n810), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(G952), .A2(G953), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n771), .B1(new_n839), .B2(new_n840), .ZN(G75));
  NOR2_X1   g655(.A1(new_n319), .A2(G952), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n807), .A2(G210), .A3(G902), .A4(new_n808), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n249), .A2(new_n253), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT118), .Z(new_n848));
  XOR2_X1   g662(.A(new_n293), .B(KEYINPUT55), .Z(new_n849));
  XOR2_X1   g663(.A(new_n848), .B(new_n849), .Z(new_n850));
  AOI21_X1  g664(.A(KEYINPUT119), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n852));
  INV_X1    g666(.A(new_n850), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n852), .B(new_n853), .C1(new_n844), .C2(new_n845), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n843), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n807), .A2(G902), .A3(new_n808), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT120), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n807), .A2(new_n858), .A3(G902), .A4(new_n808), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n311), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n860), .A2(KEYINPUT121), .A3(new_n861), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n855), .B1(new_n864), .B2(new_n865), .ZN(G51));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n807), .A2(new_n808), .ZN(new_n868));
  INV_X1    g682(.A(new_n806), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n809), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n807), .A2(KEYINPUT122), .A3(new_n806), .A4(new_n808), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n581), .B(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n578), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n857), .A2(new_n859), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n734), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n842), .B1(new_n876), .B2(new_n878), .ZN(G54));
  INV_X1    g693(.A(new_n380), .ZN(new_n880));
  INV_X1    g694(.A(new_n381), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(KEYINPUT58), .A2(G475), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n877), .A2(KEYINPUT123), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n857), .A2(new_n859), .A3(new_n883), .ZN(new_n886));
  INV_X1    g700(.A(new_n882), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n842), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(G60));
  NAND2_X1  g704(.A1(new_n598), .A2(new_n604), .ZN(new_n891));
  NAND2_X1  g705(.A1(G478), .A2(G902), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT59), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n873), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n893), .B1(new_n805), .B2(new_n809), .ZN(new_n895));
  INV_X1    g709(.A(new_n891), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n842), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n894), .A2(new_n897), .ZN(G63));
  INV_X1    g712(.A(new_n868), .ZN(new_n899));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT60), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n842), .B1(new_n903), .B2(new_n520), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n629), .A3(new_n902), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT61), .B1(new_n905), .B2(KEYINPUT124), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n904), .B(new_n905), .C1(KEYINPUT124), .C2(KEYINPUT61), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(G66));
  INV_X1    g724(.A(new_n322), .ZN(new_n911));
  OAI21_X1  g725(.A(G953), .B1(new_n911), .B2(new_n290), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n787), .A2(new_n791), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(G953), .ZN(new_n914));
  INV_X1    g728(.A(new_n848), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(G898), .B2(new_n319), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n914), .B(new_n916), .ZN(G69));
  OAI21_X1  g731(.A(new_n460), .B1(new_n461), .B2(new_n463), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(new_n375), .Z(new_n919));
  AOI21_X1  g733(.A(new_n773), .B1(new_n712), .B2(new_n715), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n714), .A2(new_n682), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n921), .A2(new_n740), .A3(new_n626), .A4(new_n646), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n922), .B(new_n720), .C1(new_n730), .C2(new_n741), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n762), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n919), .B1(new_n925), .B2(new_n319), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(G227), .B2(new_n319), .ZN(new_n927));
  INV_X1    g741(.A(new_n919), .ZN(new_n928));
  OAI21_X1  g742(.A(G900), .B1(new_n928), .B2(G227), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(G953), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n661), .A2(new_n666), .A3(new_n800), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT62), .Z(new_n932));
  INV_X1    g746(.A(new_n647), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n933), .A2(new_n669), .A3(new_n700), .A4(new_n788), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n730), .B2(new_n741), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT125), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n934), .C1(new_n730), .C2(new_n741), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n762), .A2(new_n932), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n319), .A3(new_n919), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n927), .A2(new_n930), .A3(new_n941), .ZN(G72));
  NAND4_X1  g756(.A1(new_n762), .A2(new_n932), .A3(new_n939), .A4(new_n913), .ZN(new_n943));
  XNOR2_X1  g757(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n589), .A2(new_n318), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(new_n448), .A3(new_n487), .ZN(new_n948));
  AOI22_X1  g762(.A1(new_n796), .A2(new_n804), .B1(new_n488), .B2(new_n480), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n842), .B1(new_n949), .B2(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n762), .A2(new_n924), .A3(new_n913), .A4(new_n920), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(new_n946), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n952), .B2(new_n946), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n448), .ZN(new_n956));
  INV_X1    g770(.A(new_n487), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(G57));
endmodule


