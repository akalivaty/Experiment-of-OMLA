//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  AOI211_X1 g007(.A(new_n202), .B(new_n204), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n210));
  NOR2_X1   g009(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT75), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(KEYINPUT75), .B(new_n208), .C1(new_n210), .C2(new_n211), .ZN(new_n215));
  INV_X1    g014(.A(new_n202), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT73), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n203), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT73), .B1(new_n204), .B2(new_n202), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n214), .A2(new_n215), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(new_n205), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n209), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n225));
  INV_X1    g024(.A(G113gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(KEYINPUT67), .A3(G120gat), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n224), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n226), .A2(G120gat), .ZN(new_n229));
  INV_X1    g028(.A(G120gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(G113gat), .ZN(new_n231));
  OR3_X1    g030(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT67), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n225), .B1(new_n229), .B2(new_n231), .ZN(new_n233));
  INV_X1    g032(.A(new_n224), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n228), .A2(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n223), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT5), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n238), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(new_n223), .B2(new_n235), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT79), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT74), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n206), .ZN(new_n245));
  NAND2_X1  g044(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n221), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n218), .B(new_n219), .C1(new_n247), .C2(KEYINPUT75), .ZN(new_n248));
  INV_X1    g047(.A(new_n215), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n222), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n209), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n250), .A2(new_n241), .A3(new_n235), .A4(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT80), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n240), .B1(new_n243), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n251), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n235), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT77), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n223), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n223), .B2(new_n258), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT78), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT78), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n256), .B(new_n263), .C1(new_n259), .C2(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n239), .B1(new_n254), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT82), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT82), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n223), .A2(new_n269), .A3(new_n241), .A4(new_n235), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n242), .A2(KEYINPUT81), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n268), .B(new_n270), .C1(KEYINPUT81), .C2(new_n242), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n262), .B2(new_n264), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n240), .A2(KEYINPUT5), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT83), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n275), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n279), .A2(new_n265), .A3(KEYINPUT83), .A4(new_n277), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n267), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT87), .ZN(new_n283));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT0), .ZN(new_n285));
  XNOR2_X1  g084(.A(G57gat), .B(G85gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n282), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT83), .ZN(new_n290));
  INV_X1    g089(.A(new_n264), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n250), .A2(new_n251), .A3(new_n258), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT77), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n223), .A2(new_n257), .A3(new_n258), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n263), .B1(new_n295), .B2(new_n256), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n273), .B(new_n274), .C1(new_n291), .C2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n277), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n266), .B1(new_n299), .B2(new_n280), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT6), .B1(new_n300), .B2(new_n287), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT87), .B1(new_n300), .B2(new_n287), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n289), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G8gat), .B(G36gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(G64gat), .B(G92gat), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n304), .B(new_n305), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT26), .ZN(new_n309));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n310), .A2(KEYINPUT66), .A3(new_n309), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT66), .B1(new_n310), .B2(new_n309), .ZN(new_n312));
  OAI221_X1 g111(.A(new_n308), .B1(new_n309), .B2(new_n310), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G183gat), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n314), .A2(KEYINPUT27), .ZN(new_n315));
  INV_X1    g114(.A(G190gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(KEYINPUT27), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n318), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n313), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(G183gat), .A3(G190gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n314), .A2(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n316), .A2(G183gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n327), .B2(KEYINPUT24), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n310), .A2(KEYINPUT23), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n329), .A2(new_n308), .A3(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n328), .A2(new_n332), .A3(KEYINPUT65), .A4(KEYINPUT25), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n334));
  XNOR2_X1  g133(.A(G183gat), .B(G190gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n323), .B1(new_n335), .B2(new_n322), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n329), .A2(KEYINPUT25), .A3(new_n331), .A4(new_n308), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n329), .A2(new_n308), .A3(new_n331), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n336), .B2(KEYINPUT64), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT64), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n342), .B(new_n323), .C1(new_n335), .C2(new_n322), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT25), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n321), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G197gat), .B(G204gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT70), .B(G211gat), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n350), .A2(G218gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n349), .B1(new_n351), .B2(KEYINPUT22), .ZN(new_n352));
  XNOR2_X1  g151(.A(G211gat), .B(G218gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n352), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n345), .A2(new_n356), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n348), .B(new_n355), .C1(new_n357), .C2(new_n347), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n352), .B(new_n353), .ZN(new_n359));
  INV_X1    g158(.A(new_n348), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT71), .B(KEYINPUT29), .Z(new_n361));
  AOI21_X1  g160(.A(new_n347), .B1(new_n345), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n307), .B1(new_n364), .B2(KEYINPUT37), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(KEYINPUT37), .B2(new_n364), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT38), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n358), .A2(new_n363), .A3(new_n306), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n348), .B1(new_n357), .B2(new_n347), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT37), .B1(new_n370), .B2(new_n355), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n360), .A2(new_n362), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(new_n359), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n367), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n369), .B1(new_n374), .B2(new_n365), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n282), .A2(KEYINPUT6), .A3(new_n288), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n303), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G228gat), .ZN(new_n379));
  INV_X1    g178(.A(G233gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT3), .B1(new_n355), .B2(new_n356), .ZN(new_n382));
  INV_X1    g181(.A(new_n361), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n383), .B1(new_n293), .B2(new_n294), .ZN(new_n384));
  OAI221_X1 g183(.A(new_n381), .B1(new_n382), .B2(new_n223), .C1(new_n384), .C2(new_n355), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n361), .B1(new_n259), .B2(new_n260), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n258), .B1(new_n359), .B2(new_n383), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n386), .A2(new_n359), .B1(new_n387), .B2(new_n255), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n388), .A2(KEYINPUT84), .A3(new_n381), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n390));
  INV_X1    g189(.A(new_n258), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n355), .B2(new_n361), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n384), .A2(new_n355), .B1(new_n392), .B2(new_n223), .ZN(new_n393));
  INV_X1    g192(.A(new_n381), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n385), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT85), .B1(new_n396), .B2(G22gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(G78gat), .B(G106gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT31), .B(G50gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n396), .A2(G22gat), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT84), .B1(new_n388), .B2(new_n381), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n393), .A2(new_n390), .A3(new_n394), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n403), .B1(new_n406), .B2(new_n385), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n397), .A2(new_n401), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n396), .A2(G22gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n403), .A3(new_n385), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT85), .A4(new_n400), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n289), .A2(new_n302), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n237), .A2(new_n238), .ZN(new_n414));
  OAI211_X1 g213(.A(KEYINPUT39), .B(new_n414), .C1(new_n276), .C2(new_n238), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT86), .B(KEYINPUT39), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n297), .A2(new_n240), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n287), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT40), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n415), .A2(KEYINPUT40), .A3(new_n287), .A4(new_n417), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n364), .A2(new_n307), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n369), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT72), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n369), .A2(new_n425), .A3(new_n423), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n369), .B2(new_n423), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n422), .B(new_n424), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n420), .A2(new_n421), .A3(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n378), .B(new_n412), .C1(new_n413), .C2(new_n429), .ZN(new_n430));
  XOR2_X1   g229(.A(G15gat), .B(G43gat), .Z(new_n431));
  XNOR2_X1  g230(.A(G71gat), .B(G99gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n336), .A2(KEYINPUT64), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n343), .A3(new_n332), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT25), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n436), .A2(new_n437), .B1(new_n333), .B2(new_n338), .ZN(new_n438));
  INV_X1    g237(.A(new_n321), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n236), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n235), .B(new_n321), .C1(new_n339), .C2(new_n344), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n433), .B1(new_n442), .B2(KEYINPUT33), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT32), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(new_n441), .ZN(new_n447));
  INV_X1    g246(.A(new_n434), .ZN(new_n448));
  AOI221_X4 g247(.A(new_n444), .B1(KEYINPUT33), .B2(new_n433), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n440), .A2(new_n434), .A3(new_n441), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT34), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT34), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n440), .A2(new_n453), .A3(new_n441), .A4(new_n434), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n452), .B1(new_n451), .B2(new_n454), .ZN(new_n456));
  OAI22_X1  g255(.A1(new_n446), .A2(new_n449), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT69), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n459));
  OAI221_X1 g258(.A(new_n459), .B1(new_n455), .B2(new_n456), .C1(new_n446), .C2(new_n449), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(new_n454), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n446), .A2(new_n449), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT36), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n461), .B1(new_n446), .B2(new_n449), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n466), .A2(KEYINPUT36), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n287), .B(new_n267), .C1(new_n278), .C2(new_n281), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n300), .A2(new_n287), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n377), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n428), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n408), .A2(new_n411), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n463), .B1(new_n408), .B2(new_n411), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(new_n474), .A3(new_n473), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n303), .A2(new_n377), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n428), .A2(new_n466), .A3(KEYINPUT35), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n412), .A3(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n430), .A2(new_n477), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT97), .ZN(new_n485));
  NAND2_X1  g284(.A1(G229gat), .A2(G233gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n486), .B(KEYINPUT13), .Z(new_n487));
  INV_X1    g286(.A(G1gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT16), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G22gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT93), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n403), .A2(G15gat), .ZN(new_n492));
  INV_X1    g291(.A(G15gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G22gat), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT93), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n489), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n492), .A2(new_n494), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n490), .A2(KEYINPUT93), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n488), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT94), .B(G8gat), .Z(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT95), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n496), .A2(new_n501), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G8gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n496), .A2(new_n501), .A3(new_n507), .A4(new_n502), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT90), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OR3_X1    g313(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G43gat), .B(G50gat), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n517), .A2(KEYINPUT15), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(KEYINPUT15), .ZN(new_n519));
  NAND2_X1  g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n516), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n514), .A2(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n512), .A2(KEYINPUT91), .A3(new_n513), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n517), .A2(new_n515), .A3(KEYINPUT15), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n509), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n509), .A2(new_n527), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n487), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n506), .A2(new_n508), .ZN(new_n531));
  OAI211_X1 g330(.A(KEYINPUT17), .B(new_n521), .C1(new_n525), .C2(new_n526), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT92), .B(KEYINPUT17), .ZN(new_n533));
  INV_X1    g332(.A(new_n521), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n526), .B1(new_n523), .B2(new_n524), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n531), .A2(new_n504), .A3(new_n532), .A4(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT96), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n509), .A2(new_n527), .ZN(new_n539));
  INV_X1    g338(.A(new_n486), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n530), .A2(new_n543), .ZN(new_n544));
  AOI211_X1 g343(.A(new_n541), .B(new_n540), .C1(new_n509), .C2(new_n527), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n538), .B1(new_n545), .B2(new_n537), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n485), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n537), .A2(new_n539), .A3(new_n486), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n541), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n539), .A2(new_n542), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n536), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n551), .A2(new_n509), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT96), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n553), .A2(KEYINPUT97), .A3(new_n530), .A4(new_n543), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G169gat), .B(G197gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT12), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT89), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n549), .B(new_n564), .ZN(new_n565));
  AND4_X1   g364(.A1(new_n553), .A2(new_n530), .A3(new_n543), .A4(new_n561), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT99), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n555), .A2(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT99), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT8), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(KEYINPUT102), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT102), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n578), .A2(G99gat), .A3(G106gat), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n577), .A2(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n583), .B(new_n584), .C1(new_n580), .C2(new_n581), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n580), .B2(new_n581), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT7), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n582), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G99gat), .B(G106gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n582), .A2(new_n590), .A3(new_n585), .A4(new_n588), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n527), .A2(new_n595), .B1(KEYINPUT41), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n551), .B2(new_n595), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n602), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT104), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n600), .B(new_n601), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n607), .B(new_n608), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G57gat), .B(G64gat), .Z(new_n614));
  INV_X1    g413(.A(KEYINPUT9), .ZN(new_n615));
  INV_X1    g414(.A(G71gat), .ZN(new_n616));
  INV_X1    g415(.A(G78gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G71gat), .B(G78gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n614), .A2(new_n620), .A3(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G127gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n624), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n509), .B1(KEYINPUT21), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n629), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n633));
  INV_X1    g432(.A(G155gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G183gat), .B(G211gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n632), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(G230gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n380), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n590), .A2(KEYINPUT105), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n622), .A2(new_n623), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n592), .B2(new_n594), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n622), .A2(new_n623), .A3(new_n641), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n589), .A2(new_n591), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n593), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n643), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n595), .A2(KEYINPUT10), .A3(new_n630), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n640), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n643), .A2(new_n646), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n640), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n651), .A2(new_n653), .A3(new_n657), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n613), .A2(new_n638), .A3(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n484), .A2(new_n574), .A3(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n473), .A2(KEYINPUT106), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n473), .A2(KEYINPUT106), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g469(.A1(new_n664), .A2(new_n428), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n664), .A2(KEYINPUT108), .A3(new_n428), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(G8gat), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n671), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n673), .B2(new_n674), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n675), .B(new_n678), .C1(new_n679), .C2(new_n680), .ZN(G1325gat));
  INV_X1    g480(.A(new_n466), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n664), .A2(new_n493), .A3(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n664), .A2(new_n468), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n493), .ZN(G1326gat));
  NAND2_X1  g484(.A1(new_n664), .A2(new_n476), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NOR2_X1   g487(.A1(new_n484), .A2(new_n574), .ZN(new_n689));
  INV_X1    g488(.A(new_n613), .ZN(new_n690));
  INV_X1    g489(.A(new_n638), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n691), .A3(new_n662), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT109), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G29gat), .A3(new_n667), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT45), .Z(new_n696));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n484), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n480), .A2(new_n483), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n300), .A2(new_n470), .A3(new_n287), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n282), .A2(new_n288), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n301), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n476), .B1(new_n702), .B2(new_n428), .ZN(new_n703));
  INV_X1    g502(.A(new_n468), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n303), .A2(new_n377), .A3(new_n376), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n412), .B1(new_n429), .B2(new_n413), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT111), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n698), .A2(new_n709), .A3(new_n710), .A4(new_n690), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n613), .B1(new_n699), .B2(new_n707), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n710), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n638), .B(KEYINPUT110), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(new_n571), .A3(new_n661), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n667), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n696), .A2(new_n719), .ZN(G1328gat));
  NOR3_X1   g519(.A1(new_n694), .A2(G36gat), .A3(new_n474), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n718), .B2(new_n474), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1329gat));
  NOR3_X1   g523(.A1(new_n694), .A2(G43gat), .A3(new_n466), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n715), .A2(new_n468), .A3(new_n717), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(G43gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g527(.A1(new_n476), .A2(G50gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n694), .A2(new_n412), .ZN(new_n730));
  OAI22_X1  g529(.A1(new_n718), .A2(new_n729), .B1(G50gat), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g531(.A1(new_n699), .A2(new_n707), .A3(new_n697), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n697), .B1(new_n699), .B2(new_n707), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n690), .A2(new_n691), .A3(new_n568), .A4(new_n662), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n668), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g538(.A(new_n428), .B(KEYINPUT112), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT113), .ZN(G1333gat));
  INV_X1    g545(.A(new_n737), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n466), .B(KEYINPUT114), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n616), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n737), .A2(G71gat), .A3(new_n468), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n476), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT115), .B(G78gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n568), .A2(new_n638), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n662), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n711), .B2(new_n714), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n667), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT51), .B1(new_n712), .B2(new_n756), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n756), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n668), .A2(new_n580), .A3(new_n661), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(G1336gat));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n690), .A2(new_n710), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n733), .A2(new_n734), .A3(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n740), .B(new_n758), .C1(new_n772), .C2(new_n713), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G92gat), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n775));
  INV_X1    g574(.A(new_n740), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n776), .A2(G92gat), .A3(new_n662), .ZN(new_n777));
  AND4_X1   g576(.A1(KEYINPUT51), .A2(new_n708), .A3(new_n690), .A4(new_n756), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n763), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n766), .A2(KEYINPUT116), .A3(new_n777), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n774), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n428), .B(new_n758), .C1(new_n772), .C2(new_n713), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G92gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n786), .B2(new_n779), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n770), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n581), .B1(new_n760), .B2(new_n428), .ZN(new_n789));
  INV_X1    g588(.A(new_n779), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n781), .A3(new_n782), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n792), .A3(KEYINPUT118), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n788), .A2(new_n793), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n761), .B2(new_n704), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n466), .A2(G99gat), .A3(new_n662), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n767), .B2(new_n796), .ZN(G1338gat));
  NAND2_X1  g596(.A1(new_n760), .A2(new_n476), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n412), .A2(G106gat), .A3(new_n662), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n798), .A2(G106gat), .B1(new_n766), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1339gat));
  NOR2_X1   g601(.A1(new_n663), .A2(new_n568), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n648), .A2(new_n640), .A3(new_n649), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n651), .A2(KEYINPUT54), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n650), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT119), .B1(new_n808), .B2(new_n658), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n810), .B(new_n657), .C1(new_n650), .C2(new_n807), .ZN(new_n811));
  OAI211_X1 g610(.A(KEYINPUT55), .B(new_n806), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n660), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(KEYINPUT120), .A3(new_n660), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n806), .B1(new_n809), .B2(new_n811), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n528), .A2(new_n529), .A3(new_n487), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT121), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n540), .B1(new_n552), .B2(new_n528), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n821), .A2(KEYINPUT121), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n560), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n567), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n820), .A2(new_n613), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n567), .A2(new_n661), .A3(new_n826), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n820), .B2(new_n571), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n613), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n804), .B1(new_n831), .B2(new_n716), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(new_n412), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(new_n682), .A3(new_n668), .A4(new_n776), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n834), .A2(new_n226), .A3(new_n574), .ZN(new_n835));
  INV_X1    g634(.A(new_n463), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(new_n836), .A3(new_n668), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n740), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n568), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n835), .B1(new_n839), .B2(new_n226), .ZN(G1340gat));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n230), .A3(new_n661), .ZN(new_n841));
  OAI21_X1  g640(.A(G120gat), .B1(new_n834), .B2(new_n662), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT122), .Z(G1341gat));
  INV_X1    g643(.A(G127gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n838), .A2(new_n845), .A3(new_n638), .ZN(new_n846));
  INV_X1    g645(.A(new_n716), .ZN(new_n847));
  OAI21_X1  g646(.A(G127gat), .B1(new_n834), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(G1342gat));
  OAI21_X1  g648(.A(G134gat), .B1(new_n834), .B2(new_n613), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT123), .Z(new_n851));
  NAND2_X1  g650(.A1(new_n690), .A2(new_n474), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n837), .A2(G134gat), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT56), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(G1343gat));
  INV_X1    g654(.A(G141gat), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n667), .A2(new_n468), .A3(new_n740), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n832), .A2(new_n476), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(KEYINPUT57), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n813), .B1(new_n818), .B2(new_n817), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n563), .A2(KEYINPUT99), .A3(new_n567), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT99), .B1(new_n563), .B2(new_n567), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n690), .B1(new_n864), .B2(new_n829), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n691), .B1(new_n865), .B2(new_n828), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT57), .B(new_n476), .C1(new_n867), .C2(new_n803), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n858), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n856), .B1(new_n869), .B2(new_n568), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n859), .A2(new_n857), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n574), .A2(G141gat), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n856), .B1(new_n869), .B2(new_n573), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n871), .A2(new_n872), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n874), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n873), .A2(new_n874), .B1(new_n875), .B2(new_n877), .ZN(G1344gat));
  NAND2_X1  g677(.A1(new_n869), .A2(new_n661), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n880), .A3(G148gat), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n882));
  OR3_X1    g681(.A1(new_n820), .A2(new_n613), .A3(new_n827), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n816), .A2(new_n819), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT120), .B1(new_n812), .B2(new_n660), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n884), .A2(new_n571), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n829), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n613), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n716), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(KEYINPUT57), .B(new_n476), .C1(new_n889), .C2(new_n803), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT124), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n832), .A2(new_n892), .A3(KEYINPUT57), .A4(new_n476), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n887), .B1(new_n573), .B2(new_n861), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n883), .B1(new_n897), .B2(new_n690), .ZN(new_n898));
  INV_X1    g697(.A(new_n663), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n898), .A2(new_n691), .B1(new_n574), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n895), .B(new_n896), .C1(new_n900), .C2(new_n412), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n574), .A2(new_n899), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n412), .B1(new_n866), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT125), .B1(new_n903), .B2(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n894), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n858), .A2(new_n662), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G148gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n882), .B1(new_n908), .B2(KEYINPUT59), .ZN(new_n909));
  INV_X1    g708(.A(G148gat), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n905), .B2(new_n906), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(KEYINPUT126), .A3(new_n880), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n881), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n906), .A2(new_n910), .A3(new_n859), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1345gat));
  AOI21_X1  g714(.A(G155gat), .B1(new_n871), .B2(new_n638), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n847), .A2(new_n634), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n869), .B2(new_n917), .ZN(G1346gat));
  NAND2_X1  g717(.A1(new_n869), .A2(new_n690), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G162gat), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n852), .A2(new_n468), .A3(G162gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n859), .A2(new_n668), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1347gat));
  NAND2_X1  g722(.A1(new_n667), .A2(new_n428), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n748), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n833), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(G169gat), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n926), .A2(new_n927), .A3(new_n574), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n832), .A2(new_n667), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n478), .A3(new_n740), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n568), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n928), .B1(new_n932), .B2(new_n927), .ZN(G1348gat));
  AOI21_X1  g732(.A(G176gat), .B1(new_n931), .B2(new_n661), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n833), .A2(G176gat), .A3(new_n661), .A4(new_n925), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n926), .B2(new_n847), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n638), .A2(new_n317), .A3(new_n315), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n930), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n926), .B2(new_n613), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT61), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n931), .A2(new_n316), .A3(new_n690), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1351gat));
  NOR2_X1   g746(.A1(new_n924), .A2(new_n468), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n905), .A2(G197gat), .A3(new_n573), .A4(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(G197gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n776), .A2(new_n468), .A3(new_n412), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n929), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n952), .B2(new_n571), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n949), .A2(new_n953), .ZN(G1352gat));
  NOR3_X1   g753(.A1(new_n952), .A2(G204gat), .A3(new_n662), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n905), .A2(new_n661), .A3(new_n948), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G204gat), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1353gat));
  OR3_X1    g758(.A1(new_n952), .A2(new_n350), .A3(new_n691), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n905), .A2(new_n638), .A3(new_n948), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  NAND3_X1  g763(.A1(new_n905), .A2(new_n690), .A3(new_n948), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G218gat), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n613), .A2(G218gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n952), .B2(new_n967), .ZN(G1355gat));
endmodule


