//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT73), .B(G110), .Z(new_n194));
  INV_X1    g008(.A(KEYINPUT74), .ZN(new_n195));
  OR3_X1    g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n193), .B2(new_n194), .ZN(new_n197));
  XNOR2_X1  g011(.A(G119), .B(G128), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  OAI211_X1 g013(.A(new_n196), .B(new_n197), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .A4(KEYINPUT16), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n201), .A3(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT71), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n206), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n202), .A2(new_n204), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n200), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n213), .B(new_n206), .C1(new_n207), .C2(new_n210), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n193), .A2(G110), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n199), .A2(new_n198), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT72), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT72), .ZN(new_n223));
  AOI211_X1 g037(.A(new_n223), .B(new_n220), .C1(new_n212), .C2(new_n216), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n215), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT75), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G137), .ZN(new_n227));
  INV_X1    g041(.A(G953), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  XOR2_X1   g043(.A(new_n227), .B(new_n229), .Z(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n232), .B(new_n215), .C1(new_n222), .C2(new_n224), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n226), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G902), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n217), .A2(new_n221), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n223), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n217), .A2(KEYINPUT72), .A3(new_n221), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(KEYINPUT76), .A3(new_n230), .A4(new_n215), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n230), .B(new_n215), .C1(new_n222), .C2(new_n224), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT76), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n234), .A2(new_n235), .A3(new_n240), .A4(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n240), .A2(new_n243), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(KEYINPUT25), .A3(new_n235), .A4(new_n234), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G217), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G234), .B2(new_n235), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n234), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n251), .A2(G902), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n254), .B(KEYINPUT77), .Z(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT2), .A2(G113), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NOR3_X1   g082(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G116), .B(G119), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n271), .B(new_n266), .C1(new_n268), .C2(new_n269), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n213), .A2(G143), .ZN(new_n277));
  INV_X1    g091(.A(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  NOR2_X1   g095(.A1(KEYINPUT0), .A2(G128), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT64), .ZN(new_n285));
  XNOR2_X1  g099(.A(G143), .B(G146), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(new_n281), .ZN(new_n287));
  AND4_X1   g101(.A1(new_n285), .A2(new_n277), .A3(new_n279), .A4(new_n281), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT65), .ZN(new_n290));
  INV_X1    g104(.A(G137), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT11), .B1(new_n291), .B2(G134), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(G134), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OR2_X1    g108(.A1(KEYINPUT66), .A2(G137), .ZN(new_n295));
  NAND2_X1  g109(.A1(KEYINPUT66), .A2(G137), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT11), .A2(G134), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(KEYINPUT67), .A2(G131), .ZN(new_n299));
  NOR2_X1   g113(.A1(KEYINPUT67), .A2(G131), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n294), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  AND2_X1   g116(.A1(KEYINPUT66), .A2(G137), .ZN(new_n303));
  NOR2_X1   g117(.A1(KEYINPUT66), .A2(G137), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n305), .A2(new_n297), .B1(new_n293), .B2(new_n292), .ZN(new_n306));
  INV_X1    g120(.A(G131), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n302), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n309), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n290), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT1), .B1(new_n278), .B2(G146), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n280), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n286), .A2(G128), .A3(new_n312), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(G134), .B1(new_n295), .B2(new_n296), .ZN(new_n317));
  INV_X1    g131(.A(new_n293), .ZN(new_n318));
  OAI21_X1  g132(.A(G131), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n302), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n276), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT64), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n286), .A2(new_n285), .A3(new_n281), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n323), .A2(new_n324), .B1(new_n280), .B2(new_n283), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n308), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(new_n276), .A3(new_n320), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n321), .C2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n308), .B1(new_n325), .B2(new_n309), .ZN(new_n331));
  INV_X1    g145(.A(new_n310), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n320), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n275), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n330), .B1(new_n334), .B2(new_n327), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT69), .B1(new_n327), .B2(new_n330), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n265), .B(new_n329), .C1(new_n335), .C2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT70), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n326), .A2(KEYINPUT30), .A3(new_n320), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n316), .A2(new_n302), .A3(new_n319), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n294), .A2(new_n298), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G131), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n289), .A2(KEYINPUT65), .B1(new_n344), .B2(new_n302), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n345), .B2(new_n310), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n275), .B(new_n341), .C1(new_n346), .C2(KEYINPUT30), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n264), .A3(new_n327), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT31), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(KEYINPUT31), .A3(new_n264), .A4(new_n327), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT28), .B1(new_n321), .B2(new_n328), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n336), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n354), .A2(KEYINPUT70), .A3(new_n265), .A4(new_n329), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n340), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G472), .A2(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT32), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT32), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n360), .A3(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n328), .A2(KEYINPUT28), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n326), .A2(new_n320), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n275), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n327), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n363), .B1(new_n366), .B2(KEYINPUT28), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n265), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(G902), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n347), .A2(new_n327), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n265), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n368), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n265), .B1(new_n354), .B2(new_n329), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G472), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n259), .B1(new_n362), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G214), .B1(G237), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n379));
  INV_X1    g193(.A(G113), .ZN(new_n380));
  INV_X1    g194(.A(G116), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G119), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n188), .A2(G116), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(G119), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT5), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n274), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT80), .B1(new_n390), .B2(G104), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(G104), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G101), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT3), .B1(new_n393), .B2(G107), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n390), .A3(G104), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n393), .A2(G107), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n398), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n379), .B1(new_n389), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n398), .A2(new_n400), .A3(new_n402), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G101), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n403), .A3(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n406), .B(G101), .C1(new_n408), .C2(new_n409), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n275), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT68), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT2), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n380), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n416), .A2(new_n267), .B1(KEYINPUT2), .B2(G113), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n417), .A2(new_n271), .B1(new_n384), .B2(new_n387), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(KEYINPUT84), .A3(new_n403), .A4(new_n397), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n405), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G122), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n405), .A2(new_n413), .A3(new_n421), .A4(new_n419), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(G125), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT1), .ZN(new_n427));
  AND4_X1   g241(.A1(new_n427), .A2(new_n277), .A3(new_n279), .A4(G128), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n312), .A2(G128), .B1(new_n277), .B2(new_n279), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n203), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G224), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(G953), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n431), .B(new_n433), .Z(new_n434));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n420), .A2(new_n435), .A3(new_n422), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n425), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n425), .A2(KEYINPUT85), .A3(new_n434), .A4(new_n436), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT90), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n433), .B1(new_n426), .B2(new_n430), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT7), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n418), .B1(new_n404), .B2(KEYINPUT86), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n389), .A2(new_n449), .A3(new_n403), .A4(new_n397), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n421), .B(KEYINPUT8), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT7), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n433), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n453), .B2(new_n454), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n426), .A2(new_n430), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT88), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n426), .A2(new_n459), .A3(new_n430), .A4(new_n456), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n447), .A2(new_n452), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n424), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n445), .B(new_n235), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n426), .A2(new_n430), .A3(new_n456), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n465), .A2(new_n459), .B1(new_n446), .B2(KEYINPUT7), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n466), .A2(new_n424), .A3(new_n452), .A4(new_n458), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n445), .B1(new_n467), .B2(new_n235), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n441), .A2(new_n444), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n444), .B1(new_n441), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n378), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT67), .B(G131), .ZN(new_n473));
  INV_X1    g287(.A(G237), .ZN(new_n474));
  AND4_X1   g288(.A1(G143), .A2(new_n474), .A3(new_n228), .A4(G214), .ZN(new_n475));
  AOI21_X1  g289(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT17), .B(new_n473), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT95), .B1(new_n479), .B2(new_n217), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(KEYINPUT94), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n228), .A3(G214), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n278), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n301), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n478), .A3(KEYINPUT17), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT95), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n216), .A4(new_n212), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n483), .A2(new_n484), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n473), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n491), .A2(KEYINPUT17), .A3(new_n485), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n480), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n393), .ZN(new_n496));
  INV_X1    g310(.A(new_n490), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT18), .A2(G131), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n202), .A2(new_n204), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G146), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n497), .A2(new_n498), .B1(new_n214), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n490), .A2(KEYINPUT91), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n483), .A2(new_n504), .A3(new_n484), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n498), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI211_X1 g322(.A(KEYINPUT92), .B(new_n498), .C1(new_n503), .C2(new_n505), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n501), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n494), .A2(new_n496), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n491), .ZN(new_n512));
  INV_X1    g326(.A(new_n485), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT93), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n491), .B2(new_n485), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n499), .B(KEYINPUT19), .Z(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n213), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n514), .A2(new_n212), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n496), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NOR2_X1   g338(.A1(G475), .A2(G902), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT96), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n523), .A2(KEYINPUT96), .A3(new_n524), .A4(new_n525), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n496), .B1(new_n510), .B2(new_n519), .ZN(new_n530));
  INV_X1    g344(.A(new_n501), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT91), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n504), .B1(new_n483), .B2(new_n484), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n507), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT92), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n506), .A2(new_n502), .A3(new_n507), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n531), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n477), .A2(KEYINPUT94), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n478), .B1(new_n485), .B2(KEYINPUT17), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n216), .B(new_n212), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n492), .B1(new_n540), .B2(KEYINPUT95), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n541), .B2(new_n489), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n530), .B1(new_n542), .B2(new_n496), .ZN(new_n543));
  INV_X1    g357(.A(new_n525), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT20), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n528), .A2(new_n529), .A3(new_n545), .ZN(new_n546));
  AOI211_X1 g360(.A(new_n521), .B(new_n537), .C1(new_n541), .C2(new_n489), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n496), .B1(new_n494), .B2(new_n510), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n235), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XOR2_X1   g363(.A(KEYINPUT97), .B(G475), .Z(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G128), .B(G143), .ZN(new_n552));
  INV_X1    g366(.A(G134), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT98), .ZN(new_n555));
  XOR2_X1   g369(.A(G116), .B(G122), .Z(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(G107), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(KEYINPUT13), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n278), .A2(G128), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(G134), .C1(KEYINPUT13), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n555), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n552), .B(new_n553), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n381), .A2(KEYINPUT14), .A3(G122), .ZN(new_n563));
  OAI211_X1 g377(.A(G107), .B(new_n563), .C1(new_n556), .C2(KEYINPUT14), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n562), .B(new_n564), .C1(G107), .C2(new_n556), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT9), .B(G234), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT78), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n568), .A2(new_n250), .A3(G953), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n561), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n569), .B1(new_n561), .B2(new_n565), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n235), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G478), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OAI221_X1 g389(.A(new_n235), .B1(KEYINPUT15), .B2(new_n573), .C1(new_n570), .C2(new_n571), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n228), .A2(G952), .ZN(new_n578));
  NAND2_X1  g392(.A1(G234), .A2(G237), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(G902), .A3(G953), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT21), .B(G898), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n577), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n546), .A2(new_n551), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT82), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n325), .A2(new_n411), .A3(new_n412), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n428), .A2(new_n429), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n590), .B1(new_n404), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n307), .B1(new_n294), .B2(new_n298), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n301), .B2(new_n306), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n316), .A2(KEYINPUT10), .A3(new_n403), .A4(new_n397), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n589), .A2(new_n592), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n404), .A2(new_n591), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n316), .A2(new_n403), .A3(new_n397), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n308), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT12), .B1(new_n308), .B2(KEYINPUT81), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n603));
  INV_X1    g417(.A(new_n601), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n596), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(G110), .B(G140), .ZN(new_n607));
  INV_X1    g421(.A(G227), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(G953), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n607), .B(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n589), .A2(new_n592), .A3(new_n595), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n308), .ZN(new_n612));
  INV_X1    g426(.A(new_n610), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n596), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n606), .A2(new_n610), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n588), .B(G469), .C1(new_n616), .C2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n600), .A2(new_n601), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n603), .A2(new_n604), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT83), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n596), .A2(new_n622), .A3(new_n613), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n618), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n613), .B1(new_n612), .B2(new_n596), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G469), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n628), .A3(new_n235), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n615), .A2(new_n612), .ZN(new_n630));
  INV_X1    g444(.A(new_n611), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n619), .A2(new_n620), .B1(new_n631), .B2(new_n594), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n630), .B(G469), .C1(new_n632), .C2(new_n613), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n628), .A2(new_n235), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n633), .A2(KEYINPUT82), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n617), .A2(new_n629), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(G221), .B1(new_n568), .B2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n472), .A2(new_n587), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n377), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G101), .ZN(G3));
  NAND2_X1  g456(.A1(new_n356), .A2(new_n235), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n643), .A2(G472), .B1(new_n357), .B2(new_n356), .ZN(new_n644));
  INV_X1    g458(.A(new_n251), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n246), .B2(new_n248), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n257), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n637), .A2(new_n638), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n644), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT99), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n644), .A2(new_n647), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT100), .ZN(new_n654));
  INV_X1    g468(.A(new_n585), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n378), .B(new_n655), .C1(new_n470), .C2(new_n471), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n545), .A2(new_n529), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n544), .B1(new_n511), .B2(new_n522), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT96), .B1(new_n658), .B2(new_n524), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n551), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n570), .A2(new_n571), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n573), .A2(G902), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT101), .B(G478), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n663), .A2(new_n664), .B1(new_n572), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n656), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n654), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT34), .B(G104), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G6));
  XOR2_X1   g487(.A(new_n585), .B(KEYINPUT102), .Z(new_n674));
  OAI211_X1 g488(.A(new_n378), .B(new_n674), .C1(new_n470), .C2(new_n471), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n545), .A2(new_n526), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n551), .A3(new_n577), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n654), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT104), .B(G107), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT103), .B(KEYINPUT35), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  NAND2_X1  g497(.A1(new_n643), .A2(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n358), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n226), .A2(new_n233), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n231), .A2(KEYINPUT36), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n256), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n646), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n640), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT37), .B(G110), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G12));
  NOR2_X1   g509(.A1(new_n472), .A2(new_n639), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n356), .A2(new_n360), .A3(new_n357), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n360), .B1(new_n356), .B2(new_n357), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n376), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n646), .A2(new_n690), .ZN(new_n700));
  INV_X1    g514(.A(G900), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n583), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n580), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n677), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n696), .A2(new_n699), .A3(new_n700), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  XNOR2_X1  g521(.A(new_n703), .B(KEYINPUT39), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n648), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n441), .A2(new_n469), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n443), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n441), .A2(new_n469), .A3(new_n444), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT38), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n710), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n366), .A2(new_n265), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n348), .A2(G472), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(G472), .A2(G902), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n721), .B(KEYINPUT105), .Z(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n697), .B2(new_n698), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT106), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n660), .A2(new_n577), .ZN(new_n726));
  INV_X1    g540(.A(new_n378), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n700), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n717), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G143), .ZN(G45));
  AOI211_X1 g544(.A(new_n667), .B(new_n704), .C1(new_n546), .C2(new_n551), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n696), .A2(new_n699), .A3(new_n700), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  AOI22_X1  g547(.A1(KEYINPUT83), .A2(new_n614), .B1(new_n619), .B2(new_n620), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n625), .B1(new_n734), .B2(new_n623), .ZN(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n735), .B2(G902), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n736), .A2(new_n638), .A3(new_n629), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n670), .A2(new_n647), .A3(new_n699), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND4_X1  g554(.A1(new_n678), .A2(new_n647), .A3(new_n699), .A4(new_n737), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  NOR2_X1   g556(.A1(new_n691), .A2(new_n587), .ZN(new_n743));
  INV_X1    g557(.A(new_n737), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n472), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n745), .A3(new_n699), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  OAI211_X1 g561(.A(new_n737), .B(new_n378), .C1(new_n471), .C2(new_n470), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n660), .A2(new_n577), .A3(new_n674), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n252), .A2(KEYINPUT107), .A3(new_n258), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(new_n646), .B2(new_n257), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n352), .B1(new_n264), .B2(new_n367), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n643), .A2(G472), .B1(new_n357), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n750), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  NAND4_X1  g572(.A1(new_n745), .A2(new_n700), .A3(new_n731), .A4(new_n756), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  AOI21_X1  g574(.A(KEYINPUT107), .B1(new_n252), .B2(new_n258), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n646), .A2(new_n752), .A3(new_n257), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n699), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n470), .A2(new_n471), .A3(new_n727), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n616), .A2(KEYINPUT108), .A3(G469), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n633), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n629), .A2(new_n765), .A3(new_n767), .A4(new_n635), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n638), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(KEYINPUT109), .A3(new_n638), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n731), .A2(new_n764), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT42), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n771), .A2(new_n764), .A3(new_n772), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n660), .A2(new_n668), .A3(new_n703), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(KEYINPUT42), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n377), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n307), .ZN(G33));
  NAND3_X1  g594(.A1(new_n377), .A2(new_n775), .A3(new_n705), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G134), .ZN(G36));
  NAND3_X1  g596(.A1(new_n685), .A2(new_n700), .A3(KEYINPUT110), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n644), .B2(new_n691), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n546), .A2(new_n668), .A3(new_n551), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT43), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n546), .A2(new_n668), .A3(new_n789), .A4(new_n551), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n788), .A2(new_n790), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n783), .B2(new_n785), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT112), .B1(new_n797), .B2(KEYINPUT44), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  AOI211_X1 g613(.A(new_n794), .B(new_n796), .C1(new_n785), .C2(new_n783), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n712), .A2(new_n378), .A3(new_n713), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT111), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n629), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n630), .B1(new_n632), .B2(new_n613), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n628), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n616), .A2(KEYINPUT45), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n635), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT46), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n810), .B2(new_n809), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n812), .A2(new_n638), .A3(new_n708), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n814), .B(new_n764), .C1(new_n792), .C2(new_n794), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n799), .A2(new_n802), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  NAND2_X1  g631(.A1(new_n812), .A2(new_n638), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT47), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n699), .A2(new_n647), .A3(new_n801), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n731), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  NOR2_X1   g637(.A1(new_n801), .A2(new_n744), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT120), .ZN(new_n825));
  INV_X1    g639(.A(new_n763), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n796), .A2(new_n580), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT48), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n825), .A2(new_n647), .A3(new_n581), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n660), .A3(new_n668), .A4(new_n724), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n228), .A2(G952), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n581), .A2(new_n791), .A3(new_n756), .A4(new_n754), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n745), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n829), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n715), .A2(new_n378), .A3(new_n744), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n700), .A2(new_n756), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n825), .A2(new_n842), .A3(new_n827), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n736), .A2(new_n629), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n845), .A2(new_n638), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n819), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n833), .A2(new_n764), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n660), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n830), .A2(new_n850), .A3(new_n667), .A4(new_n724), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n841), .A2(new_n843), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n829), .A2(KEYINPUT122), .A3(new_n831), .A4(new_n834), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n837), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n839), .B(KEYINPUT50), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n843), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT121), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n841), .A2(new_n858), .A3(new_n843), .A4(new_n851), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n846), .B1(new_n820), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n819), .A2(KEYINPUT119), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n848), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n857), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n854), .B1(new_n844), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n726), .A2(new_n472), .ZN(new_n866));
  INV_X1    g680(.A(new_n769), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n646), .A2(new_n690), .A3(new_n704), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n866), .A2(new_n723), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n706), .A3(new_n732), .A4(new_n759), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT52), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n774), .A2(new_n778), .A3(new_n781), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n757), .A2(new_n738), .A3(new_n741), .A4(new_n746), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n546), .A2(new_n577), .A3(new_n551), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n675), .B1(new_n669), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n650), .A2(new_n652), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n640), .B1(new_n377), .B2(new_n692), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AND4_X1   g693(.A1(new_n731), .A2(new_n764), .A3(new_n771), .A4(new_n772), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n638), .B(new_n637), .C1(new_n646), .C2(new_n690), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n575), .A2(new_n576), .A3(new_n703), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n549), .B2(new_n550), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n676), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n884), .B1(new_n676), .B2(new_n883), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n881), .A2(new_n887), .A3(new_n801), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n842), .A2(new_n880), .B1(new_n888), .B2(new_n699), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n872), .A2(new_n874), .A3(new_n879), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n871), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n877), .A2(new_n878), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n873), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(new_n872), .A3(KEYINPUT116), .A4(new_n889), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g710(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n757), .A2(new_n738), .A3(new_n746), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(new_n741), .A3(new_n877), .A4(new_n878), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n889), .A2(new_n774), .A3(new_n778), .A4(new_n781), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n891), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n870), .B(KEYINPUT52), .Z(new_n903));
  AND4_X1   g717(.A1(new_n898), .A2(new_n902), .A3(new_n895), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT54), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n903), .A3(new_n895), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n897), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n872), .A2(KEYINPUT53), .A3(new_n879), .A4(new_n889), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n873), .B(KEYINPUT118), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n871), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT54), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n907), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n865), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(G952), .B2(G953), .ZN(new_n915));
  INV_X1    g729(.A(new_n787), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n754), .A2(new_n378), .A3(new_n638), .A4(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT49), .ZN(new_n918));
  INV_X1    g732(.A(new_n845), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n917), .A2(KEYINPUT113), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(KEYINPUT113), .B2(new_n917), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT114), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n715), .B(new_n725), .C1(new_n918), .C2(new_n919), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n915), .A2(new_n926), .ZN(G75));
  AOI21_X1  g741(.A(new_n898), .B1(new_n892), .B2(new_n895), .ZN(new_n928));
  OAI211_X1 g742(.A(G902), .B(new_n443), .C1(new_n928), .C2(new_n910), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n425), .A2(new_n436), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n434), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n929), .B2(new_n930), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n228), .A2(G952), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G51));
  OAI21_X1  g751(.A(KEYINPUT54), .B1(new_n928), .B2(new_n910), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n913), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n634), .B(KEYINPUT57), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n627), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n908), .A2(new_n909), .ZN(new_n943));
  AOI22_X1  g757(.A1(new_n906), .A2(new_n897), .B1(new_n943), .B2(new_n903), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n235), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n807), .A3(new_n806), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n936), .B1(new_n942), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n543), .ZN(new_n949));
  INV_X1    g763(.A(new_n936), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n948), .A2(new_n543), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(G60));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n905), .B2(new_n913), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n950), .B1(new_n956), .B2(new_n663), .ZN(new_n957));
  INV_X1    g771(.A(new_n663), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n955), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT123), .B1(new_n939), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n961));
  INV_X1    g775(.A(new_n959), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n961), .B(new_n962), .C1(new_n938), .C2(new_n913), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n957), .A2(new_n960), .A3(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT60), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n928), .B2(new_n910), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n936), .B1(new_n968), .B2(new_n253), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n688), .A2(new_n689), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n972), .B(new_n967), .C1(new_n928), .C2(new_n910), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n253), .B1(new_n944), .B2(new_n966), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n973), .A3(new_n950), .ZN(new_n976));
  NAND2_X1  g790(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n970), .A2(new_n971), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n974), .A2(new_n979), .ZN(G66));
  OAI21_X1  g794(.A(G953), .B1(new_n584), .B2(new_n432), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n894), .B2(G953), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n931), .B1(G898), .B2(new_n228), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G69));
  MUX2_X1   g798(.A(new_n346), .B(new_n364), .S(KEYINPUT30), .Z(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(new_n517), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n706), .A2(new_n732), .A3(new_n759), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n729), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n729), .A2(KEYINPUT62), .A3(new_n987), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n801), .B(new_n709), .C1(new_n669), .C2(new_n875), .ZN(new_n992));
  AOI22_X1  g806(.A1(new_n990), .A2(new_n991), .B1(new_n377), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n993), .A2(new_n816), .A3(new_n822), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n986), .B1(new_n994), .B2(new_n228), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(G953), .B1(new_n608), .B2(new_n701), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n813), .A2(new_n826), .A3(new_n866), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n872), .A2(new_n987), .A3(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n816), .A2(new_n1000), .A3(new_n228), .A4(new_n822), .ZN(new_n1001));
  INV_X1    g815(.A(new_n986), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(G900), .B2(G953), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n996), .A2(new_n998), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1004), .ZN(new_n1007));
  OAI211_X1 g821(.A(KEYINPUT125), .B(new_n997), .C1(new_n995), .C2(new_n1007), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n1006), .A2(new_n1008), .ZN(G72));
  INV_X1    g823(.A(KEYINPUT127), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n816), .A2(new_n1000), .A3(new_n822), .A4(new_n894), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n720), .B(KEYINPUT63), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT126), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1011), .A2(KEYINPUT126), .A3(new_n1013), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n371), .A2(new_n264), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1010), .B(new_n950), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n371), .A2(new_n264), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n993), .A2(new_n816), .A3(new_n822), .A4(new_n894), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n1023), .B2(new_n1013), .ZN(new_n1024));
  OR2_X1    g838(.A1(new_n896), .A2(new_n904), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1012), .B1(new_n372), .B2(new_n348), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1020), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1028));
  OAI21_X1  g842(.A(KEYINPUT127), .B1(new_n1028), .B2(new_n936), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n1021), .A2(new_n1027), .A3(new_n1029), .ZN(G57));
endmodule


