

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U561 ( .A1(n762), .A2(n740), .ZN(n741) );
  XNOR2_X1 U562 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n746) );
  XNOR2_X1 U563 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U564 ( .A1(G651), .A2(n633), .ZN(n658) );
  XNOR2_X1 U565 ( .A(KEYINPUT86), .B(n540), .ZN(G164) );
  XNOR2_X1 U566 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n529) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XNOR2_X2 U568 ( .A(n529), .B(n528), .ZN(n898) );
  NAND2_X1 U569 ( .A1(G138), .A2(n898), .ZN(n532) );
  INV_X1 U570 ( .A(G2105), .ZN(n535) );
  AND2_X1 U571 ( .A1(n535), .A2(G2104), .ZN(n899) );
  NAND2_X1 U572 ( .A1(n899), .A2(G102), .ZN(n530) );
  XNOR2_X1 U573 ( .A(n530), .B(KEYINPUT84), .ZN(n531) );
  NAND2_X1 U574 ( .A1(n532), .A2(n531), .ZN(n534) );
  INV_X1 U575 ( .A(KEYINPUT85), .ZN(n533) );
  XNOR2_X1 U576 ( .A(n534), .B(n533), .ZN(n539) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  NAND2_X1 U578 ( .A1(G114), .A2(n894), .ZN(n537) );
  NOR2_X1 U579 ( .A1(G2104), .A2(n535), .ZN(n895) );
  NAND2_X1 U580 ( .A1(G126), .A2(n895), .ZN(n536) );
  NAND2_X1 U581 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U582 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U583 ( .A1(n894), .A2(G113), .ZN(n542) );
  NAND2_X1 U584 ( .A1(n898), .A2(G137), .ZN(n541) );
  NAND2_X1 U585 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U586 ( .A(KEYINPUT66), .B(n543), .Z(n545) );
  NAND2_X1 U587 ( .A1(n895), .A2(G125), .ZN(n544) );
  NAND2_X1 U588 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U589 ( .A1(G101), .A2(n899), .ZN(n546) );
  XNOR2_X1 U590 ( .A(KEYINPUT23), .B(n546), .ZN(n547) );
  NOR2_X1 U591 ( .A1(n548), .A2(n547), .ZN(G160) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G108), .ZN(G238) );
  INV_X1 U594 ( .A(G120), .ZN(G236) );
  INV_X1 U595 ( .A(G57), .ZN(G237) );
  INV_X1 U596 ( .A(G132), .ZN(G219) );
  INV_X1 U597 ( .A(G82), .ZN(G220) );
  INV_X1 U598 ( .A(G651), .ZN(n554) );
  NOR2_X1 U599 ( .A1(G543), .A2(n554), .ZN(n550) );
  XNOR2_X1 U600 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n549) );
  XNOR2_X1 U601 ( .A(n550), .B(n549), .ZN(n651) );
  NAND2_X1 U602 ( .A1(G64), .A2(n651), .ZN(n552) );
  XOR2_X1 U603 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  NAND2_X1 U604 ( .A1(G52), .A2(n658), .ZN(n551) );
  NAND2_X1 U605 ( .A1(n552), .A2(n551), .ZN(n560) );
  NOR2_X1 U606 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U607 ( .A1(n652), .A2(G90), .ZN(n553) );
  XNOR2_X1 U608 ( .A(n553), .B(KEYINPUT68), .ZN(n556) );
  NOR2_X1 U609 ( .A1(n633), .A2(n554), .ZN(n653) );
  NAND2_X1 U610 ( .A1(G77), .A2(n653), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U612 ( .A(KEYINPUT69), .B(n557), .ZN(n558) );
  XNOR2_X1 U613 ( .A(KEYINPUT9), .B(n558), .ZN(n559) );
  NOR2_X1 U614 ( .A1(n560), .A2(n559), .ZN(G171) );
  XNOR2_X1 U615 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n566) );
  NAND2_X1 U616 ( .A1(n652), .A2(G89), .ZN(n561) );
  XNOR2_X1 U617 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G76), .A2(n653), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U620 ( .A(n564), .B(KEYINPUT5), .ZN(n565) );
  XNOR2_X1 U621 ( .A(n566), .B(n565), .ZN(n571) );
  NAND2_X1 U622 ( .A1(G63), .A2(n651), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G51), .A2(n658), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U625 ( .A(KEYINPUT6), .B(n569), .ZN(n570) );
  NOR2_X1 U626 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U627 ( .A(KEYINPUT7), .B(KEYINPUT73), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n573), .B(n572), .ZN(G168) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U631 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U632 ( .A(G567), .ZN(n686) );
  NOR2_X1 U633 ( .A1(n686), .A2(G223), .ZN(n575) );
  XNOR2_X1 U634 ( .A(n575), .B(KEYINPUT11), .ZN(G234) );
  XOR2_X1 U635 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n577) );
  NAND2_X1 U636 ( .A1(G56), .A2(n651), .ZN(n576) );
  XNOR2_X1 U637 ( .A(n577), .B(n576), .ZN(n583) );
  NAND2_X1 U638 ( .A1(n652), .A2(G81), .ZN(n578) );
  XNOR2_X1 U639 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G68), .A2(n653), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT13), .B(n581), .Z(n582) );
  NOR2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n658), .A2(G43), .ZN(n584) );
  NAND2_X1 U645 ( .A1(n585), .A2(n584), .ZN(n1011) );
  INV_X1 U646 ( .A(G860), .ZN(n603) );
  OR2_X1 U647 ( .A1(n1011), .A2(n603), .ZN(G153) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U650 ( .A1(G79), .A2(n653), .ZN(n587) );
  NAND2_X1 U651 ( .A1(G54), .A2(n658), .ZN(n586) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G66), .A2(n651), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G92), .A2(n652), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n592), .B(KEYINPUT15), .ZN(n1012) );
  INV_X1 U658 ( .A(G868), .ZN(n670) );
  NAND2_X1 U659 ( .A1(n1012), .A2(n670), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G65), .A2(n651), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G53), .A2(n658), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U664 ( .A1(G91), .A2(n652), .ZN(n598) );
  NAND2_X1 U665 ( .A1(G78), .A2(n653), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n1026) );
  INV_X1 U668 ( .A(n1026), .ZN(G299) );
  NOR2_X1 U669 ( .A1(G286), .A2(n670), .ZN(n602) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U671 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U673 ( .A(n1012), .ZN(n618) );
  NAND2_X1 U674 ( .A1(n604), .A2(n618), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U676 ( .A1(G868), .A2(n1011), .ZN(n608) );
  NAND2_X1 U677 ( .A1(G868), .A2(n618), .ZN(n606) );
  NOR2_X1 U678 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U679 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G123), .A2(n895), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n899), .A2(G99), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G135), .A2(n898), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G111), .A2(n894), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n947) );
  XNOR2_X1 U688 ( .A(G2096), .B(n947), .ZN(n617) );
  INV_X1 U689 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(G156) );
  XNOR2_X1 U691 ( .A(n1011), .B(KEYINPUT74), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n618), .A2(G559), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n620), .B(n619), .ZN(n668) );
  NOR2_X1 U694 ( .A1(n668), .A2(G860), .ZN(n629) );
  NAND2_X1 U695 ( .A1(G67), .A2(n651), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G80), .A2(n653), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G93), .A2(n652), .ZN(n623) );
  XNOR2_X1 U699 ( .A(KEYINPUT75), .B(n623), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n658), .A2(G55), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n671) );
  XOR2_X1 U703 ( .A(n671), .B(KEYINPUT76), .Z(n628) );
  XNOR2_X1 U704 ( .A(n629), .B(n628), .ZN(G145) );
  NAND2_X1 U705 ( .A1(G49), .A2(n658), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U708 ( .A1(n651), .A2(n632), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n633), .A2(G87), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G88), .A2(n652), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G75), .A2(n653), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n642) );
  NAND2_X1 U714 ( .A1(G50), .A2(n658), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n638), .B(KEYINPUT78), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n651), .A2(G62), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U718 ( .A1(n642), .A2(n641), .ZN(G166) );
  NAND2_X1 U719 ( .A1(G61), .A2(n651), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G86), .A2(n652), .ZN(n643) );
  NAND2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G73), .A2(n653), .ZN(n645) );
  XNOR2_X1 U723 ( .A(n645), .B(KEYINPUT2), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n646), .B(KEYINPUT77), .ZN(n647) );
  NOR2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n658), .A2(G48), .ZN(n649) );
  NAND2_X1 U727 ( .A1(n650), .A2(n649), .ZN(G305) );
  AND2_X1 U728 ( .A1(n651), .A2(G60), .ZN(n657) );
  NAND2_X1 U729 ( .A1(G85), .A2(n652), .ZN(n655) );
  NAND2_X1 U730 ( .A1(G72), .A2(n653), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n658), .A2(G47), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(G290) );
  XNOR2_X1 U735 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n662) );
  XNOR2_X1 U736 ( .A(G288), .B(KEYINPUT19), .ZN(n661) );
  XNOR2_X1 U737 ( .A(n662), .B(n661), .ZN(n665) );
  XNOR2_X1 U738 ( .A(G166), .B(G305), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(n671), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(n667) );
  XNOR2_X1 U741 ( .A(G290), .B(n1026), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n667), .B(n666), .ZN(n916) );
  XNOR2_X1 U743 ( .A(n668), .B(n916), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n669), .A2(G868), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U746 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n675), .ZN(n677) );
  XOR2_X1 U750 ( .A(KEYINPUT81), .B(KEYINPUT21), .Z(n676) );
  XNOR2_X1 U751 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U752 ( .A1(n678), .A2(G2072), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n679), .B(KEYINPUT82), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U757 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U758 ( .A1(G96), .A2(n682), .ZN(n851) );
  NAND2_X1 U759 ( .A1(G2106), .A2(n851), .ZN(n683) );
  XNOR2_X1 U760 ( .A(n683), .B(KEYINPUT83), .ZN(n688) );
  NOR2_X1 U761 ( .A1(G236), .A2(G238), .ZN(n684) );
  NAND2_X1 U762 ( .A1(G69), .A2(n684), .ZN(n685) );
  NOR2_X1 U763 ( .A1(G237), .A2(n685), .ZN(n853) );
  NOR2_X1 U764 ( .A1(n686), .A2(n853), .ZN(n687) );
  NOR2_X1 U765 ( .A1(n688), .A2(n687), .ZN(G319) );
  INV_X1 U766 ( .A(G319), .ZN(n690) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U768 ( .A1(n690), .A2(n689), .ZN(n848) );
  NAND2_X1 U769 ( .A1(n848), .A2(G36), .ZN(G176) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n785) );
  INV_X1 U772 ( .A(n785), .ZN(n708) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n691) );
  XNOR2_X1 U774 ( .A(n691), .B(KEYINPUT64), .ZN(n784) );
  AND2_X2 U775 ( .A1(n708), .A2(n784), .ZN(n719) );
  INV_X1 U776 ( .A(n719), .ZN(n750) );
  NAND2_X1 U777 ( .A1(G8), .A2(n750), .ZN(n777) );
  NOR2_X1 U778 ( .A1(G1981), .A2(G305), .ZN(n692) );
  XOR2_X1 U779 ( .A(n692), .B(KEYINPUT24), .Z(n693) );
  NOR2_X1 U780 ( .A1(n777), .A2(n693), .ZN(n783) );
  XOR2_X1 U781 ( .A(G1981), .B(G305), .Z(n1020) );
  INV_X1 U782 ( .A(KEYINPUT98), .ZN(n694) );
  OR2_X1 U783 ( .A1(n694), .A2(n777), .ZN(n696) );
  NAND2_X1 U784 ( .A1(G288), .A2(G1976), .ZN(n695) );
  XNOR2_X1 U785 ( .A(n695), .B(KEYINPUT97), .ZN(n1035) );
  NOR2_X1 U786 ( .A1(n696), .A2(n1035), .ZN(n697) );
  NOR2_X1 U787 ( .A1(KEYINPUT33), .A2(n697), .ZN(n704) );
  NOR2_X1 U788 ( .A1(G1976), .A2(G288), .ZN(n698) );
  XOR2_X1 U789 ( .A(KEYINPUT96), .B(n698), .Z(n1029) );
  OR2_X1 U790 ( .A1(KEYINPUT98), .A2(n1029), .ZN(n701) );
  INV_X1 U791 ( .A(n1029), .ZN(n767) );
  NAND2_X1 U792 ( .A1(n767), .A2(KEYINPUT33), .ZN(n699) );
  NAND2_X1 U793 ( .A1(n699), .A2(KEYINPUT98), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n777), .A2(n702), .ZN(n703) );
  NOR2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U797 ( .A1(n1020), .A2(n705), .ZN(n773) );
  XNOR2_X1 U798 ( .A(KEYINPUT25), .B(G2078), .ZN(n935) );
  NOR2_X1 U799 ( .A1(n750), .A2(n935), .ZN(n707) );
  INV_X1 U800 ( .A(G1961), .ZN(n1015) );
  NOR2_X1 U801 ( .A1(n719), .A2(n1015), .ZN(n706) );
  NOR2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n743) );
  NAND2_X1 U803 ( .A1(G171), .A2(n743), .ZN(n738) );
  AND2_X1 U804 ( .A1(n708), .A2(G1996), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n784), .A2(n709), .ZN(n710) );
  XOR2_X1 U806 ( .A(n710), .B(KEYINPUT26), .Z(n711) );
  NOR2_X1 U807 ( .A1(n1011), .A2(n711), .ZN(n713) );
  NAND2_X1 U808 ( .A1(G1341), .A2(n750), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n728) );
  NOR2_X1 U810 ( .A1(n728), .A2(n1012), .ZN(n714) );
  XOR2_X1 U811 ( .A(n714), .B(KEYINPUT92), .Z(n724) );
  NAND2_X1 U812 ( .A1(G1348), .A2(n750), .ZN(n716) );
  NAND2_X1 U813 ( .A1(G2067), .A2(n719), .ZN(n715) );
  NAND2_X1 U814 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U815 ( .A(KEYINPUT93), .B(n717), .Z(n722) );
  NAND2_X1 U816 ( .A1(n719), .A2(G2072), .ZN(n718) );
  XNOR2_X1 U817 ( .A(n718), .B(KEYINPUT27), .ZN(n721) );
  INV_X1 U818 ( .A(G1956), .ZN(n994) );
  NOR2_X1 U819 ( .A1(n994), .A2(n719), .ZN(n720) );
  NOR2_X1 U820 ( .A1(n721), .A2(n720), .ZN(n725) );
  NAND2_X1 U821 ( .A1(n1026), .A2(n725), .ZN(n727) );
  AND2_X1 U822 ( .A1(n722), .A2(n727), .ZN(n723) );
  NAND2_X1 U823 ( .A1(n724), .A2(n723), .ZN(n734) );
  NOR2_X1 U824 ( .A1(n1026), .A2(n725), .ZN(n726) );
  XOR2_X1 U825 ( .A(n726), .B(KEYINPUT28), .Z(n732) );
  INV_X1 U826 ( .A(n727), .ZN(n730) );
  NAND2_X1 U827 ( .A1(n728), .A2(n1012), .ZN(n729) );
  OR2_X1 U828 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U829 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U830 ( .A1(n734), .A2(n733), .ZN(n736) );
  XOR2_X1 U831 ( .A(KEYINPUT29), .B(KEYINPUT94), .Z(n735) );
  XNOR2_X1 U832 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U833 ( .A1(n738), .A2(n737), .ZN(n749) );
  NOR2_X1 U834 ( .A1(G1966), .A2(n777), .ZN(n762) );
  NOR2_X1 U835 ( .A1(G2084), .A2(n750), .ZN(n759) );
  INV_X1 U836 ( .A(n759), .ZN(n739) );
  NAND2_X1 U837 ( .A1(G8), .A2(n739), .ZN(n740) );
  XNOR2_X1 U838 ( .A(n741), .B(KEYINPUT30), .ZN(n742) );
  NOR2_X1 U839 ( .A1(n742), .A2(G168), .ZN(n745) );
  NOR2_X1 U840 ( .A1(G171), .A2(n743), .ZN(n744) );
  NOR2_X1 U841 ( .A1(n745), .A2(n744), .ZN(n747) );
  NAND2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n760) );
  NAND2_X1 U843 ( .A1(n760), .A2(G286), .ZN(n757) );
  INV_X1 U844 ( .A(G8), .ZN(n755) );
  NOR2_X1 U845 ( .A1(G1971), .A2(n777), .ZN(n752) );
  NOR2_X1 U846 ( .A1(G2090), .A2(n750), .ZN(n751) );
  NOR2_X1 U847 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U848 ( .A1(n753), .A2(G303), .ZN(n754) );
  OR2_X1 U849 ( .A1(n755), .A2(n754), .ZN(n756) );
  AND2_X1 U850 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U851 ( .A(n758), .B(KEYINPUT32), .ZN(n766) );
  NAND2_X1 U852 ( .A1(G8), .A2(n759), .ZN(n764) );
  INV_X1 U853 ( .A(n760), .ZN(n761) );
  NOR2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n776) );
  NOR2_X1 U857 ( .A1(G1971), .A2(G303), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n770) );
  INV_X1 U859 ( .A(KEYINPUT33), .ZN(n769) );
  AND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n776), .A2(n771), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n780) );
  NOR2_X1 U863 ( .A1(G2090), .A2(G303), .ZN(n774) );
  NAND2_X1 U864 ( .A1(G8), .A2(n774), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U868 ( .A(KEYINPUT99), .B(n781), .Z(n782) );
  NOR2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n818) );
  NOR2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n830) );
  XNOR2_X1 U871 ( .A(G2067), .B(KEYINPUT37), .ZN(n828) );
  NAND2_X1 U872 ( .A1(G140), .A2(n898), .ZN(n787) );
  NAND2_X1 U873 ( .A1(G104), .A2(n899), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U875 ( .A(KEYINPUT34), .B(n788), .ZN(n793) );
  NAND2_X1 U876 ( .A1(G116), .A2(n894), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G128), .A2(n895), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U879 ( .A(n791), .B(KEYINPUT35), .Z(n792) );
  NOR2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U881 ( .A(KEYINPUT36), .B(n794), .Z(n795) );
  XNOR2_X1 U882 ( .A(KEYINPUT87), .B(n795), .ZN(n912) );
  NOR2_X1 U883 ( .A1(n828), .A2(n912), .ZN(n968) );
  NAND2_X1 U884 ( .A1(n830), .A2(n968), .ZN(n826) );
  NAND2_X1 U885 ( .A1(G105), .A2(n899), .ZN(n796) );
  XNOR2_X1 U886 ( .A(n796), .B(KEYINPUT38), .ZN(n803) );
  NAND2_X1 U887 ( .A1(G141), .A2(n898), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G117), .A2(n894), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U890 ( .A1(G129), .A2(n895), .ZN(n799) );
  XNOR2_X1 U891 ( .A(KEYINPUT89), .B(n799), .ZN(n800) );
  NOR2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U894 ( .A(KEYINPUT90), .B(n804), .ZN(n883) );
  NAND2_X1 U895 ( .A1(G1996), .A2(n883), .ZN(n805) );
  XNOR2_X1 U896 ( .A(n805), .B(KEYINPUT91), .ZN(n814) );
  NAND2_X1 U897 ( .A1(G131), .A2(n898), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G95), .A2(n899), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U900 ( .A(KEYINPUT88), .B(n808), .Z(n812) );
  NAND2_X1 U901 ( .A1(n894), .A2(G107), .ZN(n810) );
  NAND2_X1 U902 ( .A1(G119), .A2(n895), .ZN(n809) );
  AND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n909) );
  AND2_X1 U905 ( .A1(G1991), .A2(n909), .ZN(n813) );
  NOR2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n949) );
  INV_X1 U907 ( .A(n830), .ZN(n815) );
  NOR2_X1 U908 ( .A1(n949), .A2(n815), .ZN(n823) );
  INV_X1 U909 ( .A(n823), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n826), .A2(n816), .ZN(n817) );
  NOR2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n820) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n1031) );
  NAND2_X1 U913 ( .A1(n1031), .A2(n830), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n833) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n883), .ZN(n954) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n909), .ZN(n951) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n951), .A2(n821), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n954), .A2(n824), .ZN(n825) );
  XNOR2_X1 U921 ( .A(KEYINPUT39), .B(n825), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n828), .A2(n912), .ZN(n965) );
  NAND2_X1 U924 ( .A1(n829), .A2(n965), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U927 ( .A(KEYINPUT40), .B(n834), .ZN(G329) );
  XNOR2_X1 U928 ( .A(G2454), .B(G2451), .ZN(n843) );
  XNOR2_X1 U929 ( .A(G2430), .B(G2446), .ZN(n841) );
  XOR2_X1 U930 ( .A(G2435), .B(G2427), .Z(n836) );
  XNOR2_X1 U931 ( .A(KEYINPUT100), .B(G2438), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U933 ( .A(n837), .B(G2443), .Z(n839) );
  XNOR2_X1 U934 ( .A(G1341), .B(G1348), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n843), .B(n842), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n844), .A2(G14), .ZN(n920) );
  XNOR2_X1 U939 ( .A(KEYINPUT101), .B(n920), .ZN(G401) );
  INV_X1 U940 ( .A(G223), .ZN(n845) );
  NAND2_X1 U941 ( .A1(n845), .A2(G2106), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n846), .B(KEYINPUT102), .ZN(G217) );
  AND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U944 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n849), .A2(n848), .ZN(n850) );
  XOR2_X1 U947 ( .A(KEYINPUT103), .B(n850), .Z(G188) );
  INV_X1 U949 ( .A(G96), .ZN(G221) );
  INV_X1 U950 ( .A(n851), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(G261) );
  INV_X1 U952 ( .A(G261), .ZN(G325) );
  XOR2_X1 U953 ( .A(KEYINPUT41), .B(G1956), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1981), .B(G1966), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U956 ( .A(n856), .B(G2474), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U959 ( .A(G1976), .B(G1971), .Z(n860) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1961), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U963 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(G229) );
  XOR2_X1 U965 ( .A(G2096), .B(KEYINPUT43), .Z(n866) );
  XNOR2_X1 U966 ( .A(G2090), .B(G2678), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(n867), .B(KEYINPUT104), .Z(n869) );
  XNOR2_X1 U969 ( .A(G2067), .B(G2072), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U971 ( .A(KEYINPUT42), .B(G2100), .Z(n871) );
  XNOR2_X1 U972 ( .A(G2078), .B(G2084), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(G227) );
  NAND2_X1 U975 ( .A1(G112), .A2(n894), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G100), .A2(n899), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT107), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G136), .A2(n898), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n895), .A2(G124), .ZN(n879) );
  XOR2_X1 U982 ( .A(KEYINPUT44), .B(n879), .Z(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U984 ( .A(KEYINPUT108), .B(n882), .ZN(G162) );
  XNOR2_X1 U985 ( .A(n883), .B(G164), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n884), .B(G162), .ZN(n908) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n893) );
  NAND2_X1 U988 ( .A1(G139), .A2(n898), .ZN(n886) );
  NAND2_X1 U989 ( .A1(G103), .A2(n899), .ZN(n885) );
  NAND2_X1 U990 ( .A1(n886), .A2(n885), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G115), .A2(n894), .ZN(n888) );
  NAND2_X1 U992 ( .A1(G127), .A2(n895), .ZN(n887) );
  NAND2_X1 U993 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U995 ( .A1(n891), .A2(n890), .ZN(n959) );
  XNOR2_X1 U996 ( .A(n959), .B(n947), .ZN(n892) );
  XNOR2_X1 U997 ( .A(n893), .B(n892), .ZN(n906) );
  NAND2_X1 U998 ( .A1(G118), .A2(n894), .ZN(n897) );
  NAND2_X1 U999 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U1000 ( .A1(n897), .A2(n896), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G142), .A2(n898), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(G106), .A2(n899), .ZN(n900) );
  NAND2_X1 U1003 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U1004 ( .A(n902), .B(KEYINPUT45), .Z(n903) );
  NOR2_X1 U1005 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1006 ( .A(n906), .B(n905), .Z(n907) );
  XOR2_X1 U1007 ( .A(n908), .B(n907), .Z(n911) );
  XOR2_X1 U1008 ( .A(G160), .B(n909), .Z(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n914), .ZN(G395) );
  XNOR2_X1 U1012 ( .A(G286), .B(G301), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(n915), .B(n1011), .ZN(n918) );
  XOR2_X1 U1014 ( .A(n1012), .B(n916), .Z(n917) );
  XNOR2_X1 U1015 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n919), .ZN(G397) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n920), .ZN(n921) );
  XOR2_X1 U1018 ( .A(KEYINPUT109), .B(n921), .Z(n924) );
  NOR2_X1 U1019 ( .A1(G229), .A2(G227), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n922), .B(KEYINPUT49), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT110), .B(n925), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1027 ( .A(G2090), .B(G35), .Z(n941) );
  XOR2_X1 U1028 ( .A(KEYINPUT53), .B(KEYINPUT114), .Z(n939) );
  XNOR2_X1 U1029 ( .A(G2067), .B(G26), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(G33), .B(G2072), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n934) );
  XOR2_X1 U1032 ( .A(G25), .B(G1991), .Z(n930) );
  NAND2_X1 U1033 ( .A1(n930), .A2(G28), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(G32), .B(G1996), .ZN(n931) );
  NOR2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n937) );
  XOR2_X1 U1037 ( .A(G27), .B(n935), .Z(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n939), .B(n938), .ZN(n940) );
  NAND2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G34), .B(G2084), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(n942), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n976) );
  NAND2_X1 U1044 ( .A1(KEYINPUT55), .A2(n976), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(G11), .A2(n945), .ZN(n975) );
  INV_X1 U1046 ( .A(G29), .ZN(n973) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(KEYINPUT113), .ZN(n970) );
  XOR2_X1 U1048 ( .A(G2084), .B(G160), .Z(n946) );
  NOR2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G2090), .B(KEYINPUT111), .ZN(n952) );
  XNOR2_X1 U1053 ( .A(n952), .B(G162), .ZN(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n956) );
  XOR2_X1 U1055 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n955) );
  XNOR2_X1 U1056 ( .A(n956), .B(n955), .ZN(n957) );
  NAND2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n964) );
  XOR2_X1 U1058 ( .A(G2072), .B(n959), .Z(n961) );
  XOR2_X1 U1059 ( .A(G164), .B(G2078), .Z(n960) );
  NOR2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1061 ( .A(KEYINPUT50), .B(n962), .Z(n963) );
  NOR2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(n970), .B(n969), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n971), .A2(KEYINPUT55), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n980) );
  INV_X1 U1069 ( .A(n976), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(G29), .A2(KEYINPUT55), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n1043) );
  XNOR2_X1 U1073 ( .A(G5), .B(G1961), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n981), .B(KEYINPUT119), .ZN(n993) );
  XOR2_X1 U1075 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n988) );
  XNOR2_X1 U1076 ( .A(G1986), .B(G24), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(G23), .B(G1976), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1079 ( .A(G1971), .B(KEYINPUT124), .Z(n984) );
  XNOR2_X1 U1080 ( .A(G22), .B(n984), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(n988), .B(n987), .ZN(n991) );
  XOR2_X1 U1083 ( .A(G1966), .B(G21), .Z(n989) );
  XNOR2_X1 U1084 ( .A(KEYINPUT123), .B(n989), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n1007) );
  XNOR2_X1 U1087 ( .A(n994), .B(G20), .ZN(n1003) );
  XOR2_X1 U1088 ( .A(G1341), .B(G19), .Z(n998) );
  XOR2_X1 U1089 ( .A(KEYINPUT59), .B(KEYINPUT121), .Z(n995) );
  XNOR2_X1 U1090 ( .A(G4), .B(n995), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(n996), .B(G1348), .ZN(n997) );
  NAND2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(KEYINPUT120), .B(G1981), .ZN(n999) );
  XNOR2_X1 U1094 ( .A(G6), .B(n999), .ZN(n1000) );
  NOR2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1097 ( .A(n1004), .B(KEYINPUT122), .ZN(n1005) );
  XNOR2_X1 U1098 ( .A(n1005), .B(KEYINPUT60), .ZN(n1006) );
  NOR2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1100 ( .A(KEYINPUT61), .B(n1008), .Z(n1009) );
  NOR2_X1 U1101 ( .A1(G16), .A2(n1009), .ZN(n1040) );
  XOR2_X1 U1102 ( .A(G16), .B(KEYINPUT56), .Z(n1037) );
  XOR2_X1 U1103 ( .A(G1341), .B(KEYINPUT117), .Z(n1010) );
  XNOR2_X1 U1104 ( .A(n1011), .B(n1010), .ZN(n1014) );
  XNOR2_X1 U1105 ( .A(G1348), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(G303), .B(G1971), .ZN(n1017) );
  XNOR2_X1 U1108 ( .A(n1015), .B(G171), .ZN(n1016) );
  NOR2_X1 U1109 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(G1966), .B(G168), .ZN(n1021) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1113 ( .A(n1022), .B(KEYINPUT57), .ZN(n1023) );
  XNOR2_X1 U1114 ( .A(n1023), .B(KEYINPUT115), .ZN(n1024) );
  NOR2_X1 U1115 ( .A1(n1025), .A2(n1024), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(n1026), .B(G1956), .ZN(n1027) );
  XNOR2_X1 U1117 ( .A(n1027), .B(KEYINPUT116), .ZN(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1119 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1122 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1123 ( .A(n1038), .B(KEYINPUT118), .ZN(n1039) );
  NOR2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1125 ( .A(KEYINPUT126), .B(n1041), .Z(n1042) );
  NOR2_X1 U1126 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XNOR2_X1 U1127 ( .A(KEYINPUT62), .B(n1044), .ZN(G311) );
  INV_X1 U1128 ( .A(G311), .ZN(G150) );
endmodule

