//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT79), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G140), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n191), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT80), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G107), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT3), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n199), .A2(KEYINPUT80), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n201), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(G101), .B1(new_n203), .B2(new_n197), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT65), .A3(G143), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n215), .B2(G146), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n217), .A2(new_n218), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n220), .A2(new_n214), .A3(new_n222), .A4(new_n216), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT68), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(KEYINPUT82), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n220), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n213), .A2(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT82), .B1(new_n223), .B2(new_n225), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n212), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n237));
  INV_X1    g051(.A(G134), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G137), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(G137), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT11), .A3(G134), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n239), .A2(new_n242), .A3(new_n245), .A4(new_n240), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n229), .A2(G128), .B1(new_n228), .B2(new_n216), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n224), .A2(KEYINPUT68), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n224), .A2(KEYINPUT68), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n249), .B1(new_n223), .B2(new_n225), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT70), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT10), .A4(new_n212), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n228), .A2(new_n216), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n260), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n220), .A2(new_n214), .A3(new_n216), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n264), .A2(new_n265), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n202), .A2(G107), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n203), .B2(new_n205), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n204), .A2(KEYINPUT3), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n198), .B1(new_n200), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n269), .B(G101), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n268), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n271), .A2(new_n273), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n269), .B1(new_n278), .B2(new_n208), .ZN(new_n279));
  OAI21_X1  g093(.A(G101), .B1(new_n271), .B2(new_n273), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AND4_X1   g095(.A1(new_n277), .A2(new_n280), .A3(new_n209), .A4(KEYINPUT4), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n236), .A2(new_n248), .A3(new_n258), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n256), .A2(new_n211), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n234), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT12), .B1(new_n286), .B2(new_n247), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT12), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n288), .B(new_n248), .C1(new_n234), .C2(new_n285), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n284), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT83), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n195), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT83), .B(new_n284), .C1(new_n287), .C2(new_n289), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n284), .A2(new_n295), .A3(new_n195), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n236), .A2(new_n258), .A3(new_n283), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n247), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n284), .A2(new_n195), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT84), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n294), .A2(G469), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G469), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n287), .A2(new_n289), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(new_n300), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n195), .B1(new_n298), .B2(new_n284), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n304), .B(new_n305), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n304), .A2(new_n305), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n190), .B1(new_n303), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(G113), .B(G122), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(new_n202), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G125), .B(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .A4(G125), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n321), .A3(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT77), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n318), .A2(G146), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT19), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(G125), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n331), .B2(KEYINPUT88), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT88), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n317), .A2(new_n333), .A3(KEYINPUT19), .ZN(new_n334));
  AOI21_X1  g148(.A(G146), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n337));
  INV_X1    g151(.A(G237), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n192), .A3(G214), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n215), .ZN(new_n340));
  NOR2_X1   g154(.A1(G237), .A2(G953), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(G143), .A3(G214), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n337), .B1(new_n343), .B2(G131), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n340), .A2(KEYINPUT87), .A3(new_n245), .A4(new_n342), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(G131), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n336), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(KEYINPUT18), .A3(G131), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n331), .A2(G146), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n317), .A2(new_n213), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(KEYINPUT18), .A2(G131), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n340), .A2(new_n342), .A3(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n349), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT89), .B(new_n316), .C1(new_n348), .C2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT89), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n336), .B2(new_n347), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(new_n315), .ZN(new_n359));
  INV_X1    g173(.A(new_n355), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n347), .A2(KEYINPUT17), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n324), .B(new_n322), .C1(new_n331), .C2(new_n320), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n213), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n343), .A2(KEYINPUT17), .A3(G131), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n325), .A3(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n315), .B(new_n360), .C1(new_n361), .C2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n356), .A2(new_n359), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(G475), .A2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT90), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(KEYINPUT90), .A3(new_n368), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(KEYINPUT20), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT90), .B1(new_n367), .B2(new_n368), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT20), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n360), .B1(new_n361), .B2(new_n365), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT91), .A3(new_n316), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n366), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n362), .A2(new_n213), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n380), .A2(new_n326), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n381), .B(new_n364), .C1(new_n347), .C2(KEYINPUT17), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n315), .B1(new_n382), .B2(new_n360), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n305), .B(new_n377), .C1(new_n379), .C2(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n374), .A2(new_n375), .B1(G475), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n373), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OR2_X1    g201(.A1(KEYINPUT95), .A2(G952), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT95), .A2(G952), .ZN(new_n389));
  AOI21_X1  g203(.A(G953), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(G234), .A2(G237), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(KEYINPUT21), .B(G898), .Z(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(G902), .A3(G953), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT92), .ZN(new_n396));
  INV_X1    g210(.A(G122), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n396), .B1(G116), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G116), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n399), .A2(KEYINPUT92), .A3(G122), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(G122), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n196), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n402), .B1(new_n398), .B2(new_n400), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G107), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT93), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n403), .A2(KEYINPUT93), .A3(new_n405), .ZN(new_n409));
  XNOR2_X1  g223(.A(G128), .B(G143), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT13), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n221), .A2(KEYINPUT13), .A3(G143), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(new_n238), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n411), .A2(new_n413), .B1(new_n238), .B2(new_n410), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n401), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n402), .B(KEYINPUT14), .ZN(new_n417));
  OAI21_X1  g231(.A(G107), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n410), .B(new_n238), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n403), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G217), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n187), .A2(new_n422), .A3(G953), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n415), .A2(new_n420), .A3(new_n423), .ZN(new_n426));
  AOI21_X1  g240(.A(G902), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G478), .ZN(new_n428));
  OAI22_X1  g242(.A1(new_n427), .A2(KEYINPUT94), .B1(KEYINPUT15), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n426), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n423), .B1(new_n415), .B2(new_n420), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n305), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT94), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n428), .A2(KEYINPUT15), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n427), .A2(KEYINPUT94), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n387), .A2(new_n395), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT96), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n387), .A2(KEYINPUT96), .A3(new_n395), .A4(new_n438), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n313), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT32), .ZN(new_n444));
  XNOR2_X1  g258(.A(G116), .B(G119), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT2), .B(G113), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n445), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n450), .A3(KEYINPUT69), .ZN(new_n451));
  OR3_X1    g265(.A1(new_n449), .A2(KEYINPUT69), .A3(new_n445), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n247), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT67), .B1(new_n238), .B2(G137), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n240), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n238), .A2(KEYINPUT67), .A3(G137), .ZN(new_n458));
  OAI21_X1  g272(.A(G131), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n246), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n455), .B1(new_n460), .B2(new_n256), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n255), .A2(new_n464), .A3(new_n257), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n455), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n454), .B(new_n463), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n455), .A2(new_n453), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n223), .A2(new_n225), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT70), .B1(new_n470), .B2(new_n250), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n254), .B(new_n249), .C1(new_n223), .C2(new_n225), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n469), .B1(new_n473), .B2(new_n464), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n341), .A2(G210), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT26), .B(G101), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n468), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT31), .ZN(new_n483));
  INV_X1    g297(.A(new_n455), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n473), .B2(new_n464), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n454), .B1(new_n485), .B2(KEYINPUT73), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT73), .B1(new_n465), .B2(new_n455), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT28), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT72), .ZN(new_n490));
  INV_X1    g304(.A(new_n469), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n465), .A2(new_n491), .B1(new_n461), .B2(new_n454), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n461), .A2(new_n454), .ZN(new_n495));
  OAI211_X1 g309(.A(KEYINPUT72), .B(KEYINPUT28), .C1(new_n474), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n480), .B1(new_n489), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT74), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n465), .A2(KEYINPUT73), .A3(new_n455), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n453), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n493), .B1(new_n501), .B2(new_n487), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n494), .A3(new_n496), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT74), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(new_n480), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n483), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G472), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n305), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n444), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT76), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n508), .A2(new_n444), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n453), .B1(new_n465), .B2(new_n455), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT28), .B1(new_n515), .B2(new_n474), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT75), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n514), .B1(new_n517), .B2(new_n502), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n468), .A2(new_n475), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n480), .B1(new_n519), .B2(KEYINPUT29), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n481), .A2(new_n514), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n520), .B1(new_n503), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n305), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G472), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT31), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n482), .B(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n503), .A2(new_n504), .A3(new_n480), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n504), .B1(new_n503), .B2(new_n480), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT76), .A3(new_n511), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n509), .A2(new_n513), .A3(new_n524), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT78), .ZN(new_n532));
  NAND2_X1  g346(.A1(G221), .A2(G234), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT22), .B1(new_n533), .B2(G953), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT22), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n535), .A2(new_n192), .A3(G221), .A4(G234), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n536), .A3(G137), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(G137), .B1(new_n534), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n539), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT78), .A3(new_n537), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G119), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G128), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n544), .A2(G128), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n545), .B(new_n546), .C1(new_n547), .C2(KEYINPUT23), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G110), .ZN(new_n549));
  XOR2_X1   g363(.A(KEYINPUT24), .B(G110), .Z(new_n550));
  XNOR2_X1  g364(.A(G119), .B(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n363), .B2(new_n325), .ZN(new_n554));
  OAI22_X1  g368(.A1(new_n548), .A2(G110), .B1(new_n550), .B2(new_n551), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n325), .A3(new_n351), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n543), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n553), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n380), .B2(new_n326), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n538), .A2(new_n539), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n556), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n562), .A3(new_n305), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT25), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n558), .A2(new_n562), .A3(new_n565), .A4(new_n305), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n422), .B1(G234), .B2(new_n305), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n558), .A2(new_n562), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n567), .A2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n451), .A2(new_n452), .A3(new_n274), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n575));
  INV_X1    g389(.A(new_n280), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT81), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n279), .A2(new_n277), .A3(new_n280), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT5), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n544), .A3(G116), .ZN(new_n581));
  OAI211_X1 g395(.A(G113), .B(new_n581), .C1(new_n446), .C2(new_n580), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n450), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(new_n211), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(G110), .B(G122), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n586), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n579), .B2(new_n584), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(KEYINPUT6), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n268), .A2(G125), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n591), .B1(G125), .B2(new_n253), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n192), .A2(G224), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n592), .B(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT6), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n596), .B(new_n588), .C1(new_n579), .C2(new_n584), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT85), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n590), .B(new_n595), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n594), .A2(KEYINPUT86), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n592), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n593), .A2(KEYINPUT7), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n586), .B(KEYINPUT8), .Z(new_n607));
  INV_X1    g421(.A(new_n584), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n583), .A2(new_n211), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n585), .B2(new_n586), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n601), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G210), .B1(G237), .B2(G902), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n601), .A2(new_n614), .A3(new_n612), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(G214), .B1(G237), .B2(G902), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n443), .A2(new_n531), .A3(new_n573), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT97), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  NOR2_X1   g438(.A1(new_n506), .A2(new_n508), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n313), .A2(new_n625), .A3(new_n572), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n627), .B1(new_n506), .B2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n529), .A2(KEYINPUT98), .A3(new_n305), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(G472), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n618), .A2(new_n619), .A3(new_n395), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n426), .B2(KEYINPUT99), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n430), .B2(new_n431), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n425), .B(new_n426), .C1(KEYINPUT99), .C2(new_n632), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n428), .A2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT100), .B(G478), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n432), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n386), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n631), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n626), .A2(new_n630), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NAND2_X1  g460(.A1(new_n387), .A2(new_n437), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n631), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n626), .A2(new_n630), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NAND2_X1  g467(.A1(new_n529), .A2(new_n305), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n507), .B1(new_n654), .B2(new_n627), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n625), .B1(new_n655), .B2(new_n629), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n560), .A2(new_n556), .ZN(new_n658));
  OR3_X1    g472(.A1(new_n658), .A2(KEYINPUT36), .A3(new_n543), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n658), .B1(KEYINPUT36), .B2(new_n543), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n570), .A3(new_n660), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n568), .A2(KEYINPUT103), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT103), .B1(new_n568), .B2(new_n661), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n568), .A2(new_n661), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n568), .A2(KEYINPUT103), .A3(new_n661), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(KEYINPUT104), .A3(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n621), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n656), .A2(new_n443), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  OAI21_X1  g488(.A(new_n392), .B1(G900), .B2(new_n394), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT105), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  AND4_X1   g491(.A1(new_n373), .A2(new_n437), .A3(new_n385), .A4(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n670), .A2(new_n618), .A3(new_n678), .A4(new_n619), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n313), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n531), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT106), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n531), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n676), .B(KEYINPUT39), .Z(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n687), .B1(new_n313), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n312), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n292), .A2(new_n293), .B1(new_n299), .B2(new_n301), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n189), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(KEYINPUT40), .A3(new_n688), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n618), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT38), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n386), .A2(new_n619), .A3(new_n437), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n662), .A2(new_n663), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT38), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n618), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n698), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n480), .B1(new_n515), .B2(new_n474), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n482), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n507), .B1(new_n707), .B2(new_n305), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n509), .A2(new_n513), .A3(new_n530), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n696), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  AND3_X1   g526(.A1(new_n386), .A2(new_n641), .A3(new_n677), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n670), .A3(new_n619), .A4(new_n618), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n313), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n531), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT107), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  OAI21_X1  g532(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n188), .A3(new_n309), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n531), .A2(new_n573), .A3(new_n643), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT41), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G113), .ZN(G15));
  NAND4_X1  g539(.A1(new_n531), .A2(new_n573), .A3(new_n648), .A4(new_n722), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NAND2_X1  g541(.A1(new_n441), .A2(new_n442), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n671), .A2(new_n531), .A3(new_n728), .A4(new_n722), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  AOI21_X1  g544(.A(new_n507), .B1(new_n529), .B2(new_n305), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n517), .A2(new_n502), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n480), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n508), .B1(new_n733), .B2(new_n526), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n731), .A2(new_n572), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n697), .A2(new_n699), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n395), .A3(new_n722), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR3_X1   g552(.A1(new_n731), .A2(new_n700), .A3(new_n734), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n386), .A2(new_n641), .A3(new_n677), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n620), .A2(new_n721), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n303), .A2(new_n312), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n616), .A2(new_n617), .A3(new_n619), .A4(new_n188), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n531), .A2(new_n573), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n744), .B1(new_n748), .B2(new_n740), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n529), .A2(new_n511), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n509), .A2(new_n524), .A3(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n573), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n745), .A2(new_n746), .A3(new_n744), .A4(new_n740), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT108), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AND4_X1   g568(.A1(KEYINPUT108), .A2(new_n753), .A3(new_n573), .A4(new_n751), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NAND4_X1  g571(.A1(new_n531), .A2(new_n747), .A3(new_n573), .A4(new_n678), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  INV_X1    g573(.A(new_n641), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT43), .B1(new_n760), .B2(new_n386), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n387), .A2(new_n762), .A3(new_n641), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n763), .A3(new_n701), .ZN(new_n764));
  INV_X1    g578(.A(new_n625), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n764), .B1(new_n630), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT44), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n656), .B2(new_n764), .ZN(new_n773));
  INV_X1    g587(.A(new_n619), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n618), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n188), .ZN(new_n776));
  INV_X1    g590(.A(new_n309), .ZN(new_n777));
  OAI21_X1  g591(.A(G469), .B1(new_n692), .B2(KEYINPUT45), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n294), .A2(KEYINPUT45), .A3(new_n302), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n311), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT46), .B(new_n311), .C1(new_n778), .C2(new_n779), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n776), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n773), .A2(new_n688), .A3(new_n775), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n771), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT110), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n780), .A2(new_n781), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n309), .A3(new_n783), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n789), .B1(new_n791), .B2(new_n188), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n784), .A2(new_n789), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n775), .A2(new_n572), .A3(new_n713), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n531), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NAND2_X1  g612(.A1(new_n698), .A2(new_n704), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n774), .A3(new_n722), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT112), .ZN(new_n801));
  INV_X1    g615(.A(new_n392), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n761), .A2(new_n763), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n735), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(KEYINPUT113), .A3(KEYINPUT50), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n807));
  NAND3_X1  g621(.A1(new_n801), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n720), .A2(new_n309), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n746), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n739), .A2(new_n802), .A3(new_n803), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n710), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n746), .A2(new_n809), .A3(new_n572), .A4(new_n392), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n387), .A3(new_n760), .A4(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n806), .A2(new_n808), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n804), .A2(new_n775), .ZN(new_n816));
  AOI211_X1 g630(.A(KEYINPUT47), .B(new_n776), .C1(new_n782), .C2(new_n783), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n792), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n720), .A2(new_n189), .A3(new_n309), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(KEYINPUT51), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n752), .A2(new_n802), .A3(new_n803), .A4(new_n810), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT48), .Z(new_n825));
  NAND3_X1  g639(.A1(new_n804), .A2(new_n621), .A3(new_n722), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n812), .A2(new_n813), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n826), .B(new_n390), .C1(new_n642), .C2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n823), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n531), .A2(new_n715), .B1(new_n739), .B2(new_n741), .ZN(new_n831));
  INV_X1    g645(.A(new_n745), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n665), .A2(new_n776), .A3(new_n676), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n710), .A2(new_n736), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n685), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n685), .A2(KEYINPUT52), .A3(new_n831), .A4(new_n834), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n387), .A2(new_n670), .A3(new_n438), .A4(new_n677), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n531), .A2(new_n840), .A3(new_n694), .A4(new_n775), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n739), .A2(new_n713), .A3(new_n747), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n758), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n752), .A2(KEYINPUT108), .A3(new_n753), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n753), .A2(new_n751), .A3(new_n573), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT108), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n843), .B1(new_n848), .B2(new_n749), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n672), .A2(new_n723), .A3(new_n726), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n729), .A2(new_n649), .A3(new_n737), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n622), .A2(new_n644), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT111), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n853), .A2(KEYINPUT111), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n849), .A2(new_n852), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n830), .B1(new_n839), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n837), .A2(new_n838), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT53), .A4(new_n849), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n862), .A2(KEYINPUT54), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(KEYINPUT54), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n822), .A2(KEYINPUT51), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n829), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(G952), .B2(G953), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n809), .B(KEYINPUT49), .Z(new_n868));
  NAND3_X1  g682(.A1(new_n573), .A2(new_n619), .A3(new_n190), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n760), .A2(new_n386), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n799), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n867), .B1(new_n710), .B2(new_n871), .ZN(G75));
  AOI21_X1  g686(.A(new_n305), .B1(new_n857), .B2(new_n861), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(G210), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n590), .B1(new_n599), .B2(new_n600), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(new_n595), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT55), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n874), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n878), .B1(new_n874), .B2(new_n875), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n192), .A2(G952), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G51));
  AND2_X1   g696(.A1(new_n863), .A2(new_n864), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n310), .B(KEYINPUT57), .Z(new_n884));
  OAI22_X1  g698(.A1(new_n883), .A2(new_n884), .B1(new_n308), .B2(new_n307), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n778), .A2(new_n779), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT114), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n873), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n881), .B1(new_n885), .B2(new_n888), .ZN(G54));
  NAND2_X1  g703(.A1(KEYINPUT58), .A2(G475), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT115), .Z(new_n891));
  AND3_X1   g705(.A1(new_n873), .A2(new_n367), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n367), .B1(new_n873), .B2(new_n891), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n881), .ZN(G60));
  INV_X1    g708(.A(new_n881), .ZN(new_n895));
  NAND2_X1  g709(.A1(G478), .A2(G902), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT59), .Z(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n863), .B2(new_n864), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n898), .B2(new_n636), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n636), .B2(new_n898), .ZN(G63));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n901));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT60), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n857), .B2(new_n861), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n569), .B(KEYINPUT118), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n895), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n901), .B1(new_n907), .B2(KEYINPUT117), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n909));
  INV_X1    g723(.A(new_n903), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n862), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n881), .B1(new_n911), .B2(new_n905), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n659), .A2(new_n660), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT116), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n903), .B(new_n915), .C1(new_n857), .C2(new_n861), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n909), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n907), .A2(KEYINPUT119), .A3(new_n916), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n908), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT117), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT61), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT119), .B1(new_n907), .B2(new_n916), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n912), .A2(new_n909), .A3(new_n917), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n920), .A2(new_n925), .ZN(G66));
  NAND3_X1  g740(.A1(new_n393), .A2(G224), .A3(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n858), .B2(G953), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n876), .B1(G898), .B2(new_n192), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n928), .B(new_n929), .Z(G69));
  AND3_X1   g744(.A1(new_n531), .A2(new_n680), .A3(new_n683), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n683), .B1(new_n531), .B2(new_n680), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n831), .B(new_n758), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n751), .A2(new_n573), .A3(new_n736), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n784), .A2(new_n935), .A3(KEYINPUT123), .A4(new_n688), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n784), .A2(new_n688), .ZN(new_n938));
  INV_X1    g752(.A(new_n935), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n934), .A2(new_n756), .A3(new_n936), .A4(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n797), .B1(new_n771), .B2(new_n785), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n192), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n192), .A2(G900), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT122), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT120), .Z(new_n948));
  AND2_X1   g762(.A1(new_n332), .A2(new_n334), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n766), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT109), .B1(new_n766), .B2(KEYINPUT44), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n775), .B1(new_n766), .B2(KEYINPUT44), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n938), .ZN(new_n956));
  AOI22_X1  g770(.A1(new_n954), .A2(new_n956), .B1(new_n818), .B2(new_n796), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n831), .B(new_n711), .C1(new_n931), .C2(new_n932), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n685), .A2(KEYINPUT62), .A3(new_n711), .A4(new_n831), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI211_X1 g776(.A(new_n774), .B(new_n618), .C1(new_n647), .C2(new_n642), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n313), .A2(new_n689), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n531), .A2(new_n963), .A3(new_n573), .A4(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n957), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n192), .ZN(new_n967));
  INV_X1    g781(.A(new_n950), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n951), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n967), .A2(KEYINPUT121), .A3(new_n968), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n951), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n971), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n950), .B1(new_n966), .B2(new_n192), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(KEYINPUT121), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n974), .A2(new_n977), .A3(KEYINPUT124), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT121), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n971), .B1(new_n969), .B2(new_n980), .ZN(new_n981));
  AOI22_X1  g795(.A1(KEYINPUT121), .A2(new_n976), .B1(new_n946), .B2(new_n950), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n972), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(KEYINPUT125), .B(new_n972), .C1(new_n978), .C2(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(G72));
  XNOR2_X1  g802(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n507), .A2(new_n305), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n519), .A2(new_n480), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(new_n482), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n881), .B1(new_n862), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n991), .B1(new_n966), .B2(new_n858), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n519), .B(KEYINPUT127), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n996), .A2(new_n481), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n997), .A2(new_n481), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n941), .A2(new_n858), .A3(new_n942), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(new_n992), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n995), .A2(new_n998), .A3(new_n1001), .ZN(G57));
endmodule


