//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT11), .A3(G134), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT66), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(G137), .ZN(new_n194));
  AOI21_X1  g008(.A(G137), .B1(new_n191), .B2(new_n193), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n189), .B(new_n194), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G131), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G134), .ZN(new_n199));
  AOI21_X1  g013(.A(G131), .B1(new_n199), .B2(G137), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(new_n189), .C1(new_n195), .C2(new_n196), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G128), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n205), .B(new_n207), .C1(KEYINPUT1), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G107), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT82), .B1(new_n214), .B2(G104), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT82), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(G104), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G101), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n214), .A2(G104), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT80), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n217), .A2(G107), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT80), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(KEYINPUT80), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n219), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n228), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n227), .A2(new_n232), .A3(KEYINPUT81), .A4(new_n228), .ZN(new_n236));
  AOI211_X1 g050(.A(new_n213), .B(new_n222), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n236), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n228), .B1(new_n227), .B2(new_n232), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n205), .A2(new_n207), .B1(new_n243), .B2(KEYINPUT64), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  OR2_X1    g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G143), .B(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n245), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n239), .B2(new_n240), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n237), .A2(KEYINPUT10), .B1(new_n242), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n222), .B1(new_n235), .B2(new_n236), .ZN(new_n255));
  INV_X1    g069(.A(new_n213), .ZN(new_n256));
  AOI211_X1 g070(.A(KEYINPUT83), .B(KEYINPUT10), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT83), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n238), .A2(new_n256), .A3(new_n221), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT10), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n203), .B(new_n254), .C1(new_n257), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n238), .A2(new_n221), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n213), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n259), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n265), .A2(KEYINPUT84), .A3(new_n266), .A4(new_n202), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n255), .A2(new_n256), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n202), .B1(new_n268), .B2(new_n237), .ZN(new_n269));
  OR2_X1    g083(.A1(new_n266), .A2(KEYINPUT84), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(KEYINPUT84), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n262), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G110), .B(G140), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n275), .A2(G227), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n254), .B1(new_n257), .B2(new_n261), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n202), .ZN(new_n280));
  INV_X1    g094(.A(new_n277), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n262), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n187), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n280), .B2(new_n262), .ZN(new_n286));
  AND4_X1   g100(.A1(new_n262), .A2(new_n267), .A3(new_n272), .A4(new_n281), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n187), .B(new_n284), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT85), .ZN(new_n289));
  INV_X1    g103(.A(new_n262), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT83), .B1(new_n237), .B2(KEYINPUT10), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n259), .A2(new_n258), .A3(new_n260), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n203), .B1(new_n293), .B2(new_n254), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n277), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n262), .A2(new_n272), .A3(new_n267), .A4(new_n281), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT85), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n187), .A4(new_n284), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n285), .B1(new_n289), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G122), .ZN(new_n303));
  INV_X1    g117(.A(G122), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G116), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G107), .ZN(new_n307));
  XNOR2_X1  g121(.A(G116), .B(G122), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(new_n214), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n301), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(G107), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n214), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT91), .ZN(new_n313));
  XNOR2_X1  g127(.A(G128), .B(G143), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT13), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n211), .A2(KEYINPUT13), .A3(G143), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(new_n190), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n315), .A2(new_n317), .B1(new_n199), .B2(new_n314), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n310), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n302), .A2(KEYINPUT14), .A3(G122), .ZN(new_n320));
  OAI211_X1 g134(.A(G107), .B(new_n320), .C1(new_n306), .C2(KEYINPUT14), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n199), .A2(new_n314), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n199), .A2(new_n314), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n321), .B(new_n312), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT75), .B(G217), .Z(new_n326));
  XOR2_X1   g140(.A(KEYINPUT9), .B(G234), .Z(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n275), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n328), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n319), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G902), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G478), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(KEYINPUT15), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT92), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT92), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n319), .A2(new_n324), .A3(new_n330), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n330), .B1(new_n319), .B2(new_n324), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n337), .B(new_n334), .C1(new_n340), .C2(G902), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n284), .B(new_n335), .C1(new_n338), .C2(new_n339), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT93), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n329), .A2(new_n331), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n344), .A2(new_n345), .A3(new_n284), .A4(new_n335), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n336), .A2(new_n341), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(G237), .A2(G953), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(G143), .A3(G214), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(G143), .B1(new_n348), .B2(G214), .ZN(new_n351));
  OAI21_X1  g165(.A(G131), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(G214), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n206), .ZN(new_n354));
  INV_X1    g168(.A(G131), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n349), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT17), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G125), .ZN(new_n360));
  INV_X1    g174(.A(G125), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G140), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n360), .A2(new_n362), .A3(new_n363), .A4(KEYINPUT16), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT16), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT77), .B1(new_n360), .B2(KEYINPUT16), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G146), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n204), .B(new_n364), .C1(new_n365), .C2(new_n366), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n354), .A2(new_n349), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT17), .A3(G131), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n358), .A2(new_n368), .A3(new_n369), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n360), .A2(new_n362), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT90), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT90), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(G146), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n373), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n204), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT18), .A2(G131), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n354), .A2(new_n349), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n370), .A2(KEYINPUT18), .A3(G131), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(G113), .B(G122), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n217), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n372), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT19), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n375), .B2(new_n376), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n378), .A2(KEYINPUT19), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n204), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n352), .A2(new_n356), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n368), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n386), .B1(new_n393), .B2(new_n384), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(G475), .A2(G902), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT20), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT20), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n399), .B(new_n396), .C1(new_n394), .C2(new_n387), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n275), .A2(G952), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(G234), .B2(G237), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT21), .B(G898), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(G234), .A2(G237), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(G902), .A3(G953), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n386), .B1(new_n372), .B2(new_n384), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n284), .B1(new_n387), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G475), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n347), .A2(new_n401), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT94), .ZN(new_n414));
  INV_X1    g228(.A(G221), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n327), .B2(new_n284), .ZN(new_n416));
  OAI21_X1  g230(.A(G214), .B1(G237), .B2(G902), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI211_X1 g233(.A(new_n240), .B(new_n239), .C1(new_n235), .C2(new_n236), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT2), .B(G113), .Z(new_n421));
  INV_X1    g235(.A(KEYINPUT69), .ZN(new_n422));
  XNOR2_X1  g236(.A(G116), .B(G119), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G119), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G116), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n302), .A2(G119), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT2), .B(G113), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT69), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT68), .B1(new_n428), .B2(new_n429), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n421), .A2(new_n433), .A3(new_n423), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n239), .A2(new_n240), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n420), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G113), .B1(new_n426), .B2(KEYINPUT5), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(KEYINPUT5), .B2(new_n423), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT86), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n423), .A2(KEYINPUT5), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n439), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n444), .A3(new_n431), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n263), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n419), .B1(new_n438), .B2(new_n446), .ZN(new_n447));
  OAI221_X1 g261(.A(new_n418), .B1(new_n263), .B2(new_n445), .C1(new_n420), .C2(new_n437), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(KEYINPUT6), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n252), .A2(G125), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n213), .A2(new_n361), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n275), .A2(G224), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT87), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n452), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(new_n419), .C1(new_n438), .C2(new_n446), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n449), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(KEYINPUT7), .ZN(new_n459));
  AOI21_X1  g273(.A(G125), .B1(new_n210), .B2(new_n212), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n244), .A2(new_n248), .B1(new_n245), .B2(new_n250), .ZN(new_n462));
  OAI22_X1  g276(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n361), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n460), .A2(new_n461), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n459), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n450), .A2(new_n451), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT89), .A4(new_n466), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n435), .A2(new_n436), .ZN(new_n472));
  INV_X1    g286(.A(new_n445), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(new_n242), .B1(new_n473), .B2(new_n255), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n471), .B1(new_n418), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n431), .B1(new_n443), .B2(new_n439), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n255), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n418), .B(KEYINPUT8), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n477), .B(new_n478), .C1(new_n255), .C2(new_n445), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n458), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n458), .B2(new_n480), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n417), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR4_X1   g298(.A1(new_n300), .A2(new_n414), .A3(new_n416), .A4(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n326), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(G234), .B2(new_n284), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n368), .A2(new_n369), .ZN(new_n488));
  INV_X1    g302(.A(G110), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT23), .B1(new_n211), .B2(G119), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT76), .B1(new_n425), .B2(G128), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  XOR2_X1   g306(.A(G119), .B(G128), .Z(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G110), .ZN(new_n494));
  OAI221_X1 g308(.A(new_n488), .B1(new_n489), .B2(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n494), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT78), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n492), .A2(new_n489), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n368), .B(new_n379), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT22), .B(G137), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n275), .A2(G221), .A3(G234), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n495), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n495), .B2(new_n499), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT25), .B1(new_n506), .B2(new_n284), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n508));
  NOR4_X1   g322(.A1(new_n504), .A2(new_n505), .A3(new_n508), .A4(G902), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n487), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n487), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n284), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT79), .ZN(new_n513));
  INV_X1    g327(.A(new_n506), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n188), .A2(G134), .ZN(new_n516));
  OAI21_X1  g330(.A(G131), .B1(new_n195), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n189), .B1(new_n195), .B2(new_n196), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n194), .A2(new_n355), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT70), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n201), .A2(new_n522), .A3(new_n517), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n523), .A3(new_n256), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n202), .A2(new_n462), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(KEYINPUT30), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT67), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n213), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(KEYINPUT67), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n528), .A2(new_n529), .B1(new_n202), .B2(new_n462), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n526), .B(new_n435), .C1(KEYINPUT30), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  INV_X1    g346(.A(new_n435), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n524), .A2(new_n533), .A3(new_n525), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n348), .A2(G210), .ZN(new_n535));
  XOR2_X1   g349(.A(new_n535), .B(KEYINPUT27), .Z(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT26), .B(G101), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n536), .B(new_n537), .Z(new_n538));
  NAND4_X1  g352(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT71), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n524), .A2(new_n533), .A3(new_n525), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n520), .A2(new_n527), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n256), .A3(new_n529), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n533), .B1(new_n544), .B2(new_n525), .ZN(new_n545));
  OAI211_X1 g359(.A(KEYINPUT72), .B(KEYINPUT28), .C1(new_n542), .C2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n538), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n525), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n435), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n550), .B2(new_n534), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n534), .A2(new_n548), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT72), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n546), .B(new_n547), .C1(new_n551), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT73), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n531), .A2(new_n534), .A3(new_n538), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT31), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT28), .B1(new_n542), .B2(new_n545), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT72), .B1(new_n534), .B2(new_n548), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n547), .A4(new_n546), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n541), .A2(new_n556), .A3(new_n558), .A4(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT32), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n565), .A2(G472), .A3(G902), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n546), .B1(new_n551), .B2(new_n554), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT29), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n533), .B1(new_n524), .B2(new_n525), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n570), .B(KEYINPUT28), .C1(new_n542), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n524), .A2(new_n525), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n435), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n548), .B1(new_n574), .B2(new_n534), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n552), .A2(KEYINPUT74), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n572), .B(KEYINPUT29), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n569), .A2(new_n538), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n531), .A2(new_n568), .A3(new_n534), .A4(new_n547), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n579), .A2(new_n284), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n564), .A2(new_n566), .B1(new_n581), .B2(G472), .ZN(new_n582));
  NOR2_X1   g396(.A1(G472), .A2(G902), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n556), .A2(new_n558), .A3(new_n563), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n539), .A2(new_n540), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n539), .A2(new_n540), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n565), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n515), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n485), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  OAI21_X1  g406(.A(new_n284), .B1(new_n584), .B2(new_n587), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(G472), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n588), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n593), .B2(G472), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n300), .A2(new_n515), .A3(new_n416), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n409), .B(new_n417), .C1(new_n482), .C2(new_n483), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n340), .B(KEYINPUT33), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G478), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n332), .A2(new_n333), .ZN(new_n604));
  NAND2_X1  g418(.A1(G478), .A2(G902), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n401), .A2(new_n412), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n600), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  INV_X1    g427(.A(new_n347), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n398), .A2(new_n400), .B1(G475), .B2(new_n411), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n601), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n600), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT35), .B(G107), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  INV_X1    g434(.A(new_n596), .ZN(new_n621));
  INV_X1    g435(.A(new_n597), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n502), .A2(KEYINPUT36), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n495), .A2(new_n499), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n495), .B2(new_n499), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n513), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR4_X1   g443(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT96), .A4(new_n513), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n510), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n621), .A2(new_n485), .A3(new_n622), .A4(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  NAND2_X1  g449(.A1(new_n581), .A2(G472), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n566), .B1(new_n584), .B2(new_n587), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT32), .B1(new_n564), .B2(new_n583), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n632), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n289), .A2(new_n299), .ZN(new_n641));
  INV_X1    g455(.A(new_n285), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n416), .ZN(new_n644));
  INV_X1    g458(.A(new_n417), .ZN(new_n645));
  INV_X1    g459(.A(new_n483), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n458), .A2(new_n480), .A3(new_n481), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n404), .B1(G900), .B2(new_n408), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT97), .Z(new_n650));
  NOR2_X1   g464(.A1(new_n616), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n643), .A2(new_n644), .A3(new_n648), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n640), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n211), .ZN(G30));
  AND2_X1   g468(.A1(new_n531), .A2(new_n534), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n547), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n574), .A2(new_n534), .A3(new_n547), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n284), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n637), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n639), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n646), .A2(new_n647), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n646), .A2(new_n647), .A3(new_n663), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n632), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(new_n608), .A3(new_n614), .A4(new_n417), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n661), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n300), .A2(new_n416), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n650), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT99), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT99), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n672), .A2(new_n676), .A3(new_n673), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(KEYINPUT40), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n676), .A2(new_n643), .A3(new_n644), .A4(new_n673), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n676), .B1(new_n672), .B2(new_n673), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n671), .B1(new_n678), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n206), .ZN(G45));
  INV_X1    g498(.A(new_n650), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n607), .A2(new_n608), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n643), .A2(new_n644), .A3(new_n648), .A4(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n640), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n204), .ZN(G48));
  NAND2_X1  g504(.A1(new_n297), .A2(new_n284), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n289), .A2(new_n299), .B1(G469), .B2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n692), .A2(new_n610), .A3(new_n644), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n590), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT100), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n694), .B(new_n696), .ZN(G15));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  INV_X1    g512(.A(new_n515), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n638), .B2(new_n639), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n692), .A2(new_n617), .A3(new_n644), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n692), .A2(new_n617), .A3(new_n644), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n590), .A2(new_n703), .A3(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  AOI21_X1  g520(.A(new_n668), .B1(new_n582), .B2(new_n589), .ZN(new_n707));
  INV_X1    g521(.A(new_n414), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n691), .A2(G469), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n641), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n416), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n707), .A2(new_n708), .A3(new_n648), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NAND3_X1  g527(.A1(new_n608), .A2(new_n614), .A3(KEYINPUT104), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n615), .B2(new_n347), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n601), .A2(new_n717), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n692), .A2(new_n718), .A3(new_n644), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n572), .B(new_n547), .C1(new_n575), .C2(new_n576), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n558), .ZN(new_n721));
  OAI22_X1  g535(.A1(new_n721), .A2(KEYINPUT102), .B1(new_n585), .B2(new_n586), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n720), .B2(new_n558), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n583), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n725), .A2(new_n726), .B1(new_n593), .B2(G472), .ZN(new_n727));
  OAI211_X1 g541(.A(KEYINPUT103), .B(new_n583), .C1(new_n722), .C2(new_n724), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n719), .A2(new_n727), .A3(new_n699), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NAND4_X1  g544(.A1(new_n641), .A2(new_n644), .A3(new_n648), .A4(new_n709), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n686), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n632), .A3(new_n728), .A4(new_n727), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n646), .A2(new_n417), .A3(new_n647), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n643), .A2(new_n644), .A3(new_n687), .A4(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n735), .B1(new_n700), .B2(new_n738), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n300), .A2(new_n416), .A3(new_n686), .A4(new_n736), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n590), .A3(KEYINPUT42), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND4_X1  g557(.A1(new_n643), .A2(new_n644), .A3(new_n651), .A4(new_n737), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n700), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n190), .ZN(G36));
  INV_X1    g560(.A(new_n641), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n187), .A2(new_n284), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n187), .B1(new_n283), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n262), .A2(new_n281), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n753), .A2(new_n280), .B1(new_n273), .B2(new_n277), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT105), .B1(new_n754), .B2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n278), .A2(KEYINPUT45), .A3(new_n282), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT105), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n750), .B(new_n752), .C1(new_n755), .C2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n754), .A2(KEYINPUT105), .A3(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n756), .A2(new_n757), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n750), .B1(new_n763), .B2(new_n752), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n749), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n747), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n752), .B1(new_n755), .B2(new_n758), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT106), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n748), .B1(new_n769), .B2(new_n759), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT46), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n416), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n772), .A2(new_n673), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n606), .A2(new_n608), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n606), .A2(new_n608), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT108), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n777), .B2(new_n779), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n668), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n597), .B2(new_n596), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n774), .B(new_n737), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n737), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT109), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n786), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n773), .A2(new_n787), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  OAI21_X1  g606(.A(new_n641), .B1(new_n770), .B2(KEYINPUT46), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n766), .B(new_n748), .C1(new_n769), .C2(new_n759), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n644), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n644), .B(new_n799), .C1(new_n793), .C2(new_n794), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n737), .A2(new_n687), .A3(new_n515), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n801), .A2(new_n638), .A3(new_n639), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n798), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  AOI21_X1  g618(.A(new_n745), .B1(new_n739), .B2(new_n741), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n725), .A2(new_n726), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n593), .A2(G472), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n806), .A2(new_n807), .A3(new_n728), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(KEYINPUT111), .A3(new_n632), .A4(new_n740), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n806), .A2(new_n807), .A3(new_n632), .A4(new_n728), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n810), .B1(new_n811), .B2(new_n738), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n615), .A2(new_n347), .A3(new_n685), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n300), .A2(new_n416), .A3(new_n736), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n707), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n805), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n598), .B(new_n599), .C1(new_n610), .C2(new_n617), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n705), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n590), .B1(new_n485), .B2(new_n693), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n633), .A2(new_n820), .A3(new_n712), .A4(new_n729), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n692), .A2(new_n644), .A3(new_n648), .A4(new_n687), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n510), .A2(new_n631), .A3(new_n685), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n484), .A2(new_n717), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n643), .A3(new_n644), .ZN(new_n827));
  OAI22_X1  g641(.A1(new_n811), .A2(new_n824), .B1(new_n827), .B2(new_n661), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n640), .B1(new_n652), .B2(new_n688), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n823), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n300), .A2(new_n416), .A3(new_n484), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n707), .B(new_n831), .C1(new_n651), .C2(new_n687), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n672), .B(new_n826), .C1(new_n639), .C2(new_n660), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n733), .A3(KEYINPUT52), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n817), .A2(new_n822), .A3(KEYINPUT53), .A4(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n643), .A2(new_n708), .A3(new_n644), .A4(new_n648), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n692), .A2(new_n610), .A3(new_n644), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n700), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n640), .A2(new_n414), .A3(new_n731), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n839), .A2(new_n668), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n699), .A2(new_n806), .A3(new_n807), .A4(new_n728), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n598), .A2(new_n844), .B1(new_n845), .B2(new_n719), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n846), .A3(new_n705), .A4(new_n818), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n805), .A2(new_n813), .A3(new_n816), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT113), .A3(KEYINPUT53), .A4(new_n835), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n830), .A2(new_n834), .A3(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(KEYINPUT112), .B(new_n823), .C1(new_n828), .C2(new_n829), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n705), .A2(new_n818), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n633), .A2(new_n820), .A3(new_n712), .A4(new_n729), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n809), .A2(new_n812), .B1(new_n707), .B2(new_n815), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n805), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n851), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n838), .A2(new_n850), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n849), .A2(KEYINPUT53), .A3(new_n854), .A4(new_n853), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  INV_X1    g678(.A(new_n835), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n851), .B1(new_n859), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n863), .A2(new_n866), .A3(KEYINPUT114), .A4(new_n864), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n692), .A2(new_n737), .A3(new_n403), .A4(new_n644), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n871), .A2(new_n780), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n700), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT48), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n661), .A2(new_n699), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n875), .A2(new_n609), .A3(new_n871), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n402), .B(KEYINPUT116), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n403), .B1(new_n777), .B2(new_n779), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n845), .A2(new_n711), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n874), .B(new_n878), .C1(new_n484), .C2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n845), .A2(new_n737), .A3(new_n880), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n800), .B1(new_n772), .B2(new_n796), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n710), .A2(new_n644), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT50), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n727), .A2(new_n699), .A3(new_n728), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n692), .A2(new_n644), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n665), .A2(new_n645), .A3(new_n666), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n889), .A2(new_n890), .A3(new_n879), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n888), .B1(new_n892), .B2(KEYINPUT115), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n872), .A2(new_n811), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n606), .A2(new_n615), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n875), .A2(new_n871), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT115), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n898), .B(KEYINPUT50), .C1(new_n881), .C2(new_n891), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n893), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT51), .B1(new_n887), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n893), .A2(new_n897), .A3(new_n899), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT51), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n885), .B1(new_n798), .B2(new_n800), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n902), .B(new_n903), .C1(new_n904), .C2(new_n883), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n882), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n862), .A2(new_n869), .A3(new_n870), .A4(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(G952), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n275), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n515), .A2(new_n416), .A3(new_n645), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n667), .A2(new_n775), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(KEYINPUT49), .B2(new_n710), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n913), .B(new_n661), .C1(KEYINPUT49), .C2(new_n710), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT117), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n910), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(G75));
  AND2_X1   g733(.A1(new_n863), .A2(new_n866), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n284), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(G210), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n449), .A2(new_n457), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n455), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT55), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n922), .B2(new_n923), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n908), .A2(G953), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT118), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(G51));
  NAND2_X1  g746(.A1(new_n863), .A2(new_n866), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT54), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n867), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n748), .B(KEYINPUT57), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n297), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n921), .A2(new_n759), .A3(new_n769), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n931), .B1(new_n938), .B2(new_n939), .ZN(G54));
  AND3_X1   g754(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n941), .A2(new_n395), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n395), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n931), .B1(new_n942), .B2(new_n943), .ZN(G60));
  XOR2_X1   g758(.A(new_n605), .B(KEYINPUT59), .Z(new_n945));
  AOI211_X1 g759(.A(new_n602), .B(new_n945), .C1(new_n934), .C2(new_n867), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n862), .A2(new_n869), .A3(new_n870), .ZN(new_n947));
  INV_X1    g761(.A(new_n945), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI211_X1 g763(.A(new_n931), .B(new_n946), .C1(new_n602), .C2(new_n949), .ZN(G63));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT60), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT119), .B1(new_n920), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT119), .ZN(new_n955));
  INV_X1    g769(.A(new_n953), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n933), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n957), .A3(new_n514), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n930), .ZN(new_n959));
  INV_X1    g773(.A(new_n627), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n954), .B2(new_n957), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n951), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n961), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n930), .A4(new_n958), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(G66));
  INV_X1    g779(.A(G224), .ZN(new_n966));
  OAI21_X1  g780(.A(G953), .B1(new_n405), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n822), .B2(G953), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n924), .B1(G898), .B2(new_n275), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT120), .Z(new_n970));
  XNOR2_X1  g784(.A(new_n968), .B(new_n970), .ZN(G69));
  OAI21_X1  g785(.A(new_n526), .B1(KEYINPUT30), .B2(new_n530), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n389), .A2(new_n390), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT123), .Z(new_n977));
  NOR3_X1   g791(.A1(new_n680), .A2(new_n681), .A3(new_n679), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT40), .B1(new_n675), .B2(new_n677), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n670), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n832), .A2(new_n733), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n980), .A2(KEYINPUT62), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n683), .B2(new_n981), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n675), .A2(new_n677), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n736), .B1(new_n609), .B2(new_n616), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n590), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n986), .A2(new_n791), .A3(new_n803), .A4(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n977), .B1(new_n992), .B2(new_n275), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n982), .A2(new_n805), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n700), .A2(new_n484), .A3(new_n717), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n994), .B1(new_n773), .B2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n996), .A2(new_n791), .A3(new_n275), .A4(new_n803), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n976), .B1(G900), .B2(G953), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n993), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n275), .B1(G227), .B2(G900), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n999), .B(new_n1000), .Z(G72));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  NAND3_X1  g818(.A1(new_n996), .A2(new_n791), .A3(new_n803), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(new_n847), .ZN(new_n1006));
  INV_X1    g820(.A(new_n655), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1007), .A2(new_n538), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n931), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1004), .B1(new_n992), .B2(new_n847), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT124), .B1(new_n1010), .B2(new_n656), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT124), .ZN(new_n1012));
  INV_X1    g826(.A(new_n656), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n990), .B1(new_n983), .B2(new_n985), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1014), .A2(new_n791), .A3(new_n803), .A4(new_n822), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n1012), .B(new_n1013), .C1(new_n1015), .C2(new_n1004), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1009), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1008), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1018), .A2(new_n1013), .A3(new_n1004), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT125), .Z(new_n1020));
  NAND2_X1  g834(.A1(new_n861), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT126), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n861), .A2(KEYINPUT126), .A3(new_n1020), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1002), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1010), .A2(new_n656), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n1012), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1010), .A2(KEYINPUT124), .A3(new_n656), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1030), .A2(KEYINPUT127), .A3(new_n1031), .A4(new_n1009), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1026), .A2(new_n1032), .ZN(G57));
endmodule


