//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT89), .ZN(new_n189));
  OAI21_X1  g003(.A(G210), .B1(G237), .B2(G902), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n191));
  XOR2_X1   g005(.A(G110), .B(G122), .Z(new_n192));
  XOR2_X1   g006(.A(G116), .B(G119), .Z(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n193), .B(new_n194), .Z(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n197), .A2(new_n200), .A3(new_n205), .A4(new_n201), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n208), .A2(new_n203), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n202), .A2(new_n207), .A3(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT4), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT80), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n210), .A2(KEYINPUT4), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n203), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AOI211_X1 g030(.A(new_n195), .B(new_n204), .C1(new_n212), .C2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT5), .ZN(new_n218));
  INV_X1    g032(.A(G119), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G116), .ZN(new_n220));
  OAI211_X1 g034(.A(G113), .B(new_n220), .C1(new_n193), .C2(new_n218), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n193), .B2(new_n194), .ZN(new_n222));
  INV_X1    g036(.A(new_n201), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n196), .A2(G107), .ZN(new_n224));
  OAI21_X1  g038(.A(G101), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n206), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n191), .B(new_n192), .C1(new_n217), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT85), .ZN(new_n229));
  INV_X1    g043(.A(new_n192), .ZN(new_n230));
  INV_X1    g044(.A(new_n195), .ZN(new_n231));
  INV_X1    g045(.A(new_n204), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n209), .A2(KEYINPUT80), .A3(new_n211), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n214), .B1(new_n213), .B2(new_n215), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n231), .B(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n227), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n230), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT85), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n191), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n229), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n204), .B1(new_n212), .B2(new_n216), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n227), .B1(new_n241), .B2(new_n231), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT84), .B1(new_n242), .B2(new_n230), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n230), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT84), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(new_n192), .C1(new_n217), .C2(new_n227), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n243), .A2(KEYINPUT6), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G146), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT64), .B(G143), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OR2_X1    g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT64), .A2(G143), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT64), .A2(G143), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n256), .A2(new_n257), .A3(G146), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n252), .B(new_n255), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G128), .ZN(new_n266));
  AOI211_X1 g080(.A(new_n249), .B(new_n266), .C1(new_n250), .C2(G146), .ZN(new_n267));
  OR2_X1    g081(.A1(KEYINPUT64), .A2(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT64), .A2(G143), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n259), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n260), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT1), .B1(new_n248), .B2(G146), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n270), .A2(new_n271), .B1(G128), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n264), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n263), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G224), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n277), .B(KEYINPUT86), .Z(new_n278));
  XNOR2_X1  g092(.A(new_n275), .B(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n240), .A2(new_n247), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT87), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n240), .A2(new_n247), .A3(KEYINPUT87), .A4(new_n279), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(KEYINPUT7), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n275), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n226), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n222), .B(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT88), .B(KEYINPUT8), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n192), .B(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n244), .B(new_n286), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n190), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n190), .ZN(new_n296));
  AOI211_X1 g110(.A(new_n296), .B(new_n293), .C1(new_n282), .C2(new_n283), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n189), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n284), .A2(new_n190), .A3(new_n294), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT89), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n188), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G475), .A2(G902), .ZN(new_n302));
  INV_X1    g116(.A(G237), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n248), .A2(new_n303), .A3(new_n276), .A4(G214), .ZN(new_n304));
  INV_X1    g118(.A(G214), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n305), .A2(G237), .A3(G953), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n250), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G131), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(G131), .B(new_n304), .C1(new_n250), .C2(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n264), .A2(G140), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT73), .A4(KEYINPUT16), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n313), .B2(KEYINPUT16), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n315), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G146), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n313), .A2(new_n314), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT19), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n311), .B(new_n320), .C1(new_n323), .C2(G146), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n250), .A2(new_n306), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n325), .A2(KEYINPUT18), .A3(G131), .A4(new_n304), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n321), .B(new_n259), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT18), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n307), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n326), .A2(new_n327), .A3(new_n329), .A4(new_n309), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT90), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G113), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n196), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n324), .A2(KEYINPUT90), .A3(new_n330), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT91), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n319), .B(new_n259), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n325), .A2(KEYINPUT17), .A3(G131), .A4(new_n304), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n340), .B(new_n341), .C1(KEYINPUT17), .C2(new_n311), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n335), .A3(new_n330), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n338), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n339), .B1(new_n338), .B2(new_n343), .ZN(new_n345));
  OAI211_X1 g159(.A(KEYINPUT20), .B(new_n302), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n338), .A2(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n302), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT20), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n342), .A2(new_n330), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n336), .A2(KEYINPUT92), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n351), .B2(new_n352), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G475), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n346), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G122), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G116), .ZN(new_n358));
  INV_X1    g172(.A(G116), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G122), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(new_n199), .ZN(new_n362));
  OAI21_X1  g176(.A(G128), .B1(new_n256), .B2(new_n257), .ZN(new_n363));
  INV_X1    g177(.A(G134), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n363), .B(new_n364), .C1(G128), .C2(new_n248), .ZN(new_n365));
  OAI211_X1 g179(.A(KEYINPUT13), .B(G128), .C1(new_n256), .C2(new_n257), .ZN(new_n366));
  INV_X1    g180(.A(G128), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n268), .B2(new_n269), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT13), .B1(new_n248), .B2(G128), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n366), .B(KEYINPUT93), .C1(new_n368), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n363), .A2(new_n369), .ZN(new_n373));
  OAI21_X1  g187(.A(G134), .B1(new_n373), .B2(KEYINPUT93), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n362), .B(new_n365), .C1(new_n372), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n248), .A2(G128), .ZN(new_n376));
  OAI21_X1  g190(.A(G134), .B1(new_n368), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n365), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n361), .A2(new_n199), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT94), .B1(new_n360), .B2(KEYINPUT14), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n360), .A2(KEYINPUT14), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT94), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT14), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n359), .A4(G122), .ZN(new_n384));
  AND4_X1   g198(.A1(new_n358), .A2(new_n380), .A3(new_n381), .A4(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n378), .B(new_n379), .C1(new_n199), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT9), .B(G234), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n388), .A2(new_n389), .A3(G953), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n375), .A2(new_n386), .A3(new_n390), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT70), .B(G902), .Z(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G478), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n398), .A2(KEYINPUT15), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n397), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(G234), .A2(G237), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n402), .A2(G952), .A3(new_n276), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n395), .A2(G953), .A3(new_n402), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT21), .B(G898), .Z(new_n406));
  OAI21_X1  g220(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n356), .A2(new_n401), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT25), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT22), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(G137), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n413), .B(KEYINPUT75), .Z(new_n414));
  NOR2_X1   g228(.A1(new_n367), .A2(G119), .ZN(new_n415));
  OR3_X1    g229(.A1(new_n219), .A2(KEYINPUT23), .A3(G128), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT23), .B1(new_n219), .B2(G128), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G110), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT24), .B(G110), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n219), .A2(G128), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n420), .A2(new_n423), .B1(new_n259), .B2(new_n321), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n320), .ZN(new_n425));
  OR3_X1    g239(.A1(new_n421), .A2(new_n415), .A3(new_n422), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G110), .B1(new_n418), .B2(new_n427), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n425), .B1(new_n340), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT74), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n425), .B(KEYINPUT74), .C1(new_n340), .C2(new_n430), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n414), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n413), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n435), .A2(new_n395), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n410), .B1(new_n438), .B2(KEYINPUT76), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n434), .ZN(new_n440));
  INV_X1    g254(.A(new_n414), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n437), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n396), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT76), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT25), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n389), .B1(new_n396), .B2(G234), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n439), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n439), .A2(new_n446), .A3(KEYINPUT77), .A4(new_n447), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n435), .A2(new_n437), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n447), .A2(G902), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(G101), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n303), .A2(new_n276), .A3(G210), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT11), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n364), .B2(G137), .ZN(new_n461));
  INV_X1    g275(.A(G137), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(KEYINPUT11), .A3(G134), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n364), .A2(G137), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n461), .A2(new_n463), .A3(new_n308), .A4(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n364), .A2(G137), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n465), .B(new_n468), .C1(new_n267), .C2(new_n273), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n461), .A2(new_n464), .A3(new_n463), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G131), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n254), .A3(new_n261), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n469), .A2(new_n473), .A3(new_n195), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n195), .B1(new_n469), .B2(new_n473), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT28), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(new_n473), .A3(new_n195), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT28), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(KEYINPUT68), .A3(new_n478), .ZN(new_n482));
  AND4_X1   g296(.A1(new_n459), .A2(new_n476), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT69), .B1(new_n483), .B2(KEYINPUT29), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n476), .A2(new_n481), .A3(new_n459), .A4(new_n482), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT29), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n396), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT71), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(KEYINPUT71), .B(new_n396), .C1(new_n484), .C2(new_n488), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n469), .A2(new_n473), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n469), .B2(new_n473), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n231), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT65), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT65), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n498), .B(new_n231), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n474), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n487), .B(new_n485), .C1(new_n500), .C2(new_n459), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n491), .A2(new_n492), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G472), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT67), .ZN(new_n504));
  INV_X1    g318(.A(new_n459), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT66), .B1(new_n474), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n477), .A2(new_n507), .A3(new_n459), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n497), .A2(new_n499), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT31), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n469), .A2(new_n473), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT30), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n469), .A2(new_n473), .A3(new_n493), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n498), .B1(new_n516), .B2(new_n231), .ZN(new_n517));
  INV_X1    g331(.A(new_n499), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n509), .A2(new_n510), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n476), .A2(new_n481), .A3(new_n482), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n505), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n511), .A2(new_n520), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(G472), .A2(G902), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT32), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT32), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n528), .A3(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n455), .B1(new_n503), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G469), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT82), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n367), .B1(new_n270), .B2(KEYINPUT1), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n534), .A2(new_n251), .ZN(new_n535));
  INV_X1    g349(.A(new_n267), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n226), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n287), .A2(new_n267), .A3(new_n273), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n533), .B(new_n472), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT83), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT83), .B(new_n472), .C1(new_n537), .C2(new_n538), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n539), .B2(new_n540), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n241), .A2(new_n262), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n537), .A2(KEYINPUT10), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n287), .B(KEYINPUT10), .C1(new_n267), .C2(new_n273), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n472), .B(KEYINPUT81), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  XOR2_X1   g365(.A(G110), .B(G140), .Z(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT78), .ZN(new_n553));
  INV_X1    g367(.A(G227), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(G953), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n553), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n546), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n472), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n556), .B1(new_n560), .B2(new_n551), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n532), .B(new_n396), .C1(new_n558), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(G469), .A2(G902), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n551), .B1(new_n544), .B2(new_n545), .ZN(new_n564));
  INV_X1    g378(.A(new_n556), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n551), .A3(new_n556), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(G469), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n562), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G221), .B1(new_n388), .B2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n301), .A2(new_n409), .A3(new_n531), .A4(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G101), .ZN(G3));
  AND3_X1   g388(.A1(new_n235), .A2(new_n230), .A3(new_n236), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n192), .B1(new_n217), .B2(new_n227), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(KEYINPUT84), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n191), .B1(new_n237), .B2(new_n245), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n577), .A2(new_n578), .B1(new_n229), .B2(new_n239), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT87), .B1(new_n579), .B2(new_n279), .ZN(new_n580));
  INV_X1    g394(.A(new_n283), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n294), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n296), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n188), .B1(new_n583), .B2(new_n299), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n394), .A2(new_n398), .A3(new_n396), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n375), .A2(new_n386), .A3(new_n390), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n390), .B1(new_n375), .B2(new_n386), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT33), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n392), .A2(new_n589), .A3(new_n393), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n395), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n585), .B1(new_n591), .B2(new_n398), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT95), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n594), .B(new_n585), .C1(new_n591), .C2(new_n398), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n356), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n584), .A2(new_n407), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n524), .A2(new_n396), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n526), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n604), .A2(new_n455), .A3(new_n571), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  NAND2_X1  g422(.A1(new_n346), .A2(new_n355), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n302), .B1(new_n344), .B2(new_n345), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n349), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n584), .A2(new_n401), .A3(new_n407), .A4(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n605), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NOR2_X1   g430(.A1(new_n441), .A2(KEYINPUT36), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(new_n440), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n453), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n450), .A2(new_n451), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n604), .A2(new_n571), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n301), .A2(new_n409), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT37), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n419), .ZN(G12));
  OAI211_X1 g438(.A(new_n187), .B(new_n620), .C1(new_n295), .C2(new_n297), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n609), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n610), .A2(new_n349), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n405), .A2(G900), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n629), .A2(KEYINPUT96), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(KEYINPUT96), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n404), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT97), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n627), .A2(new_n401), .A3(new_n628), .A4(new_n633), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n634), .B(new_n571), .C1(new_n530), .C2(new_n503), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n626), .A2(new_n635), .A3(KEYINPUT98), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n530), .A2(new_n503), .ZN(new_n638));
  INV_X1    g452(.A(new_n634), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n572), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n637), .B1(new_n640), .B2(new_n625), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  NOR2_X1   g457(.A1(new_n297), .A2(new_n189), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n583), .A2(new_n299), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(new_n189), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT38), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n620), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n505), .B1(new_n474), .B2(new_n475), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n519), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n292), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n527), .A2(new_n529), .B1(G472), .B2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n652), .A2(new_n400), .A3(new_n598), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n633), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n572), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT40), .Z(new_n656));
  NAND4_X1  g470(.A1(new_n648), .A2(new_n187), .A3(new_n653), .A4(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(new_n250), .Z(G45));
  AOI21_X1  g472(.A(new_n571), .B1(new_n530), .B2(new_n503), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n596), .A2(new_n356), .A3(new_n633), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n596), .A2(new_n356), .A3(KEYINPUT99), .A4(new_n633), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n584), .A2(new_n659), .A3(new_n620), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n259), .ZN(G48));
  INV_X1    g481(.A(new_n531), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n558), .A2(new_n561), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n396), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G469), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n671), .A2(new_n570), .A3(new_n562), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n601), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND2_X1  g491(.A1(new_n613), .A2(new_n674), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  NAND3_X1  g493(.A1(new_n626), .A2(new_n638), .A3(new_n672), .ZN(new_n680));
  INV_X1    g494(.A(new_n409), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n219), .ZN(G21));
  NOR2_X1   g497(.A1(new_n598), .A2(new_n400), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n584), .A2(KEYINPUT101), .A3(new_n684), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n187), .B(new_n684), .C1(new_n295), .C2(new_n297), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n673), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n455), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n497), .A2(new_n499), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n510), .B1(new_n692), .B2(new_n512), .ZN(new_n693));
  INV_X1    g507(.A(new_n523), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(KEYINPUT100), .B(new_n523), .C1(new_n509), .C2(new_n510), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n521), .A3(new_n696), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n602), .A2(G472), .B1(new_n697), .B2(new_n525), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n690), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n689), .A2(new_n407), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n689), .A2(KEYINPUT102), .A3(new_n407), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT103), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n357), .ZN(G24));
  AND3_X1   g520(.A1(new_n698), .A2(new_n662), .A3(new_n663), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n584), .A2(new_n707), .A3(new_n620), .A4(new_n672), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n626), .A2(KEYINPUT104), .A3(new_n672), .A4(new_n707), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n563), .B(KEYINPUT105), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n562), .A2(new_n568), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n570), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n188), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n298), .A2(new_n300), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n721), .A2(new_n668), .A3(new_n664), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n714), .A2(KEYINPUT42), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n716), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n646), .A2(new_n531), .A3(new_n718), .A4(new_n720), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n715), .B1(new_n726), .B2(new_n664), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  NOR2_X1   g543(.A1(new_n726), .A2(new_n634), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n364), .ZN(G36));
  INV_X1    g545(.A(new_n646), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n188), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n598), .A2(new_n596), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT43), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n604), .A3(new_n620), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n734), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n566), .A2(new_n567), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT46), .B1(new_n743), .B2(new_n717), .ZN(new_n744));
  INV_X1    g558(.A(new_n562), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n717), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n719), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(new_n654), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n740), .B(new_n749), .C1(new_n735), .C2(new_n739), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  XNOR2_X1  g565(.A(new_n748), .B(KEYINPUT47), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n638), .A2(new_n664), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n455), .A3(new_n733), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n450), .A2(new_n718), .A3(new_n451), .A4(new_n619), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n633), .A2(new_n570), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT110), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n757), .A2(KEYINPUT110), .A3(new_n758), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n652), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT101), .B1(new_n584), .B2(new_n684), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n686), .A2(new_n687), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n759), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n666), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n712), .A2(new_n764), .A3(new_n642), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT111), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n666), .B1(new_n636), .B2(new_n641), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n769), .A3(new_n712), .A4(new_n764), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n756), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n767), .A2(new_n756), .A3(new_n770), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n400), .B(KEYINPUT107), .Z(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n598), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n408), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT89), .B1(new_n583), .B2(new_n299), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n187), .B(new_n777), .C1(new_n778), .C2(new_n644), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT108), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n301), .A2(new_n781), .A3(new_n777), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n780), .A2(new_n605), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n301), .A2(new_n407), .A3(new_n599), .A4(new_n605), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n573), .A2(new_n622), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT109), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n573), .A2(new_n784), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n780), .A2(new_n782), .A3(new_n605), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n622), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n659), .A2(new_n298), .A3(new_n187), .A4(new_n300), .ZN(new_n792));
  INV_X1    g606(.A(new_n775), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n611), .A3(new_n633), .ZN(new_n794));
  INV_X1    g608(.A(new_n707), .ZN(new_n795));
  OAI22_X1  g609(.A1(new_n792), .A2(new_n794), .B1(new_n721), .B2(new_n795), .ZN(new_n796));
  AOI221_X4 g610(.A(new_n730), .B1(new_n620), .B2(new_n796), .C1(new_n725), .C2(new_n727), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n678), .B(new_n675), .C1(new_n681), .C2(new_n680), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(new_n702), .B2(new_n703), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n791), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n774), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n768), .A2(new_n712), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(KEYINPUT52), .A3(new_n764), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n773), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n791), .A2(new_n797), .A3(new_n799), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n801), .A2(new_n807), .A3(KEYINPUT54), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n774), .A2(new_n800), .A3(KEYINPUT53), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n806), .B1(new_n804), .B2(new_n805), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(KEYINPUT54), .B2(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n734), .A2(new_n404), .A3(new_n673), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n531), .A3(new_n738), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT48), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n690), .A2(new_n652), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n734), .A2(new_n404), .A3(new_n673), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n599), .ZN(new_n818));
  INV_X1    g632(.A(G952), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n738), .A2(new_n699), .A3(new_n403), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n673), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n819), .B(G953), .C1(new_n821), .C2(new_n584), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n815), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT112), .Z(new_n824));
  AND2_X1   g638(.A1(new_n671), .A2(new_n562), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n752), .B1(new_n719), .B2(new_n825), .ZN(new_n826));
  OR3_X1    g640(.A1(new_n826), .A2(new_n734), .A3(new_n820), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n647), .A2(new_n188), .A3(new_n821), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT50), .Z(new_n829));
  NAND4_X1  g643(.A1(new_n813), .A2(new_n620), .A3(new_n698), .A4(new_n738), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n817), .A2(new_n598), .A3(new_n597), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n827), .A2(new_n829), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT51), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n812), .A2(new_n824), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(G952), .B2(G953), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT49), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n825), .A2(new_n836), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n736), .B(new_n816), .C1(new_n836), .C2(new_n825), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n647), .A2(new_n720), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n839), .ZN(G75));
  NOR2_X1   g654(.A1(new_n801), .A2(new_n807), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n396), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT56), .B1(new_n842), .B2(new_n296), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n579), .B(new_n279), .Z(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT55), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n843), .B(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n276), .A2(G952), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT113), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n846), .A2(new_n848), .ZN(G51));
  XOR2_X1   g663(.A(new_n669), .B(KEYINPUT115), .Z(new_n850));
  XNOR2_X1  g664(.A(new_n841), .B(KEYINPUT54), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n717), .B(KEYINPUT114), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT57), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n850), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n842), .A2(G469), .A3(new_n742), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n847), .B1(new_n854), .B2(new_n855), .ZN(G54));
  NAND3_X1  g670(.A1(new_n842), .A2(KEYINPUT58), .A3(G475), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n344), .A2(new_n345), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n857), .B(new_n858), .Z(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n847), .ZN(G60));
  AND2_X1   g674(.A1(new_n588), .A2(new_n590), .ZN(new_n861));
  NAND2_X1  g675(.A1(G478), .A2(G902), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT59), .Z(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(new_n812), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n848), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n861), .A2(new_n863), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n864), .B(new_n865), .C1(new_n851), .C2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(G63));
  NAND2_X1  g682(.A1(G217), .A2(G902), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT60), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n801), .B2(new_n807), .ZN(new_n872));
  INV_X1    g686(.A(new_n452), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n767), .A2(new_n756), .A3(new_n770), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n771), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n806), .B1(new_n876), .B2(new_n805), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n773), .A2(new_n803), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n800), .A2(KEYINPUT53), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n870), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n618), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n874), .A2(new_n881), .A3(KEYINPUT61), .A4(new_n865), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n883));
  OAI211_X1 g697(.A(KEYINPUT116), .B(new_n865), .C1(new_n880), .C2(new_n452), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n881), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT116), .B1(new_n874), .B2(new_n865), .ZN(new_n886));
  OAI211_X1 g700(.A(KEYINPUT117), .B(new_n883), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n865), .B1(new_n880), .B2(new_n452), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n884), .A3(new_n881), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT117), .B1(new_n892), .B2(new_n883), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n882), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT118), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n896), .B(new_n882), .C1(new_n888), .C2(new_n893), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(new_n897), .ZN(G66));
  AOI21_X1  g712(.A(new_n276), .B1(new_n406), .B2(G224), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n791), .A2(new_n799), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n276), .ZN(new_n901));
  INV_X1    g715(.A(G898), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n579), .B1(new_n902), .B2(G953), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n901), .B(new_n903), .ZN(G69));
  XOR2_X1   g718(.A(new_n802), .B(KEYINPUT121), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n657), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(KEYINPUT122), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n906), .B(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n750), .A2(new_n754), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(KEYINPUT122), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n734), .A2(new_n655), .ZN(new_n912));
  INV_X1    g726(.A(new_n776), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n912), .B(new_n531), .C1(new_n599), .C2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(G953), .ZN(new_n917));
  XOR2_X1   g731(.A(KEYINPUT119), .B(KEYINPUT120), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n323), .B(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n516), .B(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(G900), .ZN(new_n921));
  OAI21_X1  g735(.A(G953), .B1(new_n554), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(G953), .B1(new_n921), .B2(G227), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n730), .B1(new_n725), .B2(new_n727), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n749), .B(new_n531), .C1(new_n762), .C2(new_n763), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n910), .A2(new_n905), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n924), .B1(new_n927), .B2(G953), .ZN(new_n928));
  OAI22_X1  g742(.A1(new_n917), .A2(new_n923), .B1(new_n920), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT123), .ZN(G72));
  NAND2_X1  g744(.A1(G472), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT63), .Z(new_n932));
  NOR2_X1   g746(.A1(new_n500), .A2(new_n459), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT127), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(new_n509), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n811), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n927), .A2(new_n900), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n932), .B(KEYINPUT124), .Z(new_n938));
  OAI211_X1 g752(.A(new_n505), .B(new_n500), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(G952), .B2(new_n276), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT126), .Z(new_n941));
  INV_X1    g755(.A(new_n900), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n938), .B1(new_n916), .B2(new_n942), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n943), .A2(new_n505), .A3(new_n500), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n946));
  AOI211_X1 g760(.A(new_n936), .B(new_n941), .C1(new_n945), .C2(new_n946), .ZN(G57));
endmodule


