//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n539, new_n540, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159, new_n1160;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT67), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(KEYINPUT3), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(G137), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n458), .A2(new_n459), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  NAND3_X1  g047(.A1(new_n460), .A2(new_n467), .A3(new_n462), .ZN(new_n473));
  INV_X1    g048(.A(G136), .ZN(new_n474));
  OR3_X1    g049(.A1(new_n473), .A2(KEYINPUT69), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n460), .A2(new_n462), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n467), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT69), .B1(new_n473), .B2(new_n474), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n475), .A2(new_n478), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT70), .Z(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT71), .ZN(G162));
  NAND4_X1  g059(.A1(new_n460), .A2(G126), .A3(G2105), .A4(new_n462), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n460), .A2(G138), .A3(new_n467), .A4(new_n462), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n491), .A2(new_n492), .A3(new_n467), .A4(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n491), .B2(new_n492), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n490), .A2(KEYINPUT4), .B1(new_n468), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n486), .B1(new_n485), .B2(new_n488), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n489), .A2(new_n495), .A3(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n500));
  XOR2_X1   g075(.A(KEYINPUT74), .B(G651), .Z(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G50), .ZN(new_n503));
  INV_X1    g078(.A(new_n501), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G75), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n498), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT75), .B(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n504), .A2(G62), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n506), .A2(new_n512), .ZN(G166));
  AOI22_X1  g088(.A1(new_n502), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(new_n508), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n502), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n515), .B1(G51), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(G168));
  NAND2_X1  g096(.A1(new_n502), .A2(new_n507), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G90), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(G52), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(new_n501), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(new_n525), .A3(new_n527), .ZN(G301));
  INV_X1    g103(.A(G301), .ZN(G171));
  NAND2_X1  g104(.A1(G68), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G56), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n508), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n517), .A2(G43), .B1(new_n504), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(G81), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  AND3_X1   g111(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G36), .ZN(G176));
  NAND2_X1  g113(.A1(G1), .A2(G3), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT8), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n537), .A2(new_n540), .ZN(G188));
  NAND2_X1  g116(.A1(G78), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G65), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n508), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  INV_X1    g120(.A(G91), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n522), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G53), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n516), .A2(new_n549), .B1(KEYINPUT76), .B2(KEYINPUT9), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT76), .B(KEYINPUT9), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n502), .A2(G53), .A3(G543), .A4(new_n551), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n550), .A2(KEYINPUT77), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(KEYINPUT77), .B1(new_n550), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(G299));
  INV_X1    g130(.A(G168), .ZN(G286));
  INV_X1    g131(.A(G166), .ZN(G303));
  OAI21_X1  g132(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n558));
  INV_X1    g133(.A(G87), .ZN(new_n559));
  INV_X1    g134(.A(G49), .ZN(new_n560));
  OAI221_X1 g135(.A(new_n558), .B1(new_n522), .B2(new_n559), .C1(new_n560), .C2(new_n516), .ZN(G288));
  NAND2_X1  g136(.A1(G73), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G61), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n508), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n517), .A2(G48), .B1(new_n504), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n523), .A2(G86), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(G305));
  AOI22_X1  g142(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT78), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(new_n504), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n517), .A2(G47), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n523), .A2(G85), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G290));
  INV_X1    g148(.A(G868), .ZN(new_n574));
  NOR2_X1   g149(.A1(G171), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT10), .ZN(new_n576));
  INV_X1    g151(.A(G92), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n522), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n502), .A2(KEYINPUT10), .A3(G92), .A4(new_n507), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n516), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n502), .A2(new_n582), .A3(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(G54), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n507), .A2(G66), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT80), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n580), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n580), .A2(new_n584), .A3(KEYINPUT81), .A4(new_n588), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n575), .B1(new_n593), .B2(new_n574), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT82), .ZN(G284));
  XOR2_X1   g170(.A(new_n594), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g171(.A1(G299), .A2(new_n574), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n574), .B2(G168), .ZN(G280));
  XOR2_X1   g173(.A(G280), .B(KEYINPUT84), .Z(G297));
  INV_X1    g174(.A(new_n593), .ZN(new_n600));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G860), .ZN(G148));
  NOR2_X1   g177(.A1(new_n535), .A2(G868), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(KEYINPUT85), .A3(new_n601), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT85), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n593), .B2(G559), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n603), .B1(new_n607), .B2(G868), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT86), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT87), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g186(.A1(new_n464), .A2(new_n468), .A3(new_n467), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n477), .A2(G123), .ZN(new_n616));
  INV_X1    g191(.A(new_n473), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G135), .ZN(new_n618));
  NOR2_X1   g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n616), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2435), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2438), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(G1341), .B(G1348), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT88), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n632), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2072), .B(G2078), .Z(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n640), .B1(new_n644), .B2(KEYINPUT18), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2096), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n642), .A2(new_n643), .ZN(new_n649));
  AOI21_X1  g224(.A(KEYINPUT18), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n647), .B(new_n650), .Z(G227));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT89), .ZN(new_n653));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n653), .A2(new_n654), .ZN(new_n660));
  AOI22_X1  g235(.A1(new_n658), .A2(new_n659), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  OR3_X1    g236(.A1(new_n655), .A2(new_n660), .A3(new_n657), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n661), .B(new_n662), .C1(new_n659), .C2(new_n658), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT90), .B(KEYINPUT91), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1991), .B(G1996), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT21), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT22), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n668), .B(new_n670), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G229));
  MUX2_X1   g247(.A(G6), .B(G305), .S(G16), .Z(new_n673));
  XOR2_X1   g248(.A(KEYINPUT32), .B(G1981), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G22), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G166), .B2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(KEYINPUT94), .B1(G16), .B2(G23), .ZN(new_n681));
  OR3_X1    g256(.A1(KEYINPUT94), .A2(G16), .A3(G23), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n681), .B(new_n682), .C1(G288), .C2(new_n676), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT95), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT33), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n675), .A2(new_n680), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT34), .Z(new_n688));
  NOR2_X1   g263(.A1(G25), .A2(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n477), .A2(G119), .ZN(new_n690));
  OR2_X1    g265(.A1(G95), .A2(G2105), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n691), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G131), .ZN(new_n694));
  OAI21_X1  g269(.A(KEYINPUT92), .B1(new_n473), .B2(new_n694), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n473), .A2(KEYINPUT92), .A3(new_n694), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n689), .B1(new_n698), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT93), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT35), .B(G1991), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G16), .A2(G24), .ZN(new_n704));
  INV_X1    g279(.A(G290), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n688), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT36), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT103), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n676), .A2(G20), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n550), .A2(new_n552), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT77), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n550), .A2(KEYINPUT77), .A3(new_n552), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n547), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n714), .B1(new_n719), .B2(new_n676), .ZN(new_n720));
  INV_X1    g295(.A(G1956), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g297(.A(G1956), .B(new_n714), .C1(new_n719), .C2(new_n676), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n617), .A2(G139), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(new_n467), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT25), .Z(new_n729));
  NAND3_X1  g304(.A1(new_n725), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(KEYINPUT99), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT99), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n725), .A2(new_n727), .A3(new_n732), .A4(new_n729), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n731), .A2(G29), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G2072), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT100), .Z(new_n739));
  AOI21_X1  g314(.A(new_n735), .B1(new_n734), .B2(new_n737), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n477), .A2(G129), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n617), .A2(G141), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n464), .A2(G105), .A3(new_n467), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT26), .Z(new_n745));
  NAND4_X1  g320(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G32), .B(new_n746), .S(G29), .Z(new_n747));
  XOR2_X1   g322(.A(KEYINPUT27), .B(G1996), .Z(new_n748));
  AOI21_X1  g323(.A(new_n740), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT30), .B(G28), .Z(new_n750));
  MUX2_X1   g325(.A(new_n750), .B(new_n621), .S(G29), .Z(new_n751));
  NAND4_X1  g326(.A1(new_n724), .A2(new_n739), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G21), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G168), .B2(G16), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(G171), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G5), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1961), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n736), .A2(G27), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G164), .B2(new_n736), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n755), .B(new_n759), .C1(G2078), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(G2078), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n754), .A2(G1966), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n752), .A2(new_n762), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT31), .B(G11), .ZN(new_n767));
  INV_X1    g342(.A(G34), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(KEYINPUT24), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(KEYINPUT24), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  MUX2_X1   g346(.A(new_n771), .B(G160), .S(G29), .Z(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n757), .A2(new_n758), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n747), .A2(new_n748), .B1(new_n773), .B2(new_n772), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n766), .A2(new_n767), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT101), .B1(new_n779), .B2(G29), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n779), .A2(KEYINPUT101), .A3(G29), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n780), .B(new_n781), .C1(G162), .C2(new_n736), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT29), .B(G2090), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n593), .A2(G16), .ZN(new_n786));
  INV_X1    g361(.A(G4), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT96), .B(G1348), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n676), .A2(G19), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n535), .B2(new_n676), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1341), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n736), .A2(G26), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT97), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n477), .A2(G128), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n617), .A2(G140), .ZN(new_n799));
  OR2_X1    g374(.A1(G104), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n736), .ZN(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n786), .B(new_n789), .C1(new_n787), .C2(G16), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n791), .A2(new_n794), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT98), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n711), .B1(new_n785), .B2(new_n810), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n778), .A2(new_n809), .A3(new_n784), .A4(KEYINPUT103), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n710), .B1(new_n811), .B2(new_n812), .ZN(G150));
  INV_X1    g388(.A(KEYINPUT104), .ZN(new_n814));
  NAND2_X1  g389(.A1(G150), .A2(new_n814), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n710), .B(KEYINPUT104), .C1(new_n811), .C2(new_n812), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(G311));
  NAND2_X1  g392(.A1(G80), .A2(G543), .ZN(new_n818));
  INV_X1    g393(.A(G67), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n508), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n517), .A2(G55), .B1(new_n504), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n523), .A2(G93), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n535), .A2(new_n823), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n533), .A2(new_n534), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n827), .A2(new_n822), .A3(new_n821), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n593), .A2(new_n601), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n825), .B1(new_n833), .B2(G860), .ZN(G145));
  INV_X1    g409(.A(KEYINPUT106), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n731), .A2(new_n733), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n494), .A2(new_n468), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n839), .A2(new_n485), .A3(new_n488), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n746), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n802), .ZN(new_n842));
  MUX2_X1   g417(.A(new_n836), .B(new_n730), .S(new_n842), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n697), .B(new_n613), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n847), .B(new_n848), .C1(G118), .C2(new_n467), .ZN(new_n849));
  INV_X1    g424(.A(G142), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n473), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G130), .B2(new_n477), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n844), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n843), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n621), .B(G160), .Z(new_n856));
  XNOR2_X1  g431(.A(G162), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n835), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(G37), .B1(new_n855), .B2(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n854), .A2(KEYINPUT106), .A3(new_n857), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g438(.A(new_n607), .B(new_n829), .ZN(new_n864));
  INV_X1    g439(.A(new_n589), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n719), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(G299), .A2(new_n589), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(KEYINPUT41), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(KEYINPUT41), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n864), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n868), .B(KEYINPUT107), .Z(new_n874));
  AOI22_X1  g449(.A1(new_n872), .A2(KEYINPUT108), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n873), .A2(KEYINPUT108), .A3(new_n874), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT42), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G166), .B(G288), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G305), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n705), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n873), .A2(KEYINPUT108), .A3(new_n874), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n873), .A2(new_n874), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT108), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n864), .B2(new_n871), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n877), .A2(new_n880), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n880), .B1(new_n877), .B2(new_n886), .ZN(new_n888));
  OAI21_X1  g463(.A(G868), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n823), .A2(new_n574), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(G295));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n890), .ZN(G331));
  NAND3_X1  g467(.A1(new_n826), .A2(new_n828), .A3(G301), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(G301), .B1(new_n826), .B2(new_n828), .ZN(new_n895));
  OAI21_X1  g470(.A(G286), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(G168), .A3(new_n893), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n871), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n896), .A2(new_n898), .A3(new_n867), .A4(new_n866), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n880), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT109), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n869), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n870), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n868), .A2(new_n905), .A3(KEYINPUT41), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n899), .A3(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n874), .A2(new_n899), .ZN(new_n910));
  INV_X1    g485(.A(new_n880), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n904), .A2(KEYINPUT43), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n902), .A2(new_n903), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n880), .B1(new_n900), .B2(new_n901), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT44), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT110), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n914), .B1(new_n921), .B2(new_n915), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  INV_X1    g498(.A(new_n916), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n904), .A2(KEYINPUT43), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n919), .A2(new_n920), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n920), .B1(new_n919), .B2(new_n926), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(G397));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n485), .A2(new_n488), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n495), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(G160), .A2(G40), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n802), .B(G2067), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT111), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n746), .B(G1996), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n702), .A3(new_n698), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n803), .A2(new_n805), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n936), .B1(new_n940), .B2(new_n746), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n937), .B2(G1996), .ZN(new_n948));
  OR3_X1    g523(.A1(new_n937), .A2(new_n947), .A3(G1996), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  NAND2_X1  g526(.A1(new_n697), .A2(new_n701), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n698), .A2(new_n702), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n942), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n936), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n705), .A2(new_n707), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(new_n937), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT48), .Z(new_n958));
  AOI211_X1 g533(.A(new_n945), .B(new_n951), .C1(new_n955), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT126), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT57), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n715), .A2(new_n961), .A3(new_n548), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(G299), .B2(KEYINPUT57), .ZN(new_n964));
  OAI211_X1 g539(.A(KEYINPUT45), .B(new_n930), .C1(new_n495), .C2(new_n931), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n931), .A2(KEYINPUT72), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n839), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT45), .B1(new_n969), .B2(new_n930), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(G160), .A2(G40), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n489), .A2(new_n496), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n974), .B2(new_n839), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT112), .B1(new_n975), .B2(KEYINPUT45), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT56), .B(G2072), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n972), .A2(new_n973), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n969), .A2(new_n979), .A3(new_n930), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n932), .A2(KEYINPUT50), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n973), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n721), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n964), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n978), .A2(new_n964), .A3(new_n983), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n935), .A2(new_n932), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(G2067), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n969), .A2(new_n930), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n979), .B(new_n930), .C1(new_n495), .C2(new_n931), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n973), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1348), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n985), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n984), .B1(new_n996), .B2(new_n600), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n978), .A2(new_n983), .ZN(new_n998));
  INV_X1    g573(.A(new_n964), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n978), .A2(new_n964), .A3(new_n983), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(KEYINPUT61), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT117), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1000), .A2(new_n1004), .A3(KEYINPUT61), .A4(new_n1001), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n591), .A2(new_n1007), .A3(new_n592), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(new_n995), .A3(KEYINPUT60), .A4(new_n989), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT60), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n979), .B1(new_n969), .B2(new_n930), .ZN(new_n1012));
  INV_X1    g587(.A(new_n992), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1012), .A2(new_n935), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(G1348), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1011), .B1(new_n1015), .B2(new_n988), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1015), .A2(new_n1011), .A3(new_n988), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n593), .A2(KEYINPUT118), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1008), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1010), .B(new_n1016), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT61), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n985), .B2(new_n984), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT58), .B(G1341), .Z(new_n1024));
  NAND2_X1  g599(.A1(new_n987), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n971), .B(new_n933), .C1(G164), .C2(G1384), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n976), .A2(new_n973), .A3(new_n1026), .A4(new_n965), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT116), .B(G1996), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1023), .B1(new_n1029), .B2(new_n535), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1029), .A2(new_n1023), .A3(new_n535), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1020), .B(new_n1022), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n997), .B1(new_n1006), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT119), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1026), .A2(new_n965), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n973), .B1(new_n970), .B2(new_n971), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n679), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n982), .A2(G2090), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1035), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G303), .A2(G8), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1042), .B(KEYINPUT55), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT113), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G2090), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1014), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1035), .B1(new_n1038), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1044), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT49), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n565), .A2(new_n1051), .A3(new_n566), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n565), .B2(new_n566), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1050), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT49), .A3(new_n1052), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n986), .A2(new_n1035), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n987), .B(G8), .C1(new_n1060), .C2(G288), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT52), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1058), .B(new_n1063), .C1(new_n1060), .C2(G288), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1059), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1039), .B1(new_n1027), .B2(new_n679), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1066), .B(new_n1043), .C1(new_n1067), .C2(new_n1035), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1045), .A2(new_n1049), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1027), .B2(G2078), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n993), .A2(new_n758), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n973), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G2078), .B1(new_n935), .B2(KEYINPUT123), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n965), .A3(new_n934), .A4(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1071), .A2(G301), .A3(new_n1072), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n935), .B1(new_n933), .B2(new_n932), .ZN(new_n1080));
  INV_X1    g655(.A(G2078), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n969), .A2(KEYINPUT45), .A3(new_n930), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1080), .A2(KEYINPUT122), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(KEYINPUT53), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1071), .A2(new_n1072), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1079), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1069), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1071), .A2(new_n1072), .A3(new_n1076), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1071), .A2(new_n1087), .A3(G301), .A4(new_n1072), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(KEYINPUT54), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT125), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT125), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1095), .A2(new_n1099), .A3(KEYINPUT54), .A4(new_n1096), .ZN(new_n1100));
  NOR4_X1   g675(.A1(new_n1012), .A2(new_n1013), .A3(G2084), .A4(new_n935), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1966), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1102));
  OAI21_X1  g677(.A(G8), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G286), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(KEYINPUT120), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G286), .A2(G8), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1103), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1966), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1082), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n934), .A2(new_n973), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n991), .A2(new_n773), .A3(new_n973), .A4(new_n992), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(G8), .B(new_n1107), .C1(new_n1116), .C2(G286), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1106), .A2(KEYINPUT120), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1110), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1098), .A2(new_n1100), .B1(new_n1105), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1121), .B(new_n997), .C1(new_n1006), .C2(new_n1032), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1034), .A2(new_n1093), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1104), .A2(new_n1125), .A3(G168), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT114), .B1(new_n1103), .B2(G286), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1124), .B1(new_n1069), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1065), .B1(new_n1048), .B2(new_n1044), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1065), .B(KEYINPUT115), .C1(new_n1048), .C2(new_n1044), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1132), .A2(new_n1049), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1049), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1052), .B1(new_n1138), .B2(G288), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1137), .A2(new_n1065), .B1(new_n1058), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1069), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1119), .A2(new_n1105), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT62), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1119), .A2(new_n1144), .A3(new_n1105), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1089), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1136), .A2(new_n1140), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1123), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n954), .B1(G1986), .B2(G290), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n937), .B1(new_n1150), .B2(new_n956), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n960), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g728(.A(KEYINPUT126), .B(new_n1151), .C1(new_n1123), .C2(new_n1148), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n959), .B1(new_n1153), .B2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g730(.A(G227), .ZN(new_n1157));
  NAND3_X1  g731(.A1(new_n638), .A2(new_n456), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g732(.A(new_n1158), .B(KEYINPUT127), .Z(new_n1159));
  NOR2_X1   g733(.A1(new_n1159), .A2(G229), .ZN(new_n1160));
  NAND4_X1  g734(.A1(new_n1160), .A2(new_n862), .A3(new_n922), .A4(new_n925), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


