//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G141gat), .B(G148gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(new_n207), .B2(KEYINPUT2), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT78), .A2(G155gat), .A3(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT78), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT80), .B(G155gat), .Z(new_n219));
  OAI21_X1  g018(.A(KEYINPUT2), .B1(new_n219), .B2(new_n213), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n209), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n206), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT29), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT85), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT72), .B(G197gat), .Z(new_n229));
  INV_X1    g028(.A(G204gat), .ZN(new_n230));
  INV_X1    g029(.A(G211gat), .ZN(new_n231));
  INV_X1    g030(.A(G218gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI22_X1  g032(.A1(new_n229), .A2(new_n230), .B1(KEYINPUT22), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(new_n230), .B2(new_n229), .ZN(new_n235));
  XOR2_X1   g034(.A(G211gat), .B(G218gat), .Z(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n237), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n227), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n228), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT29), .B1(new_n238), .B2(new_n239), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n223), .B1(new_n244), .B2(KEYINPUT3), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n205), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n205), .B1(new_n226), .B2(new_n240), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(G22gat), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  INV_X1    g050(.A(G22gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n242), .A2(new_n241), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n226), .A2(new_n227), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n245), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(new_n204), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT31), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G50gat), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n250), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n250), .B2(new_n257), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G15gat), .B(G43gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(G71gat), .B(G99gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  NOR3_X1   g068(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT26), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR4_X1   g071(.A1(KEYINPUT66), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT67), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n276), .B(new_n268), .C1(new_n272), .C2(new_n273), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  AND2_X1   g077(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n281), .B(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n275), .A2(new_n277), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G183gat), .B(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(KEYINPUT24), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G169gat), .ZN(new_n290));
  INV_X1    g089(.A(G176gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT23), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n294), .A3(new_n269), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(G183gat), .A3(G190gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(new_n287), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n289), .A2(new_n296), .A3(KEYINPUT25), .A4(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n286), .B2(new_n297), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(new_n295), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309));
  INV_X1    g108(.A(G113gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G120gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(G120gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n313), .B1(KEYINPUT69), .B2(new_n311), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(KEYINPUT69), .B2(new_n311), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(new_n309), .A3(new_n306), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n305), .B(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G227gat), .A2(G233gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(KEYINPUT70), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT33), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(KEYINPUT32), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n267), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n320), .A2(new_n321), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT34), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT32), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n266), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n327), .B1(new_n266), .B2(new_n336), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n326), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n331), .A2(new_n334), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n333), .B1(new_n343), .B2(new_n330), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n263), .A2(new_n345), .A3(KEYINPUT87), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT35), .ZN(new_n347));
  XOR2_X1   g146(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n348));
  XNOR2_X1  g147(.A(G1gat), .B(G29gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G57gat), .B(G85gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  NAND2_X1  g151(.A1(new_n223), .A2(KEYINPUT3), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n319), .B1(new_n223), .B2(KEYINPUT3), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT81), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n224), .A2(new_n225), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT81), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n353), .A4(new_n319), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n319), .A2(new_n223), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n319), .A2(new_n223), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n361), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n365), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n369), .B(KEYINPUT84), .C1(new_n363), .C2(new_n362), .ZN(new_n370));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(KEYINPUT5), .ZN(new_n373));
  AND4_X1   g172(.A1(new_n360), .A2(new_n367), .A3(new_n370), .A4(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n319), .A2(new_n223), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n372), .B1(new_n375), .B2(new_n362), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n362), .A2(new_n365), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n319), .A2(new_n223), .A3(new_n363), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n378), .A2(new_n372), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n377), .B1(new_n360), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n352), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n352), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n360), .A2(new_n367), .A3(new_n370), .A4(new_n373), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n380), .A2(new_n360), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n383), .B(new_n384), .C1(new_n385), .C2(new_n377), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(KEYINPUT6), .B(new_n352), .C1(new_n374), .C2(new_n381), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n305), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n285), .A2(new_n396), .A3(new_n304), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n396), .B1(new_n285), .B2(new_n304), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n397), .A2(new_n398), .A3(new_n391), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n395), .B1(new_n399), .B2(KEYINPUT74), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n305), .A2(KEYINPUT73), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n285), .A2(new_n396), .A3(new_n304), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT74), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(KEYINPUT75), .B(new_n241), .C1(new_n400), .C2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n394), .B1(new_n403), .B2(new_n404), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n399), .A2(KEYINPUT74), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n240), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT75), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n392), .A2(KEYINPUT29), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n401), .A2(new_n402), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n285), .A2(new_n392), .A3(new_n304), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n418), .B2(new_n240), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n406), .B(new_n410), .C1(new_n413), .C2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT30), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n413), .A2(new_n419), .ZN(new_n426));
  AOI211_X1 g225(.A(new_n414), .B(new_n240), .C1(new_n411), .C2(new_n412), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT76), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT76), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n406), .B(new_n429), .C1(new_n413), .C2(new_n419), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n409), .A3(new_n430), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n423), .A2(new_n425), .A3(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n346), .A2(new_n347), .A3(new_n390), .A4(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n345), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n261), .A2(new_n262), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n423), .A2(new_n431), .A3(new_n390), .A4(new_n425), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT35), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n436), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n360), .A2(new_n367), .A3(new_n370), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n372), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n443), .A2(KEYINPUT39), .ZN(new_n444));
  OR3_X1    g243(.A1(new_n375), .A2(new_n362), .A3(new_n372), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(KEYINPUT39), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n383), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT40), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n444), .A2(KEYINPUT40), .A3(new_n383), .A4(new_n446), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n382), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT38), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n420), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n428), .A2(KEYINPUT37), .A3(new_n430), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n406), .B(new_n455), .C1(new_n413), .C2(new_n419), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n456), .A2(new_n409), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n453), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n388), .A2(new_n389), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n409), .A2(new_n452), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n416), .A2(new_n241), .A3(new_n417), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT86), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n411), .A2(new_n240), .A3(new_n412), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n462), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n460), .B1(new_n466), .B2(KEYINPUT37), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n456), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  OAI22_X1  g268(.A1(new_n432), .A2(new_n451), .B1(new_n458), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n441), .B1(new_n470), .B2(new_n436), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT36), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT36), .B1(new_n342), .B2(new_n344), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n440), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G113gat), .B(G141gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(G197gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT11), .B(G169gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n479), .B(KEYINPUT12), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G50gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G43gat), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT15), .B1(new_n483), .B2(KEYINPUT88), .ZN(new_n484));
  INV_X1    g283(.A(G43gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(G50gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n484), .B(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(G29gat), .A2(G36gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n489), .B(KEYINPUT14), .Z(new_n490));
  NAND2_X1  g289(.A1(G29gat), .A2(G36gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT89), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  AOI211_X1 g294(.A(new_n495), .B(new_n487), .C1(new_n490), .C2(new_n491), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n498), .A2(G1gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT16), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n500), .B2(G1gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G8gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n499), .B(new_n501), .C1(new_n503), .C2(G8gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n497), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n497), .A2(KEYINPUT17), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT91), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n497), .A2(KEYINPUT17), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n512), .A2(new_n508), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT18), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n497), .B(new_n508), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n515), .B(KEYINPUT13), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n518), .B1(new_n514), .B2(new_n515), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n481), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n525), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n527), .A2(new_n523), .A3(new_n519), .A4(new_n480), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT7), .ZN(new_n534));
  OAI211_X1 g333(.A(G85gat), .B(G92gat), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT97), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(KEYINPUT96), .B2(KEYINPUT7), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n535), .B(KEYINPUT97), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n539), .A2(new_n533), .A3(new_n534), .ZN(new_n540));
  NOR2_X1   g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n542), .A2(KEYINPUT98), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT8), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n542), .B2(KEYINPUT98), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n541), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n538), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G99gat), .B(G106gat), .Z(new_n548));
  OR2_X1    g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(G57gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G64gat), .ZN(new_n554));
  AND2_X1   g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(KEYINPUT9), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n559));
  AND2_X1   g358(.A1(G57gat), .A2(G64gat), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n555), .A2(new_n556), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n554), .A2(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n551), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT10), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n567), .A2(new_n566), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT99), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n532), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT99), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n531), .B1(new_n565), .B2(new_n567), .ZN(new_n575));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT100), .ZN(new_n577));
  XNOR2_X1  g376(.A(G120gat), .B(G148gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n532), .B1(new_n568), .B2(new_n569), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n580), .B1(new_n583), .B2(new_n575), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n530), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT21), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n564), .B1(new_n508), .B2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n508), .A2(new_n587), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n590), .A2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n593), .B2(new_n594), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G183gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G211gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT94), .B(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G134gat), .B(G162gat), .Z(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n511), .A2(new_n512), .A3(new_n551), .ZN(new_n612));
  INV_X1    g411(.A(new_n551), .ZN(new_n613));
  INV_X1    g412(.A(new_n497), .ZN(new_n614));
  AND2_X1   g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n613), .A2(new_n614), .B1(KEYINPUT41), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n611), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n615), .A2(KEYINPUT41), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n612), .A2(new_n616), .A3(new_n611), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  INV_X1    g423(.A(new_n622), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n624), .B1(new_n625), .B2(new_n617), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  AND4_X1   g426(.A1(new_n475), .A2(new_n586), .A3(new_n609), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n459), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g429(.A1(new_n423), .A2(new_n431), .A3(new_n425), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT42), .B1(new_n632), .B2(new_n505), .ZN(new_n633));
  NAND2_X1  g432(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n500), .A2(new_n505), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  MUX2_X1   g435(.A(KEYINPUT42), .B(new_n633), .S(new_n636), .Z(G1325gat));
  AOI21_X1  g436(.A(G15gat), .B1(new_n628), .B2(new_n434), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT101), .B1(new_n472), .B2(new_n473), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n345), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n342), .A2(new_n344), .A3(KEYINPUT36), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT102), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n639), .A2(new_n644), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n650), .A2(G15gat), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n638), .B1(new_n628), .B2(new_n651), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n628), .A2(new_n263), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT103), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT43), .B(G22gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  AND2_X1   g455(.A1(new_n623), .A2(new_n626), .ZN(new_n657));
  INV_X1    g456(.A(new_n609), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n586), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n475), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G29gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n662), .A3(new_n459), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT45), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  INV_X1    g464(.A(new_n440), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n471), .B2(new_n645), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n390), .B1(new_n456), .B2(new_n467), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n454), .A2(new_n457), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n669), .B1(new_n670), .B2(new_n453), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n631), .A2(new_n382), .A3(new_n450), .A4(new_n449), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n263), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(KEYINPUT104), .B(new_n647), .C1(new_n673), .C2(new_n441), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n666), .B1(new_n668), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n665), .B1(new_n675), .B2(new_n627), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n475), .A2(KEYINPUT44), .A3(new_n657), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(new_n390), .A3(new_n659), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n664), .B1(new_n679), .B2(new_n662), .ZN(G1328gat));
  NAND4_X1  g479(.A1(new_n676), .A2(new_n631), .A3(new_n660), .A4(new_n677), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G36gat), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n432), .A2(G36gat), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n475), .A2(new_n657), .A3(new_n660), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT46), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT105), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n682), .B(new_n686), .C1(KEYINPUT46), .C2(new_n684), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT106), .ZN(G1329gat));
  NAND3_X1  g487(.A1(new_n661), .A2(new_n485), .A3(new_n434), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT107), .Z(new_n690));
  NAND4_X1  g489(.A1(new_n676), .A2(new_n645), .A3(new_n660), .A4(new_n677), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n692));
  OAI21_X1  g491(.A(G43gat), .B1(new_n691), .B2(KEYINPUT108), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n690), .B(KEYINPUT47), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n676), .A2(new_n677), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n650), .A3(new_n660), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G43gat), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n697), .A2(new_n690), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n694), .B1(new_n698), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g498(.A1(new_n661), .A2(new_n482), .A3(new_n263), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n678), .A2(new_n436), .A3(new_n659), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n482), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1331gat));
  INV_X1    g503(.A(new_n585), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n609), .A2(new_n627), .ZN(new_n706));
  NOR4_X1   g505(.A1(new_n675), .A2(new_n529), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n459), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n631), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT49), .B(G64gat), .Z(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n710), .B2(new_n712), .ZN(G1333gat));
  NAND2_X1  g512(.A1(new_n707), .A2(new_n650), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n345), .A2(G71gat), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n714), .A2(G71gat), .B1(new_n707), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g516(.A1(new_n707), .A2(new_n263), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g518(.A1(new_n668), .A2(new_n674), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n627), .B1(new_n720), .B2(new_n440), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n609), .A2(new_n529), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT51), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724));
  INV_X1    g523(.A(new_n722), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n675), .A2(new_n724), .A3(new_n627), .A4(new_n725), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n723), .A2(new_n726), .A3(KEYINPUT110), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(KEYINPUT110), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n705), .A2(G85gat), .A3(new_n390), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n722), .A2(new_n585), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(KEYINPUT109), .Z(new_n732));
  AND3_X1   g531(.A1(new_n676), .A2(new_n677), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734), .B2(new_n390), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n730), .A2(new_n735), .ZN(G1336gat));
  NOR2_X1   g535(.A1(new_n723), .A2(new_n726), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n432), .A2(new_n705), .A3(G92gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(G92gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n733), .B2(new_n631), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT52), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n742), .A2(KEYINPUT52), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n727), .A2(new_n728), .A3(new_n738), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(G1337gat));
  XOR2_X1   g545(.A(KEYINPUT111), .B(G99gat), .Z(new_n747));
  NOR3_X1   g546(.A1(new_n705), .A2(new_n345), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n727), .A2(new_n728), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n650), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n747), .B1(new_n734), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1338gat));
  NOR3_X1   g551(.A1(new_n705), .A2(G106gat), .A3(new_n436), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT113), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n723), .B2(new_n726), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n676), .A2(new_n263), .A3(new_n677), .A4(new_n732), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G106gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT112), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n761), .A3(G106gat), .ZN(new_n762));
  OAI211_X1 g561(.A(KEYINPUT114), .B(new_n754), .C1(new_n723), .C2(new_n726), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n757), .A2(new_n760), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT53), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n727), .A2(new_n728), .A3(new_n753), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n767), .A3(new_n759), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770));
  OAI21_X1  g569(.A(KEYINPUT54), .B1(new_n570), .B2(new_n531), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n572), .B2(new_n573), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n773));
  AOI21_X1  g572(.A(new_n579), .B1(new_n583), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n573), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT99), .B1(new_n568), .B2(new_n569), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n777), .A2(new_n778), .A3(new_n532), .ZN(new_n779));
  OAI211_X1 g578(.A(KEYINPUT55), .B(new_n774), .C1(new_n779), .C2(new_n771), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n776), .A2(new_n780), .A3(new_n529), .A4(new_n582), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n514), .A2(new_n515), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n521), .A2(new_n522), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n479), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n524), .A2(new_n525), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n480), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n657), .B1(new_n585), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n776), .A2(new_n786), .A3(new_n780), .A4(new_n582), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n657), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n790), .A3(new_n658), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n705), .A2(new_n530), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n706), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n432), .A2(new_n459), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n434), .A2(new_n436), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n530), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(new_n310), .ZN(G1340gat));
  NOR2_X1   g600(.A1(new_n799), .A2(new_n705), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g602(.A1(new_n799), .A2(new_n658), .ZN(new_n804));
  XOR2_X1   g603(.A(KEYINPUT116), .B(G127gat), .Z(new_n805));
  XNOR2_X1  g604(.A(new_n804), .B(new_n805), .ZN(G1342gat));
  NAND3_X1  g605(.A1(new_n795), .A2(new_n657), .A3(new_n798), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(G134gat), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(G134gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(G1343gat));
  NOR2_X1   g612(.A1(new_n650), .A2(new_n796), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n609), .B1(new_n781), .B2(new_n787), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n793), .B1(new_n815), .B2(new_n790), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n436), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n818), .A2(G141gat), .A3(new_n530), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n819), .B(new_n820), .ZN(new_n821));
  XOR2_X1   g620(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n822));
  NOR2_X1   g621(.A1(new_n645), .A2(new_n796), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT57), .B1(new_n795), .B2(new_n263), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n816), .A2(new_n825), .A3(new_n436), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n530), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(G141gat), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n821), .B(new_n822), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n827), .A2(KEYINPUT117), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n836), .B(new_n823), .C1(new_n824), .C2(new_n826), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n529), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n819), .B1(new_n839), .B2(G141gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n833), .B1(new_n834), .B2(new_n840), .ZN(G1344gat));
  OR3_X1    g640(.A1(new_n818), .A2(G148gat), .A3(new_n705), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n263), .B1(new_n816), .B2(KEYINPUT121), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845));
  AOI211_X1 g644(.A(new_n845), .B(new_n793), .C1(new_n815), .C2(new_n790), .ZN(new_n846));
  OAI211_X1 g645(.A(KEYINPUT122), .B(new_n825), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n826), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n795), .A2(new_n845), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n816), .A2(KEYINPUT121), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n851), .A3(new_n263), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT122), .B1(new_n852), .B2(new_n825), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n585), .B(new_n823), .C1(new_n849), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n843), .B1(new_n854), .B2(G148gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n843), .A2(G148gat), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n838), .B2(new_n585), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n842), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT123), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(new_n842), .C1(new_n855), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1345gat));
  NOR2_X1   g661(.A1(new_n658), .A2(new_n219), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n814), .A2(new_n609), .A3(new_n817), .ZN(new_n864));
  AOI22_X1  g663(.A1(new_n838), .A2(new_n863), .B1(new_n864), .B2(new_n219), .ZN(G1346gat));
  NOR3_X1   g664(.A1(new_n818), .A2(G162gat), .A3(new_n627), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT124), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n627), .B1(new_n835), .B2(new_n837), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n213), .B2(new_n868), .ZN(G1347gat));
  NOR3_X1   g668(.A1(new_n797), .A2(new_n432), .A3(new_n459), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n795), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n530), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(new_n290), .ZN(G1348gat));
  NOR2_X1   g672(.A1(new_n871), .A2(new_n705), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(new_n291), .ZN(G1349gat));
  NOR2_X1   g674(.A1(new_n871), .A2(new_n658), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n280), .B2(new_n279), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT125), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(KEYINPUT125), .ZN(new_n879));
  INV_X1    g678(.A(new_n876), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT126), .B1(new_n880), .B2(G183gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g682(.A1(new_n871), .A2(new_n627), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n278), .ZN(new_n886));
  XOR2_X1   g685(.A(KEYINPUT61), .B(G190gat), .Z(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n884), .B2(new_n887), .ZN(G1351gat));
  INV_X1    g687(.A(G197gat), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n849), .A2(new_n853), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n650), .A2(new_n459), .A3(new_n432), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n892), .B2(new_n529), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n817), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(G197gat), .A3(new_n530), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n893), .A2(new_n895), .ZN(G1352gat));
  NOR3_X1   g695(.A1(new_n894), .A2(G204gat), .A3(new_n705), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT62), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n585), .A3(new_n891), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n900), .B2(new_n230), .ZN(G1353gat));
  NAND3_X1  g700(.A1(new_n890), .A2(new_n609), .A3(new_n891), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n902), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT63), .B1(new_n902), .B2(G211gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n609), .A2(new_n231), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n903), .A2(new_n904), .B1(new_n894), .B2(new_n905), .ZN(G1354gat));
  OAI21_X1  g705(.A(new_n232), .B1(new_n894), .B2(new_n627), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT127), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n627), .A2(new_n232), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n892), .B2(new_n909), .ZN(G1355gat));
endmodule


