

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585;

  AND2_X2 U320 ( .A1(n508), .A2(n543), .ZN(n509) );
  XNOR2_X2 U321 ( .A(G99GAT), .B(G106GAT), .ZN(n369) );
  XNOR2_X1 U322 ( .A(n479), .B(KEYINPUT64), .ZN(n504) );
  XNOR2_X2 U323 ( .A(n289), .B(n369), .ZN(n413) );
  XOR2_X2 U324 ( .A(G85GAT), .B(G92GAT), .Z(n289) );
  XNOR2_X2 U325 ( .A(n430), .B(n429), .ZN(n478) );
  XNOR2_X1 U326 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U327 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n288) );
  INV_X1 U328 ( .A(KEYINPUT65), .ZN(n370) );
  XNOR2_X1 U329 ( .A(n371), .B(n370), .ZN(n372) );
  NAND2_X1 U330 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U331 ( .A(n413), .B(n372), .ZN(n373) );
  XNOR2_X1 U332 ( .A(n428), .B(n427), .ZN(n429) );
  NOR2_X1 U333 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U334 ( .A(n458), .B(n457), .ZN(n583) );
  XNOR2_X1 U335 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U336 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n291) );
  XNOR2_X1 U337 ( .A(G1GAT), .B(G57GAT), .ZN(n290) );
  XNOR2_X1 U338 ( .A(n291), .B(n290), .ZN(n309) );
  XOR2_X1 U339 ( .A(G148GAT), .B(G162GAT), .Z(n293) );
  XNOR2_X1 U340 ( .A(G141GAT), .B(G120GAT), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n295) );
  XOR2_X1 U342 ( .A(G29GAT), .B(G85GAT), .Z(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n305) );
  XOR2_X1 U344 ( .A(G127GAT), .B(KEYINPUT0), .Z(n297) );
  XNOR2_X1 U345 ( .A(G113GAT), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n341) );
  XOR2_X1 U347 ( .A(G155GAT), .B(KEYINPUT2), .Z(n299) );
  XNOR2_X1 U348 ( .A(KEYINPUT93), .B(KEYINPUT3), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n327) );
  XNOR2_X1 U350 ( .A(n341), .B(n327), .ZN(n303) );
  XOR2_X1 U351 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n301) );
  XNOR2_X1 U352 ( .A(KEYINPUT97), .B(KEYINPUT4), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n307) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n465) );
  INV_X1 U359 ( .A(n465), .ZN(n567) );
  XOR2_X1 U360 ( .A(KEYINPUT23), .B(G106GAT), .Z(n311) );
  XNOR2_X1 U361 ( .A(G50GAT), .B(G218GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U363 ( .A(G204GAT), .B(KEYINPUT90), .Z(n313) );
  XNOR2_X1 U364 ( .A(KEYINPUT22), .B(KEYINPUT96), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U367 ( .A(G141GAT), .B(G22GAT), .Z(n439) );
  XOR2_X1 U368 ( .A(G148GAT), .B(G78GAT), .Z(n428) );
  XOR2_X1 U369 ( .A(KEYINPUT75), .B(G162GAT), .Z(n383) );
  XOR2_X1 U370 ( .A(n428), .B(n383), .Z(n317) );
  NAND2_X1 U371 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n439), .B(n318), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U375 ( .A(KEYINPUT91), .B(KEYINPUT95), .Z(n322) );
  XNOR2_X1 U376 ( .A(KEYINPUT94), .B(KEYINPUT24), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U378 ( .A(n324), .B(n323), .Z(n329) );
  XOR2_X1 U379 ( .A(G211GAT), .B(KEYINPUT21), .Z(n326) );
  XNOR2_X1 U380 ( .A(G197GAT), .B(KEYINPUT92), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n335) );
  XNOR2_X1 U382 ( .A(n327), .B(n335), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n548) );
  XOR2_X1 U384 ( .A(n548), .B(KEYINPUT28), .Z(n474) );
  XOR2_X1 U385 ( .A(G190GAT), .B(G218GAT), .Z(n382) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(G204GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n330), .B(G64GAT), .ZN(n424) );
  XOR2_X1 U388 ( .A(G183GAT), .B(KEYINPUT81), .Z(n389) );
  XOR2_X1 U389 ( .A(n424), .B(n389), .Z(n333) );
  XOR2_X1 U390 ( .A(G169GAT), .B(G8GAT), .Z(n436) );
  XNOR2_X1 U391 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n331), .B(KEYINPUT17), .ZN(n344) );
  XNOR2_X1 U393 ( .A(n436), .B(n344), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U395 ( .A(n334), .B(G92GAT), .Z(n337) );
  XNOR2_X1 U396 ( .A(G36GAT), .B(n335), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U398 ( .A(n382), .B(n338), .Z(n340) );
  NAND2_X1 U399 ( .A1(G226GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n545) );
  XNOR2_X1 U401 ( .A(n545), .B(KEYINPUT27), .ZN(n361) );
  NAND2_X1 U402 ( .A1(n465), .A2(n361), .ZN(n531) );
  NOR2_X1 U403 ( .A1(n474), .A2(n531), .ZN(n517) );
  XOR2_X1 U404 ( .A(G120GAT), .B(G71GAT), .Z(n419) );
  XOR2_X1 U405 ( .A(n419), .B(n341), .Z(n343) );
  NAND2_X1 U406 ( .A1(G227GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n345) );
  XOR2_X1 U408 ( .A(n345), .B(n344), .Z(n347) );
  XNOR2_X1 U409 ( .A(G169GAT), .B(G15GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n355) );
  XOR2_X1 U411 ( .A(KEYINPUT20), .B(G190GAT), .Z(n349) );
  XNOR2_X1 U412 ( .A(G43GAT), .B(G99GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U414 ( .A(G176GAT), .B(G183GAT), .Z(n351) );
  XNOR2_X1 U415 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U417 ( .A(n353), .B(n352), .Z(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n551) );
  NAND2_X1 U419 ( .A1(n517), .A2(n551), .ZN(n356) );
  XOR2_X1 U420 ( .A(KEYINPUT99), .B(n356), .Z(n366) );
  INV_X1 U421 ( .A(n551), .ZN(n471) );
  NAND2_X1 U422 ( .A1(n471), .A2(n545), .ZN(n357) );
  NAND2_X1 U423 ( .A1(n548), .A2(n357), .ZN(n358) );
  XOR2_X1 U424 ( .A(KEYINPUT25), .B(n358), .Z(n363) );
  XNOR2_X1 U425 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n360) );
  NOR2_X1 U426 ( .A1(n471), .A2(n548), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n568) );
  NAND2_X1 U428 ( .A1(n568), .A2(n361), .ZN(n362) );
  NAND2_X1 U429 ( .A1(n363), .A2(n362), .ZN(n364) );
  NAND2_X1 U430 ( .A1(n567), .A2(n364), .ZN(n365) );
  NAND2_X1 U431 ( .A1(n366), .A2(n365), .ZN(n459) );
  XOR2_X1 U432 ( .A(KEYINPUT79), .B(KEYINPUT11), .Z(n368) );
  XNOR2_X1 U433 ( .A(KEYINPUT9), .B(KEYINPUT76), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n374) );
  NAND2_X1 U435 ( .A1(G232GAT), .A2(G233GAT), .ZN(n371) );
  XOR2_X1 U436 ( .A(n374), .B(n373), .Z(n387) );
  XNOR2_X1 U437 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n375), .B(G29GAT), .ZN(n376) );
  XOR2_X1 U439 ( .A(n376), .B(KEYINPUT8), .Z(n378) );
  XNOR2_X1 U440 ( .A(G43GAT), .B(G50GAT), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n434) );
  XOR2_X1 U442 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n380) );
  XNOR2_X1 U443 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n434), .B(n381), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n384) );
  INV_X1 U447 ( .A(n388), .ZN(n543) );
  XOR2_X1 U448 ( .A(KEYINPUT80), .B(n543), .Z(n562) );
  INV_X1 U449 ( .A(n562), .ZN(n458) );
  XOR2_X1 U450 ( .A(n389), .B(G211GAT), .Z(n391) );
  XOR2_X1 U451 ( .A(G15GAT), .B(G1GAT), .Z(n435) );
  XNOR2_X1 U452 ( .A(n435), .B(G155GAT), .ZN(n390) );
  XNOR2_X1 U453 ( .A(n391), .B(n390), .ZN(n396) );
  XNOR2_X1 U454 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n392), .B(KEYINPUT72), .ZN(n423) );
  XOR2_X1 U456 ( .A(n423), .B(KEYINPUT15), .Z(n394) );
  NAND2_X1 U457 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U459 ( .A(n396), .B(n395), .Z(n398) );
  XNOR2_X1 U460 ( .A(G22GAT), .B(G78GAT), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U462 ( .A(G64GAT), .B(G127GAT), .Z(n400) );
  XNOR2_X1 U463 ( .A(G8GAT), .B(G71GAT), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U465 ( .A(n402), .B(n401), .Z(n410) );
  XOR2_X1 U466 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n404) );
  XNOR2_X1 U467 ( .A(KEYINPUT82), .B(KEYINPUT84), .ZN(n403) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U469 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n406) );
  XNOR2_X1 U470 ( .A(KEYINPUT86), .B(KEYINPUT12), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U472 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n578) );
  NAND2_X1 U474 ( .A1(n458), .A2(n578), .ZN(n411) );
  XOR2_X1 U475 ( .A(KEYINPUT16), .B(n411), .Z(n412) );
  AND2_X1 U476 ( .A1(n459), .A2(n412), .ZN(n480) );
  XNOR2_X1 U477 ( .A(n413), .B(KEYINPUT32), .ZN(n416) );
  INV_X1 U478 ( .A(n416), .ZN(n415) );
  INV_X1 U479 ( .A(KEYINPUT73), .ZN(n414) );
  NAND2_X1 U480 ( .A1(n415), .A2(n414), .ZN(n418) );
  NAND2_X1 U481 ( .A1(n416), .A2(KEYINPUT73), .ZN(n417) );
  NAND2_X1 U482 ( .A1(n418), .A2(n417), .ZN(n422) );
  XNOR2_X1 U483 ( .A(n419), .B(KEYINPUT31), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n420), .B(KEYINPUT33), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n430) );
  NAND2_X1 U488 ( .A1(G230GAT), .A2(G233GAT), .ZN(n427) );
  XOR2_X1 U489 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n432) );
  XNOR2_X1 U490 ( .A(KEYINPUT69), .B(KEYINPUT66), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n447) );
  XOR2_X1 U493 ( .A(G113GAT), .B(G197GAT), .Z(n438) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U496 ( .A(n440), .B(n439), .Z(n445) );
  XOR2_X1 U497 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n442) );
  NAND2_X1 U498 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U500 ( .A(KEYINPUT29), .B(n443), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n570) );
  XNOR2_X1 U503 ( .A(n570), .B(KEYINPUT71), .ZN(n554) );
  INV_X1 U504 ( .A(n554), .ZN(n512) );
  NOR2_X1 U505 ( .A1(n478), .A2(n512), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n448), .B(KEYINPUT74), .ZN(n462) );
  NAND2_X1 U507 ( .A1(n480), .A2(n462), .ZN(n454) );
  NOR2_X1 U508 ( .A1(n567), .A2(n454), .ZN(n449) );
  XOR2_X1 U509 ( .A(KEYINPUT34), .B(n449), .Z(n450) );
  XNOR2_X1 U510 ( .A(G1GAT), .B(n450), .ZN(G1324GAT) );
  INV_X1 U511 ( .A(n545), .ZN(n494) );
  NOR2_X1 U512 ( .A1(n494), .A2(n454), .ZN(n451) );
  XOR2_X1 U513 ( .A(G8GAT), .B(n451), .Z(G1325GAT) );
  NOR2_X1 U514 ( .A1(n551), .A2(n454), .ZN(n453) );
  XNOR2_X1 U515 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n452) );
  XNOR2_X1 U516 ( .A(n453), .B(n452), .ZN(G1326GAT) );
  INV_X1 U517 ( .A(n474), .ZN(n501) );
  NOR2_X1 U518 ( .A1(n501), .A2(n454), .ZN(n456) );
  XNOR2_X1 U519 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n455) );
  XNOR2_X1 U520 ( .A(n456), .B(n455), .ZN(G1327GAT) );
  XOR2_X1 U521 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n467) );
  XNOR2_X1 U522 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n457) );
  NOR2_X1 U523 ( .A1(n583), .A2(n578), .ZN(n460) );
  NAND2_X1 U524 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U525 ( .A(KEYINPUT37), .B(n461), .ZN(n492) );
  NAND2_X1 U526 ( .A1(n462), .A2(n492), .ZN(n463) );
  XNOR2_X1 U527 ( .A(n463), .B(KEYINPUT38), .ZN(n464) );
  XNOR2_X1 U528 ( .A(KEYINPUT103), .B(n464), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n475), .A2(n465), .ZN(n466) );
  XNOR2_X1 U530 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U531 ( .A(G29GAT), .B(n468), .ZN(G1328GAT) );
  XOR2_X1 U532 ( .A(G36GAT), .B(KEYINPUT105), .Z(n470) );
  NAND2_X1 U533 ( .A1(n545), .A2(n475), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(G1329GAT) );
  NAND2_X1 U535 ( .A1(n475), .A2(n471), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n472), .B(KEYINPUT40), .ZN(n473) );
  XNOR2_X1 U537 ( .A(G43GAT), .B(n473), .ZN(G1330GAT) );
  NAND2_X1 U538 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(KEYINPUT106), .ZN(n477) );
  XNOR2_X1 U540 ( .A(G50GAT), .B(n477), .ZN(G1331GAT) );
  XNOR2_X1 U541 ( .A(n478), .B(KEYINPUT41), .ZN(n479) );
  XOR2_X1 U542 ( .A(n504), .B(KEYINPUT108), .Z(n557) );
  AND2_X1 U543 ( .A1(n570), .A2(n557), .ZN(n491) );
  NAND2_X1 U544 ( .A1(n491), .A2(n480), .ZN(n488) );
  NOR2_X1 U545 ( .A1(n567), .A2(n488), .ZN(n485) );
  XOR2_X1 U546 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n482) );
  XNOR2_X1 U547 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n481) );
  XNOR2_X1 U548 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U549 ( .A(KEYINPUT107), .B(n483), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n485), .B(n484), .ZN(G1332GAT) );
  NOR2_X1 U551 ( .A1(n494), .A2(n488), .ZN(n486) );
  XOR2_X1 U552 ( .A(G64GAT), .B(n486), .Z(G1333GAT) );
  NOR2_X1 U553 ( .A1(n551), .A2(n488), .ZN(n487) );
  XOR2_X1 U554 ( .A(G71GAT), .B(n487), .Z(G1334GAT) );
  NOR2_X1 U555 ( .A1(n501), .A2(n488), .ZN(n490) );
  XNOR2_X1 U556 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n489) );
  XNOR2_X1 U557 ( .A(n490), .B(n489), .ZN(G1335GAT) );
  NAND2_X1 U558 ( .A1(n492), .A2(n491), .ZN(n500) );
  NOR2_X1 U559 ( .A1(n567), .A2(n500), .ZN(n493) );
  XOR2_X1 U560 ( .A(G85GAT), .B(n493), .Z(G1336GAT) );
  NOR2_X1 U561 ( .A1(n494), .A2(n500), .ZN(n495) );
  XOR2_X1 U562 ( .A(G92GAT), .B(n495), .Z(G1337GAT) );
  NOR2_X1 U563 ( .A1(n551), .A2(n500), .ZN(n497) );
  XNOR2_X1 U564 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n496) );
  XNOR2_X1 U565 ( .A(n497), .B(n496), .ZN(G1338GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n499) );
  XNOR2_X1 U567 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n498) );
  XNOR2_X1 U568 ( .A(n499), .B(n498), .ZN(n503) );
  NOR2_X1 U569 ( .A1(n501), .A2(n500), .ZN(n502) );
  XOR2_X1 U570 ( .A(n503), .B(n502), .Z(G1339GAT) );
  XNOR2_X1 U571 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n521) );
  NOR2_X1 U572 ( .A1(n570), .A2(n504), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n505), .B(KEYINPUT46), .ZN(n506) );
  NOR2_X2 U574 ( .A1(n506), .A2(n578), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n507), .B(KEYINPUT114), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(KEYINPUT47), .ZN(n515) );
  INV_X1 U577 ( .A(n578), .ZN(n539) );
  NOR2_X1 U578 ( .A1(n583), .A2(n539), .ZN(n510) );
  XOR2_X1 U579 ( .A(KEYINPUT45), .B(n510), .Z(n511) );
  NOR2_X1 U580 ( .A1(n478), .A2(n511), .ZN(n513) );
  NAND2_X1 U581 ( .A1(n513), .A2(n512), .ZN(n514) );
  NAND2_X1 U582 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X2 U583 ( .A(n516), .B(KEYINPUT48), .ZN(n546) );
  NAND2_X1 U584 ( .A1(n546), .A2(n517), .ZN(n518) );
  NOR2_X1 U585 ( .A1(n551), .A2(n518), .ZN(n519) );
  XOR2_X1 U586 ( .A(KEYINPUT115), .B(n519), .Z(n528) );
  NAND2_X1 U587 ( .A1(n528), .A2(n554), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n523) );
  NAND2_X1 U590 ( .A1(n528), .A2(n557), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U592 ( .A(G120GAT), .B(n524), .Z(G1341GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n526) );
  NAND2_X1 U594 ( .A1(n528), .A2(n578), .ZN(n525) );
  XNOR2_X1 U595 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U596 ( .A(G127GAT), .B(n527), .Z(G1342GAT) );
  XOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT51), .Z(n530) );
  NAND2_X1 U598 ( .A1(n528), .A2(n562), .ZN(n529) );
  XNOR2_X1 U599 ( .A(n530), .B(n529), .ZN(G1343GAT) );
  INV_X1 U600 ( .A(n568), .ZN(n532) );
  NOR2_X1 U601 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U602 ( .A1(n546), .A2(n533), .ZN(n542) );
  NOR2_X1 U603 ( .A1(n570), .A2(n542), .ZN(n535) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n534) );
  XNOR2_X1 U605 ( .A(n535), .B(n534), .ZN(G1344GAT) );
  NOR2_X1 U606 ( .A1(n504), .A2(n542), .ZN(n537) );
  XNOR2_X1 U607 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n536) );
  XNOR2_X1 U608 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(n538), .ZN(G1345GAT) );
  NOR2_X1 U610 ( .A1(n539), .A2(n542), .ZN(n540) );
  XOR2_X1 U611 ( .A(KEYINPUT120), .B(n540), .Z(n541) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(n541), .ZN(G1346GAT) );
  NOR2_X1 U613 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U614 ( .A(G162GAT), .B(n544), .Z(G1347GAT) );
  XOR2_X1 U615 ( .A(G169GAT), .B(KEYINPUT123), .Z(n556) );
  XNOR2_X1 U616 ( .A(n547), .B(n288), .ZN(n566) );
  AND2_X1 U617 ( .A1(n567), .A2(n548), .ZN(n549) );
  NAND2_X1 U618 ( .A1(n566), .A2(n549), .ZN(n550) );
  XOR2_X1 U619 ( .A(n550), .B(KEYINPUT55), .Z(n552) );
  XNOR2_X1 U620 ( .A(KEYINPUT122), .B(n553), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n563), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n559) );
  NAND2_X1 U624 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n578), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  AND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n582) );
  NOR2_X1 U634 ( .A1(n570), .A2(n582), .ZN(n575) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT59), .B(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U641 ( .A(n582), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n579), .A2(n478), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

