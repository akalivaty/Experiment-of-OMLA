//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  INV_X1    g000(.A(G101), .ZN(new_n187));
  INV_X1    g001(.A(G107), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G104), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G107), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n187), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT76), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT76), .ZN(new_n194));
  AOI211_X1 g008(.A(new_n194), .B(new_n187), .C1(new_n189), .C2(new_n191), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n188), .A3(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT3), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n197), .A2(new_n200), .A3(new_n188), .A4(G104), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n199), .A2(new_n187), .A3(new_n201), .A4(new_n191), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT2), .B(G113), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G116), .B(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(KEYINPUT5), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT5), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G116), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT80), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n212), .A2(new_n208), .A3(new_n209), .A4(G116), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(G113), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n196), .A2(new_n202), .A3(new_n206), .A4(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n199), .A2(new_n201), .A3(new_n191), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G101), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n217), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n219), .A3(G101), .ZN(new_n220));
  INV_X1    g034(.A(new_n205), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n203), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n206), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n215), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G110), .B(G122), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n215), .B(new_n226), .C1(new_n218), .C2(new_n224), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n228), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(KEYINPUT6), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n217), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n220), .A3(new_n223), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n226), .B1(new_n233), .B2(new_n215), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT6), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n225), .A2(new_n236), .A3(new_n227), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT81), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n230), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n245), .A2(new_n248), .A3(KEYINPUT64), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT64), .B1(new_n245), .B2(new_n248), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  XNOR2_X1  g065(.A(G143), .B(G146), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(new_n246), .ZN(new_n253));
  AND4_X1   g067(.A1(new_n251), .A2(new_n242), .A3(new_n244), .A4(new_n246), .ZN(new_n254));
  OAI22_X1  g068(.A1(new_n249), .A2(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G125), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n257));
  AND4_X1   g071(.A1(new_n257), .A2(new_n242), .A3(new_n244), .A4(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT1), .B1(new_n243), .B2(G146), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n259), .A2(G128), .B1(new_n242), .B2(new_n244), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G125), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G224), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n264), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n240), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(G210), .B1(G237), .B2(G902), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n270), .B(KEYINPUT84), .Z(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n256), .A2(KEYINPUT83), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(KEYINPUT7), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n264), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n192), .A2(KEYINPUT76), .ZN(new_n276));
  XNOR2_X1  g090(.A(G104), .B(G107), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n194), .B1(new_n277), .B2(new_n187), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n202), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n206), .A3(new_n214), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n226), .B(KEYINPUT8), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n211), .A2(G113), .A3(new_n213), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n282), .A2(KEYINPUT82), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n282), .A2(KEYINPUT82), .B1(KEYINPUT5), .B2(new_n205), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n283), .A2(new_n284), .B1(new_n205), .B2(new_n204), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n280), .B(new_n281), .C1(new_n285), .C2(new_n279), .ZN(new_n286));
  INV_X1    g100(.A(new_n274), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n256), .B(new_n263), .C1(KEYINPUT83), .C2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n275), .A2(new_n286), .A3(new_n229), .A4(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n269), .A2(new_n272), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n238), .B(new_n237), .C1(new_n231), .C2(new_n234), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n267), .B1(new_n295), .B2(new_n230), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n271), .B1(new_n296), .B2(new_n291), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n272), .B1(new_n269), .B2(new_n292), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT85), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT9), .B(G234), .ZN(new_n304));
  OAI21_X1  g118(.A(G221), .B1(new_n304), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G110), .B(G140), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n265), .A2(G227), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT11), .ZN(new_n310));
  INV_X1    g124(.A(G134), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(G137), .ZN(new_n312));
  INV_X1    g126(.A(G137), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT11), .A3(G134), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(G137), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G131), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT66), .B(G131), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(new_n314), .A3(new_n312), .A4(new_n315), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT10), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n259), .A2(G128), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n245), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n252), .A2(G128), .A3(new_n259), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n196), .A2(new_n321), .A3(new_n202), .A4(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT67), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT67), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n258), .B2(new_n260), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n279), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n330), .B2(new_n321), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT64), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT0), .B(G128), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n252), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n245), .A2(new_n248), .A3(KEYINPUT64), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT65), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n252), .A2(new_n251), .A3(new_n246), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n220), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n332), .B1(new_n342), .B2(new_n232), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n335), .A2(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n344));
  AND4_X1   g158(.A1(new_n332), .A2(new_n232), .A3(new_n220), .A4(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n320), .B(new_n331), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n279), .A2(new_n261), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n325), .A2(new_n202), .A3(new_n276), .A4(new_n278), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n317), .A2(new_n319), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT12), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT12), .ZN(new_n353));
  AOI211_X1 g167(.A(new_n353), .B(new_n320), .C1(new_n348), .C2(new_n349), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n309), .B1(new_n347), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n309), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n346), .A2(KEYINPUT77), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n331), .B1(new_n343), .B2(new_n345), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n351), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT77), .B1(new_n346), .B2(new_n357), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n356), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n290), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G469), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(G469), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n350), .A2(new_n351), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n353), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n350), .A2(KEYINPUT12), .A3(new_n351), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT79), .B1(new_n352), .B2(new_n354), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n346), .A4(new_n357), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n357), .B1(new_n360), .B2(new_n346), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n290), .B(new_n366), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n306), .B1(new_n365), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT13), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT89), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(G128), .B2(new_n243), .ZN(new_n380));
  INV_X1    g194(.A(G128), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n381), .A2(KEYINPUT89), .A3(G143), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n378), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n243), .A2(G128), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT89), .B1(new_n381), .B2(G143), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n379), .A2(new_n243), .A3(G128), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT90), .A4(KEYINPUT13), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT13), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G134), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n387), .ZN(new_n394));
  AND4_X1   g208(.A1(KEYINPUT91), .A2(new_n394), .A3(new_n311), .A4(new_n385), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT91), .B1(new_n396), .B2(new_n311), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G122), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT88), .B1(new_n399), .B2(G116), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n401));
  INV_X1    g215(.A(G116), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(G116), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n188), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n188), .A3(new_n405), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n393), .A2(new_n398), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n404), .A2(KEYINPUT14), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n400), .A2(new_n403), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n413), .A3(new_n405), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G107), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n396), .B(new_n311), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n408), .ZN(new_n417));
  INV_X1    g231(.A(G217), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n304), .A2(new_n418), .A3(G953), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n410), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n410), .B2(new_n417), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n290), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT92), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n423), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n389), .ZN(new_n430));
  INV_X1    g244(.A(new_n392), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n311), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n394), .A2(new_n311), .A3(new_n385), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT91), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n396), .A2(KEYINPUT91), .A3(new_n311), .ZN(new_n436));
  INV_X1    g250(.A(new_n408), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n435), .B(new_n436), .C1(new_n437), .C2(new_n406), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n417), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n419), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n410), .A2(new_n417), .A3(new_n419), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n428), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n290), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n429), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G113), .B(G122), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(new_n190), .ZN(new_n448));
  INV_X1    g262(.A(G237), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n265), .A3(G214), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(G143), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(G237), .A2(G953), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n454), .B(G214), .C1(new_n451), .C2(G143), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT18), .A3(G131), .ZN(new_n457));
  NOR2_X1   g271(.A1(G125), .A2(G140), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(G125), .A2(G140), .ZN(new_n460));
  AOI21_X1  g274(.A(G146), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n460), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n462), .A2(new_n458), .A3(new_n241), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT87), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G125), .B(G140), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n241), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(G146), .A3(new_n460), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(KEYINPUT18), .A2(G131), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n453), .A2(new_n455), .A3(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n457), .A2(new_n464), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n453), .A2(new_n455), .A3(new_n318), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n318), .B1(new_n453), .B2(new_n455), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT17), .ZN(new_n476));
  INV_X1    g290(.A(new_n318), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n456), .A2(KEYINPUT17), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT16), .B1(new_n462), .B2(new_n458), .ZN(new_n479));
  OR3_X1    g293(.A1(new_n262), .A2(KEYINPUT16), .A3(G140), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n241), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(G146), .A3(new_n480), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n478), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n448), .B(new_n472), .C1(new_n476), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n456), .A2(new_n477), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n473), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n489), .A2(new_n482), .A3(new_n483), .A4(new_n478), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n448), .B1(new_n490), .B2(new_n472), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n290), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G475), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n465), .A2(KEYINPUT19), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT19), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n459), .B2(new_n460), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n241), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n474), .B2(new_n475), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n483), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n479), .A2(KEYINPUT72), .A3(G146), .A4(new_n480), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n472), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n448), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n485), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n494), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  AOI211_X1 g324(.A(KEYINPUT20), .B(new_n510), .C1(new_n506), .C2(new_n485), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n493), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n265), .A2(G952), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(G234), .B2(G237), .ZN(new_n514));
  AOI211_X1 g328(.A(new_n290), .B(new_n265), .C1(G234), .C2(G237), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT21), .B(G898), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n446), .A2(new_n512), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n303), .A2(new_n377), .A3(KEYINPUT93), .A4(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n520));
  INV_X1    g334(.A(G469), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(new_n363), .B2(new_n290), .ZN(new_n522));
  INV_X1    g336(.A(new_n376), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n518), .B(new_n305), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n520), .B1(new_n524), .B2(new_n302), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n418), .B1(G234), .B2(new_n290), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n482), .A2(new_n483), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT69), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n381), .B2(G119), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n209), .A2(KEYINPUT69), .A3(G128), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n529), .A2(new_n530), .B1(G119), .B2(new_n381), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT24), .B(G110), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G110), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n381), .A2(G119), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n209), .A2(G128), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(KEYINPUT23), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(KEYINPUT23), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT23), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT70), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n540), .A2(new_n542), .A3(G119), .A4(new_n381), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n527), .B(new_n534), .C1(new_n535), .C2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(G110), .B1(new_n539), .B2(new_n543), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n531), .A2(new_n533), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT71), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n531), .A2(new_n533), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n550), .B1(new_n551), .B2(new_n546), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n501), .A2(new_n466), .A3(new_n502), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n545), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT73), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT22), .B(G137), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n545), .B(new_n559), .C1(new_n553), .C2(new_n554), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n290), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n526), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n561), .A2(new_n562), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n526), .A2(G902), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n223), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n337), .A2(new_n351), .A3(new_n341), .ZN(new_n574));
  INV_X1    g388(.A(new_n315), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n311), .A2(G137), .ZN(new_n576));
  OAI21_X1  g390(.A(G131), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n325), .A2(new_n319), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n573), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT68), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n319), .A2(new_n577), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n344), .A2(new_n351), .B1(new_n582), .B2(new_n325), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT68), .B1(new_n583), .B2(new_n573), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n329), .A2(new_n327), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n585), .A2(new_n582), .B1(new_n344), .B2(new_n351), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n573), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n581), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT28), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT28), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n454), .A2(G210), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT27), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT26), .B(G101), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n578), .B1(new_n255), .B2(new_n320), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT30), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n258), .A2(new_n260), .A3(new_n328), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT67), .B1(new_n323), .B2(new_n324), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n582), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(KEYINPUT30), .A3(new_n574), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n600), .A2(new_n604), .A3(new_n223), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n587), .A3(new_n596), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT31), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n605), .A2(KEYINPUT31), .A3(new_n587), .A4(new_n596), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n592), .A2(new_n597), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(G472), .A2(G902), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT32), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n609), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n580), .A2(new_n579), .B1(new_n586), .B2(new_n573), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n590), .B1(new_n615), .B2(new_n584), .ZN(new_n616));
  INV_X1    g430(.A(new_n591), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n597), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT32), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n611), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n613), .A2(new_n621), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n586), .A2(new_n573), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n587), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n617), .B1(new_n624), .B2(KEYINPUT28), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n596), .A2(KEYINPUT29), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n605), .A2(new_n587), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT29), .B1(new_n628), .B2(new_n597), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n629), .B1(new_n592), .B2(new_n597), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G472), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n572), .B1(new_n622), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n519), .A2(new_n525), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT94), .B(G101), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G3));
  INV_X1    g450(.A(new_n572), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n619), .A2(new_n611), .ZN(new_n638));
  OAI21_X1  g452(.A(G472), .B1(new_n610), .B2(G902), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT95), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n377), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n305), .B1(new_n522), .B2(new_n523), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT95), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n296), .A2(new_n271), .A3(new_n291), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n301), .B1(new_n299), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n290), .A2(G478), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT96), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n650), .A2(KEYINPUT96), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n651), .B(new_n652), .C1(new_n420), .C2(new_n421), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n441), .A2(KEYINPUT96), .A3(new_n650), .A4(new_n442), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(G478), .B1(new_n443), .B2(new_n290), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n517), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n659), .A3(new_n512), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n646), .A2(new_n648), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT34), .B(G104), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  NAND2_X1  g477(.A1(new_n487), .A2(new_n473), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n664), .A2(new_n501), .A3(new_n502), .A4(new_n498), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n448), .B1(new_n665), .B2(new_n472), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n508), .B1(new_n486), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT20), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n507), .A2(new_n494), .A3(new_n508), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n668), .A2(new_n669), .B1(G475), .B2(new_n492), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n446), .ZN(new_n671));
  NOR4_X1   g485(.A1(new_n646), .A2(new_n517), .A3(new_n648), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT97), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT35), .B(G107), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  NAND2_X1  g489(.A1(new_n639), .A2(new_n638), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n560), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n555), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n570), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n567), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n519), .A2(new_n525), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT37), .B(G110), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G12));
  AOI21_X1  g501(.A(new_n681), .B1(new_n622), .B2(new_n632), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n514), .B1(new_n515), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n670), .A2(new_n446), .A3(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n692), .B(new_n301), .C1(new_n299), .C2(new_n647), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n694));
  INV_X1    g508(.A(new_n301), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n293), .B2(new_n297), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n697), .A3(new_n692), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n688), .A2(new_n377), .A3(new_n694), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  XOR2_X1   g514(.A(new_n690), .B(KEYINPUT39), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n377), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT40), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n298), .A2(new_n300), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n628), .A2(new_n596), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n709), .B(new_n290), .C1(new_n596), .C2(new_n624), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n613), .A2(new_n621), .B1(G472), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n444), .B1(new_n443), .B2(new_n290), .ZN(new_n712));
  AOI211_X1 g526(.A(G902), .B(new_n428), .C1(new_n441), .C2(new_n442), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n670), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n301), .ZN(new_n716));
  OR3_X1    g530(.A1(new_n716), .A2(new_n680), .A3(KEYINPUT102), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT102), .B1(new_n716), .B2(new_n680), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n711), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n704), .A2(new_n708), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  OAI211_X1 g535(.A(new_n512), .B(new_n691), .C1(new_n655), .C2(new_n656), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n648), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n688), .A2(new_n377), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G146), .ZN(G48));
  INV_X1    g539(.A(new_n660), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n360), .A2(new_n346), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n309), .ZN(new_n728));
  AOI21_X1  g542(.A(G902), .B1(new_n728), .B2(new_n373), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n376), .B(new_n305), .C1(new_n729), .C2(new_n521), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n648), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n633), .A2(new_n726), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND2_X1  g548(.A1(new_n622), .A2(new_n632), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n671), .A2(new_n517), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n731), .A2(new_n735), .A3(new_n637), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT103), .B(G116), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G18));
  AND2_X1   g553(.A1(new_n680), .A2(new_n518), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n731), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  OAI21_X1  g556(.A(KEYINPUT105), .B1(new_n714), .B2(new_n670), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT105), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n446), .A2(new_n512), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n730), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n625), .A2(new_n596), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n612), .B1(new_n748), .B2(new_n614), .ZN(new_n749));
  AOI21_X1  g563(.A(G902), .B1(new_n614), .B2(new_n618), .ZN(new_n750));
  INV_X1    g564(.A(G472), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT104), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(G472), .C1(new_n610), .C2(G902), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n749), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  AOI211_X1 g569(.A(new_n695), .B(new_n517), .C1(new_n293), .C2(new_n297), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n747), .A2(new_n755), .A3(new_n637), .A4(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT106), .B(G122), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G24));
  XNOR2_X1  g573(.A(new_n722), .B(KEYINPUT107), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n731), .A2(new_n755), .A3(new_n680), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  NAND2_X1  g576(.A1(new_n705), .A2(new_n301), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n644), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(KEYINPUT42), .A3(new_n633), .A4(new_n760), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n695), .B1(new_n298), .B2(new_n300), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n633), .A2(new_n377), .A3(new_n760), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT108), .B(G131), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G33));
  NAND3_X1  g586(.A1(new_n633), .A2(new_n377), .A3(new_n766), .ZN(new_n773));
  INV_X1    g587(.A(new_n692), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n311), .ZN(G36));
  NAND2_X1  g590(.A1(G469), .A2(G902), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n346), .A2(new_n357), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT77), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n358), .A3(new_n360), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n781), .B2(new_n356), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT109), .B1(new_n782), .B2(new_n521), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n521), .B1(new_n363), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n363), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT45), .ZN(new_n789));
  AND4_X1   g603(.A1(KEYINPUT110), .A2(new_n783), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n785), .A2(new_n786), .B1(new_n788), .B2(KEYINPUT45), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT110), .B1(new_n791), .B2(new_n783), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n777), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n523), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n791), .A2(new_n783), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(KEYINPUT110), .A3(new_n783), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(KEYINPUT111), .A3(KEYINPUT46), .A4(new_n777), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT46), .B(new_n777), .C1(new_n790), .C2(new_n792), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n795), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n658), .A2(new_n670), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n806), .A2(KEYINPUT43), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(KEYINPUT43), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n676), .A3(new_n680), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n811), .A2(new_n812), .A3(new_n763), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n805), .A2(new_n305), .A3(new_n701), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  OR3_X1    g629(.A1(new_n735), .A2(new_n637), .A3(new_n722), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n763), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n305), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT47), .B1(new_n805), .B2(new_n305), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  AND3_X1   g635(.A1(new_n807), .A2(new_n514), .A3(new_n808), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n637), .A3(new_n755), .ZN(new_n823));
  INV_X1    g637(.A(new_n730), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n824), .B(new_n695), .C1(KEYINPUT116), .C2(KEYINPUT50), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n823), .A2(new_n708), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n637), .A2(new_n514), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n766), .A3(new_n824), .A4(new_n711), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n830), .A2(new_n512), .A3(new_n658), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT117), .Z(new_n832));
  NAND3_X1  g646(.A1(new_n822), .A2(new_n824), .A3(new_n766), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n834), .A2(new_n680), .A3(new_n755), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n828), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n729), .A2(new_n521), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n523), .A3(new_n305), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n818), .A2(new_n819), .A3(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n823), .A2(new_n763), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(KEYINPUT51), .B(new_n836), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n732), .A2(new_n757), .A3(new_n737), .A4(new_n741), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n377), .A2(new_n735), .A3(new_n766), .A4(new_n637), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n755), .A2(new_n680), .A3(new_n760), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n847), .A2(new_n692), .B1(new_n848), .B2(new_n764), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n688), .A2(new_n377), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n446), .A2(new_n512), .A3(new_n690), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n766), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n766), .A2(new_n851), .A3(new_n852), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n770), .A2(new_n846), .A3(new_n849), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n303), .A2(KEYINPUT112), .A3(new_n736), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT112), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n670), .A2(new_n446), .A3(new_n659), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n302), .B2(new_n860), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n858), .A2(new_n861), .B1(new_n303), .B2(new_n726), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n634), .B(new_n683), .C1(new_n862), .C2(new_n646), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n699), .A2(new_n724), .A3(new_n761), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n648), .A2(new_n746), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n710), .A2(G472), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n620), .B1(new_n619), .B2(new_n611), .ZN(new_n868));
  AOI211_X1 g682(.A(KEYINPUT32), .B(new_n612), .C1(new_n614), .C2(new_n618), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n567), .A2(new_n679), .A3(new_n691), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n377), .A2(new_n866), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT114), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n711), .A2(new_n871), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n377), .A4(new_n866), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n865), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT52), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n865), .A2(new_n878), .A3(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n864), .A2(new_n883), .A3(KEYINPUT53), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n864), .A2(new_n883), .A3(KEYINPUT115), .A4(KEYINPUT53), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  INV_X1    g702(.A(new_n855), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n889), .A2(new_n850), .A3(new_n853), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n732), .A2(new_n757), .A3(new_n737), .A4(new_n741), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n755), .A2(new_n760), .A3(new_n680), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n377), .A2(new_n766), .ZN(new_n893));
  OAI22_X1  g707(.A1(new_n773), .A2(new_n774), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n862), .A2(new_n646), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n634), .A2(new_n683), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n895), .A2(new_n770), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n865), .A2(new_n878), .A3(KEYINPUT52), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT52), .B1(new_n865), .B2(new_n878), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n888), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n886), .A2(new_n887), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n905), .A3(new_n884), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n834), .A2(new_n633), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT48), .Z(new_n908));
  XOR2_X1   g722(.A(new_n513), .B(KEYINPUT118), .Z(new_n909));
  NAND2_X1  g723(.A1(new_n658), .A2(new_n512), .ZN(new_n910));
  INV_X1    g724(.A(new_n731), .ZN(new_n911));
  OAI221_X1 g725(.A(new_n909), .B1(new_n910), .B2(new_n830), .C1(new_n823), .C2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n904), .A2(new_n906), .A3(new_n913), .ZN(new_n914));
  OAI22_X1  g728(.A1(new_n845), .A2(new_n914), .B1(G952), .B2(G953), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n806), .A2(new_n572), .A3(new_n695), .A4(new_n306), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT49), .B1(new_n837), .B2(new_n523), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n837), .A2(new_n523), .A3(KEYINPUT49), .ZN(new_n919));
  OR4_X1    g733(.A1(new_n708), .A2(new_n918), .A3(new_n870), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n915), .A2(new_n920), .ZN(G75));
  XOR2_X1   g735(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n864), .A2(new_n883), .A3(KEYINPUT53), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT53), .B1(new_n864), .B2(new_n883), .ZN(new_n925));
  OAI211_X1 g739(.A(G902), .B(new_n271), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n240), .B(new_n268), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT120), .Z(new_n929));
  AND3_X1   g743(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n926), .B2(new_n927), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n929), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n290), .B(new_n272), .C1(new_n902), .C2(new_n884), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(KEYINPUT56), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n922), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n265), .A2(G952), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n932), .A2(new_n937), .A3(new_n939), .ZN(G51));
  XOR2_X1   g754(.A(new_n777), .B(KEYINPUT57), .Z(new_n941));
  INV_X1    g755(.A(new_n906), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n905), .B1(new_n902), .B2(new_n884), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n375), .B2(new_n374), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n902), .A2(new_n884), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(G902), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(new_n800), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n938), .B1(new_n945), .B2(new_n948), .ZN(G54));
  NAND2_X1  g763(.A1(KEYINPUT58), .A2(G475), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT121), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n485), .B(new_n506), .C1(new_n947), .C2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n946), .A2(G902), .A3(new_n507), .A4(new_n951), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n953), .A2(new_n939), .A3(new_n954), .ZN(G60));
  AND2_X1   g769(.A1(new_n653), .A2(new_n654), .ZN(new_n956));
  NAND2_X1  g770(.A1(G478), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT59), .Z(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n942), .B2(new_n943), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n939), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n942), .B1(KEYINPUT54), .B2(new_n903), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(new_n958), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n961), .B1(new_n963), .B2(new_n956), .ZN(G63));
  INV_X1    g778(.A(KEYINPUT61), .ZN(new_n965));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT60), .Z(new_n967));
  AND2_X1   g781(.A1(new_n946), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n678), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n939), .B1(new_n968), .B2(new_n569), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n965), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n968), .A2(new_n569), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n969), .A3(KEYINPUT61), .A4(new_n939), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(G66));
  INV_X1    g789(.A(new_n516), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n265), .B1(new_n976), .B2(G224), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n863), .A2(new_n891), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT122), .Z(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n980), .B2(new_n265), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n295), .B(new_n230), .C1(G898), .C2(new_n265), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n981), .B(new_n982), .Z(G69));
  AOI21_X1  g797(.A(new_n265), .B1(G227), .B2(G900), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n633), .A2(new_n866), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n805), .A2(new_n305), .A3(new_n701), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n775), .B1(new_n765), .B2(new_n769), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n699), .A2(new_n724), .A3(new_n761), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT123), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n814), .A2(new_n986), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n820), .A3(new_n265), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n600), .A2(new_n604), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n495), .A2(new_n497), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(G900), .B2(G953), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n984), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n817), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n805), .A2(new_n305), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT47), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n305), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n720), .B1(new_n990), .B2(new_n991), .ZN(new_n1010));
  XNOR2_X1  g824(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  OAI221_X1 g828(.A(new_n720), .B1(KEYINPUT124), .B2(new_n1014), .C1(new_n990), .C2(new_n991), .ZN(new_n1015));
  INV_X1    g829(.A(new_n702), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n910), .A2(new_n671), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1016), .A2(new_n633), .A3(new_n766), .A4(new_n1017), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1013), .A2(new_n814), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n265), .B1(new_n1009), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n999), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n1001), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1003), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1021), .B(new_n1001), .C1(new_n1002), .C2(new_n984), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1023), .A2(new_n1024), .ZN(G72));
  AND4_X1   g839(.A1(new_n814), .A2(new_n1013), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n979), .A3(new_n820), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  AOI21_X1  g843(.A(new_n709), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1030), .A2(new_n938), .ZN(new_n1031));
  INV_X1    g845(.A(new_n628), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1032), .A2(new_n596), .ZN(new_n1033));
  INV_X1    g847(.A(new_n606), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1029), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT126), .Z(new_n1036));
  NAND2_X1  g850(.A1(new_n903), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT127), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT127), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n903), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n979), .A2(new_n994), .A3(new_n820), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1029), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n597), .B(new_n1032), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AND3_X1   g858(.A1(new_n1031), .A2(new_n1041), .A3(new_n1044), .ZN(G57));
endmodule


