//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n212, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G87), .ZN(G355));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n214), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n214), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n206), .A2(new_n207), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n222), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT65), .ZN(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n244), .B(new_n248), .Z(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n227), .ZN(new_n251));
  OAI21_X1  g0051(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR3_X1   g0053(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n207), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n259), .A2(new_n260), .B1(new_n228), .B2(G68), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n251), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT11), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(KEYINPUT11), .B(new_n251), .C1(new_n256), .C2(new_n261), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT74), .B1(new_n268), .B2(G68), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT12), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n268), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n251), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n267), .A2(G20), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(G68), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n271), .A2(KEYINPUT75), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(KEYINPUT75), .B1(new_n271), .B2(new_n275), .ZN(new_n278));
  NOR3_X1   g0078(.A1(new_n266), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT14), .ZN(new_n281));
  AND2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  OAI211_X1 g0083(.A(G232), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT73), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n257), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT73), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(G232), .A4(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G97), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n289), .A2(G226), .A3(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n285), .A2(new_n291), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(G1), .A3(G13), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n297), .A3(G274), .ZN(new_n302));
  INV_X1    g0102(.A(G238), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n297), .A2(new_n300), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT13), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT13), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n299), .A2(new_n309), .A3(new_n306), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n281), .B1(new_n311), .B2(G169), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n309), .B1(new_n299), .B2(new_n306), .ZN(new_n313));
  AOI211_X1 g0113(.A(KEYINPUT13), .B(new_n305), .C1(new_n295), .C2(new_n298), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n281), .B(G169), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n308), .A2(G179), .A3(new_n310), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n280), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n308), .A2(G190), .A3(new_n310), .ZN(new_n319));
  OAI21_X1  g0119(.A(G200), .B1(new_n313), .B2(new_n314), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n279), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT8), .B(G58), .Z(new_n323));
  AND2_X1   g0123(.A1(new_n323), .A2(new_n274), .ZN(new_n324));
  INV_X1    g0124(.A(new_n323), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(new_n273), .B1(new_n325), .B2(new_n272), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n251), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n282), .A2(new_n283), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT7), .B1(new_n329), .B2(new_n228), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  NOR4_X1   g0131(.A1(new_n282), .A2(new_n283), .A3(new_n331), .A4(G20), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n334));
  OR3_X1    g0134(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n252), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n334), .A2(G20), .B1(new_n336), .B2(G159), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n328), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT76), .B1(new_n282), .B2(new_n283), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT76), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n287), .A2(new_n342), .A3(new_n288), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n343), .A3(new_n228), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n332), .B1(new_n344), .B2(new_n331), .ZN(new_n345));
  OAI211_X1 g0145(.A(KEYINPUT16), .B(new_n337), .C1(new_n345), .C2(new_n203), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n327), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(G223), .B(new_n293), .C1(new_n282), .C2(new_n283), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT77), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n293), .B1(new_n287), .B2(new_n288), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G226), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT77), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n289), .A2(new_n352), .A3(G223), .A4(new_n293), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G87), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n349), .A2(new_n351), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n298), .ZN(new_n356));
  INV_X1    g0156(.A(G190), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n297), .A2(G232), .A3(new_n300), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT78), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT78), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n297), .A2(new_n300), .A3(new_n361), .A4(G232), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n302), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT79), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT79), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n360), .A2(new_n365), .A3(new_n302), .A4(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n363), .B1(new_n355), .B2(new_n298), .ZN(new_n368));
  OAI22_X1  g0168(.A1(new_n358), .A2(new_n367), .B1(new_n368), .B2(G200), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n347), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT17), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(KEYINPUT80), .A2(KEYINPUT18), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n356), .A2(new_n374), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n375), .A2(new_n367), .B1(new_n368), .B2(G169), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n373), .B1(new_n347), .B2(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n364), .A2(new_n366), .ZN(new_n378));
  AOI21_X1  g0178(.A(G179), .B1(new_n355), .B2(new_n298), .ZN(new_n379));
  INV_X1    g0179(.A(new_n363), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n356), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G169), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n378), .A2(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n331), .B1(new_n289), .B2(G20), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n203), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n202), .A2(new_n203), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n206), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n336), .A2(G159), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n339), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n251), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n344), .A2(new_n331), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n203), .B1(new_n393), .B2(new_n385), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n337), .A2(KEYINPUT16), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n326), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(KEYINPUT80), .A2(KEYINPUT18), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n373), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n383), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n347), .A2(new_n369), .A3(KEYINPUT17), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n372), .A2(new_n377), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n322), .A2(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n336), .A2(G150), .B1(new_n323), .B2(new_n258), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n208), .A2(G20), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n328), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n273), .A2(G50), .A3(new_n274), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(G50), .B2(new_n268), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n302), .ZN(new_n411));
  INV_X1    g0211(.A(new_n304), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(G226), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n350), .A2(G223), .B1(new_n329), .B2(G77), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n289), .A2(G222), .A3(new_n293), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n413), .B1(new_n416), .B2(new_n297), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n410), .B1(new_n417), .B2(new_n382), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G179), .B2(new_n417), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n410), .A2(KEYINPUT9), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT71), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT10), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n410), .A2(KEYINPUT9), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n417), .A2(G200), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n417), .A2(new_n357), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n421), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n422), .B1(new_n421), .B2(new_n426), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n419), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n273), .A2(G77), .A3(new_n274), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(G77), .B2(new_n268), .ZN(new_n431));
  XOR2_X1   g0231(.A(KEYINPUT15), .B(G87), .Z(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n258), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT69), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n336), .A2(new_n323), .B1(G20), .B2(G77), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n431), .B1(new_n436), .B2(new_n251), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n293), .A2(G232), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n303), .A2(new_n293), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n289), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n211), .B2(new_n289), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT68), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n297), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n443), .B2(new_n442), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n411), .B1(G244), .B2(new_n412), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n438), .B(KEYINPUT70), .C1(new_n447), .C2(G169), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT70), .ZN(new_n449));
  AOI21_X1  g0249(.A(G169), .B1(new_n445), .B2(new_n446), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(new_n437), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n374), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n447), .A2(G190), .ZN(new_n454));
  INV_X1    g0254(.A(G200), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n437), .C1(new_n455), .C2(new_n447), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n429), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT72), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT72), .B1(new_n429), .B2(new_n457), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n404), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n228), .B(G87), .C1(new_n282), .C2(new_n283), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT22), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT22), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n289), .A2(new_n466), .A3(new_n228), .A4(G87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT24), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G116), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G20), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n228), .B2(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n211), .A2(KEYINPUT23), .A3(G20), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n468), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n469), .B1(new_n468), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n251), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n267), .A2(G33), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n273), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT25), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n268), .B2(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n272), .A2(KEYINPUT25), .A3(new_n211), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n481), .A2(G107), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(G257), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n487));
  OAI211_X1 g0287(.A(G250), .B(new_n293), .C1(new_n282), .C2(new_n283), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G294), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n298), .ZN(new_n491));
  INV_X1    g0291(.A(G274), .ZN(new_n492));
  INV_X1    g0292(.A(new_n227), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(new_n493), .B2(new_n296), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT5), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(G41), .ZN(new_n497));
  INV_X1    g0297(.A(G41), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n267), .B(G45), .C1(new_n498), .C2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT83), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G45), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(G1), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n496), .A2(G41), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT83), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n494), .B(new_n500), .C1(new_n503), .C2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n496), .A2(G41), .ZN(new_n509));
  OAI211_X1 g0309(.A(G264), .B(new_n297), .C1(new_n501), .C2(new_n509), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n491), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n357), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n508), .A2(new_n510), .ZN(new_n513));
  AOI21_X1  g0313(.A(G200), .B1(new_n513), .B2(new_n491), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT90), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n511), .A2(KEYINPUT90), .A3(new_n357), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n486), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n485), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n468), .A2(new_n475), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT24), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n468), .A2(new_n469), .A3(new_n475), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n519), .B1(new_n523), .B2(new_n251), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n511), .A2(new_n374), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n491), .A2(new_n508), .A3(new_n510), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n382), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT91), .B1(new_n518), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n515), .B1(new_n526), .B2(new_n455), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n526), .A2(G190), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n517), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n524), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n486), .A2(new_n525), .A3(new_n527), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT91), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n505), .A2(new_n492), .ZN(new_n539));
  INV_X1    g0339(.A(G250), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n504), .B2(G1), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n297), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n303), .A2(new_n293), .ZN(new_n544));
  INV_X1    g0344(.A(G244), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G1698), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n544), .B(new_n546), .C1(new_n282), .C2(new_n283), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n470), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n297), .B1(new_n548), .B2(KEYINPUT85), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT85), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n550), .A3(new_n470), .ZN(new_n551));
  AOI211_X1 g0351(.A(KEYINPUT86), .B(new_n543), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT86), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(KEYINPUT85), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n298), .A3(new_n551), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(new_n542), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n382), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n547), .A2(new_n550), .A3(new_n470), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n550), .B1(new_n547), .B2(new_n470), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n558), .A2(new_n559), .A3(new_n297), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT86), .B1(new_n560), .B2(new_n543), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n555), .A2(new_n553), .A3(new_n542), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n374), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n259), .B2(new_n210), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n289), .A2(new_n228), .A3(G68), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n228), .B1(new_n292), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(G87), .B2(new_n212), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n251), .ZN(new_n570));
  INV_X1    g0370(.A(new_n432), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n272), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n572), .C1(new_n571), .C2(new_n480), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n557), .A2(new_n563), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n552), .B2(new_n556), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n561), .A2(G190), .A3(new_n562), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n572), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(G87), .B2(new_n481), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT87), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT87), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n574), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(G244), .B(new_n293), .C1(new_n282), .C2(new_n283), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT4), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G283), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n289), .A2(G250), .A3(G1698), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(KEYINPUT4), .A2(G244), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n293), .B(new_n590), .C1(new_n282), .C2(new_n283), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n289), .A2(KEYINPUT82), .A3(new_n293), .A4(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n298), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(G257), .B(new_n297), .C1(new_n501), .C2(new_n509), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n508), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G200), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n600), .A2(new_n210), .A3(G107), .ZN(new_n601));
  XNOR2_X1  g0401(.A(G97), .B(G107), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n603), .A2(new_n228), .B1(new_n260), .B2(new_n255), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n211), .B1(new_n384), .B2(new_n385), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n251), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n268), .A2(G97), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n607), .B(KEYINPUT81), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(G97), .B2(new_n481), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n597), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n350), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n613), .A2(new_n586), .A3(new_n593), .A4(new_n594), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n614), .B2(new_n298), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(G190), .A3(new_n508), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n599), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n598), .A2(new_n382), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n374), .A3(new_n508), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(new_n619), .A3(new_n610), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(G270), .B(new_n297), .C1(new_n501), .C2(new_n509), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n508), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n273), .A2(G116), .A3(new_n479), .ZN(new_n624));
  OR3_X1    g0424(.A1(new_n268), .A2(KEYINPUT88), .A3(G116), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT88), .B1(new_n268), .B2(G116), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G116), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n250), .A2(new_n227), .B1(G20), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n587), .B(new_n228), .C1(G33), .C2(new_n210), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n629), .A2(KEYINPUT20), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT20), .B1(new_n629), .B2(new_n630), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n624), .B(new_n627), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(G257), .B(new_n293), .C1(new_n282), .C2(new_n283), .ZN(new_n634));
  OAI211_X1 g0434(.A(G264), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n287), .A2(G303), .A3(new_n288), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n298), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n623), .A2(new_n633), .A3(G179), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n508), .A3(new_n622), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT89), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT21), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n640), .A2(new_n633), .A3(G169), .A4(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n633), .B1(new_n640), .B2(G200), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n357), .B2(new_n640), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n640), .A2(new_n633), .A3(G169), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n641), .A3(new_n642), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n645), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n621), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n581), .A2(new_n583), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n463), .A2(new_n538), .A3(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n419), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT94), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n347), .B2(new_n376), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n383), .A2(new_n397), .A3(KEYINPUT94), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT18), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n318), .ZN(new_n663));
  INV_X1    g0463(.A(new_n453), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n321), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n372), .A2(new_n401), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT95), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n427), .A2(new_n428), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n669), .B1(new_n667), .B2(KEYINPUT95), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n654), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n610), .B1(G200), .B2(new_n598), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n598), .A2(new_n382), .B1(new_n606), .B2(new_n609), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n672), .A2(new_n616), .B1(new_n673), .B2(new_n619), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n555), .A2(new_n542), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n382), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n563), .A2(new_n676), .A3(new_n573), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(G200), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n576), .A2(new_n578), .A3(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n674), .A2(new_n534), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n649), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n639), .A2(new_n644), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT92), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT92), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n645), .A2(new_n684), .A3(new_n649), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n529), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT93), .B1(new_n680), .B2(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n681), .A2(new_n682), .A3(KEYINPUT92), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n684), .B1(new_n645), .B2(new_n649), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n535), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n677), .A2(new_n679), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n621), .A2(new_n518), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n690), .A2(new_n691), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n620), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n677), .A3(new_n679), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n677), .B1(new_n697), .B2(KEYINPUT26), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n581), .A2(new_n583), .A3(new_n696), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(KEYINPUT26), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n462), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n671), .A2(new_n702), .ZN(G369));
  NAND3_X1  g0503(.A1(new_n267), .A2(new_n228), .A3(G13), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT96), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n535), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n486), .A2(new_n710), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n530), .A2(new_n537), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n529), .A2(new_n710), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT97), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT97), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n713), .A2(new_n717), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n681), .A2(new_n682), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n710), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n711), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n710), .A2(new_n633), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n647), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n683), .A2(new_n685), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n724), .B1(new_n725), .B2(new_n723), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n719), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n722), .A2(new_n729), .ZN(G399));
  INV_X1    g0530(.A(new_n223), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G41), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n212), .A2(G87), .A3(G116), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(G1), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n226), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(new_n733), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  INV_X1    g0538(.A(new_n710), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n701), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n720), .A2(new_n535), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n693), .A2(new_n692), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n677), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n697), .B2(KEYINPUT26), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n574), .A2(new_n579), .A3(new_n582), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n582), .B1(new_n574), .B2(new_n579), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT26), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(new_n751), .A3(new_n696), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n710), .B1(new_n747), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT99), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(new_n754), .A3(KEYINPUT29), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n699), .A2(KEYINPUT26), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n744), .A2(new_n746), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n739), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT99), .B1(new_n758), .B2(new_n741), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n742), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n534), .A2(new_n536), .A3(new_n535), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n536), .B1(new_n534), .B2(new_n535), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n750), .A2(new_n763), .A3(new_n651), .A4(new_n739), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n638), .A2(G179), .A3(new_n508), .A4(new_n622), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n526), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n766), .A2(new_n561), .A3(new_n562), .A4(new_n615), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT30), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n596), .A2(new_n597), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n770), .A2(new_n526), .A3(new_n765), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n552), .A2(new_n556), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT30), .ZN(new_n773));
  AOI21_X1  g0573(.A(G179), .B1(new_n555), .B2(new_n542), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n598), .A2(new_n774), .A3(new_n526), .A4(new_n640), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n769), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  AND3_X1   g0576(.A1(new_n776), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n777));
  AOI21_X1  g0577(.A(KEYINPUT31), .B1(new_n776), .B2(new_n710), .ZN(new_n778));
  OAI21_X1  g0578(.A(KEYINPUT98), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n764), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G330), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n760), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n738), .B1(new_n783), .B2(G1), .ZN(G364));
  AOI21_X1  g0584(.A(new_n227), .B1(G20), .B2(new_n382), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G179), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n210), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n228), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n786), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G159), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n790), .B1(KEYINPUT32), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n228), .A2(new_n374), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n796), .A2(new_n357), .A3(G200), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(KEYINPUT32), .B2(new_n794), .C1(new_n203), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n228), .A2(new_n357), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n455), .A2(G179), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT104), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT104), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G87), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n374), .A2(G200), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n791), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n329), .B1(new_n809), .B2(G77), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n799), .A2(new_n807), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n791), .A2(new_n800), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G58), .A2(new_n812), .B1(new_n814), .B2(G107), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n806), .A2(new_n810), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n796), .A2(G190), .A3(G200), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT103), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n817), .A2(new_n818), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n798), .B(new_n816), .C1(G50), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n289), .B1(new_n812), .B2(G322), .ZN(new_n825));
  INV_X1    g0625(.A(G294), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT33), .B(G317), .Z(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n789), .C1(new_n797), .C2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G311), .A2(new_n809), .B1(new_n793), .B2(G329), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  INV_X1    g0630(.A(G303), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n830), .B2(new_n813), .C1(new_n804), .C2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n828), .B(new_n832), .C1(G326), .C2(new_n823), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n785), .B1(new_n824), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n228), .A2(G13), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n267), .B1(new_n835), .B2(G45), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n732), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(G13), .A2(G33), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(G20), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n731), .A2(new_n329), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT100), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(G355), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT100), .B1(new_n212), .B2(G87), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n845), .A2(new_n846), .B1(G116), .B2(new_n223), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n248), .A2(G45), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n341), .A2(new_n343), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n731), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n504), .B2(new_n226), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n847), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n842), .B(new_n785), .C1(new_n853), .C2(KEYINPUT101), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n839), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n834), .B1(new_n856), .B2(KEYINPUT102), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(KEYINPUT102), .B2(new_n856), .ZN(new_n858));
  INV_X1    g0658(.A(new_n842), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n726), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n728), .A2(new_n838), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(G330), .B2(new_n726), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G396));
  NOR2_X1   g0664(.A1(new_n739), .A2(new_n437), .ZN(new_n865));
  MUX2_X1   g0665(.A(new_n457), .B(new_n453), .S(new_n865), .Z(new_n866));
  NAND2_X1  g0666(.A1(new_n740), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n457), .A2(new_n710), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n687), .A2(new_n694), .ZN(new_n869));
  INV_X1    g0669(.A(new_n698), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n748), .A2(new_n749), .A3(new_n620), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(new_n751), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n868), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  OR3_X1    g0674(.A1(new_n874), .A2(KEYINPUT105), .A3(new_n782), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT105), .B1(new_n874), .B2(new_n782), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n838), .B1(new_n874), .B2(new_n782), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n866), .A2(new_n840), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n785), .A2(new_n840), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n838), .B1(G77), .B2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(G143), .A2(new_n812), .B1(new_n809), .B2(G159), .ZN(new_n883));
  INV_X1    g0683(.A(G150), .ZN(new_n884));
  INV_X1    g0684(.A(G137), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n883), .B1(new_n884), .B2(new_n797), .C1(new_n822), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT34), .ZN(new_n887));
  AOI22_X1  g0687(.A1(G68), .A2(new_n814), .B1(new_n793), .B2(G132), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n888), .B(new_n849), .C1(new_n202), .C2(new_n789), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(G50), .B2(new_n805), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n822), .A2(new_n831), .ZN(new_n892));
  INV_X1    g0692(.A(G311), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n329), .B1(new_n792), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n797), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n894), .B(new_n790), .C1(G283), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n814), .A2(G87), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n826), .B2(new_n811), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(G116), .B2(new_n809), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n896), .B(new_n899), .C1(new_n211), .C2(new_n804), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n891), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n882), .B1(new_n901), .B2(new_n785), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n877), .A2(new_n878), .B1(new_n879), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(G384));
  XNOR2_X1  g0704(.A(new_n603), .B(KEYINPUT106), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT35), .ZN(new_n906));
  OAI211_X1 g0706(.A(G116), .B(new_n229), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n906), .B2(new_n905), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT36), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n226), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n207), .A2(G68), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n267), .B(G13), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n453), .A2(new_n710), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n873), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT37), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n339), .B1(new_n394), .B2(new_n390), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n251), .A3(new_n346), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n326), .ZN(new_n921));
  INV_X1    g0721(.A(new_n708), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n921), .A2(new_n922), .B1(new_n347), .B2(new_n369), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n383), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n397), .A2(new_n922), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n370), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n347), .A2(new_n376), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT37), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n920), .A2(new_n326), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n708), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n402), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(KEYINPUT108), .B(new_n917), .C1(new_n930), .C2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n917), .B1(new_n930), .B2(new_n933), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n402), .A2(new_n932), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n937), .B(KEYINPUT38), .C1(new_n925), .C2(new_n929), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT107), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n313), .A2(new_n314), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT14), .B1(new_n941), .B2(new_n382), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n321), .A2(new_n942), .A3(new_n316), .A4(new_n315), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n279), .A2(new_n739), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n944), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n318), .A2(new_n321), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n318), .A2(new_n940), .A3(new_n321), .A4(new_n946), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n916), .A2(new_n934), .A3(new_n939), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n660), .A2(new_n661), .A3(new_n708), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n938), .A2(new_n936), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n370), .B1(new_n931), .B2(new_n708), .ZN(new_n954));
  INV_X1    g0754(.A(new_n924), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT37), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n927), .A2(KEYINPUT37), .A3(new_n928), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT38), .B1(new_n958), .B2(new_n937), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n934), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT39), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n666), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n926), .B1(new_n662), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n927), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n918), .B1(new_n965), .B2(new_n658), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(new_n929), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n917), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n938), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT39), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n962), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n663), .A2(new_n739), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n951), .B(new_n952), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n742), .A2(new_n462), .A3(new_n759), .A4(new_n755), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n671), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n974), .B(new_n976), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n960), .A2(KEYINPUT40), .A3(new_n961), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n777), .A2(new_n778), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n764), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n664), .A2(new_n865), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n457), .B2(new_n865), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n950), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n948), .A2(new_n949), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(new_n866), .ZN(new_n985));
  INV_X1    g0785(.A(new_n661), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT18), .B1(new_n656), .B2(new_n657), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n963), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(new_n397), .A3(new_n922), .ZN(new_n989));
  INV_X1    g0789(.A(new_n967), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT38), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n938), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n985), .B(new_n980), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n978), .A2(new_n983), .B1(new_n993), .B2(KEYINPUT40), .ZN(new_n994));
  INV_X1    g0794(.A(new_n980), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n463), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT40), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n983), .A2(new_n997), .A3(new_n934), .A4(new_n939), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n666), .B1(new_n660), .B2(new_n661), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n999), .A2(new_n926), .B1(new_n929), .B2(new_n966), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n992), .B1(new_n917), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n950), .A2(new_n980), .A3(new_n982), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT40), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1004), .A2(new_n462), .A3(new_n980), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n996), .A2(G330), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n977), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n267), .B2(new_n835), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n977), .A2(new_n1006), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n913), .B1(new_n1008), .B2(new_n1009), .ZN(G367));
  INV_X1    g0810(.A(new_n783), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n713), .A2(new_n717), .A3(new_n714), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n717), .B1(new_n713), .B2(new_n714), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n721), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n711), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT45), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n674), .B1(new_n611), .B2(new_n739), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n696), .A2(new_n710), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NOR3_X1   g0821(.A1(new_n1016), .A2(new_n1017), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(KEYINPUT45), .B1(new_n722), .B2(new_n1020), .ZN(new_n1023));
  AOI21_X1  g0823(.A(KEYINPUT44), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT44), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1025), .B(new_n1020), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n1022), .A2(new_n1023), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n729), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1025), .B1(new_n722), .B2(new_n1020), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1016), .A2(KEYINPUT44), .A3(new_n1021), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n729), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n719), .A2(new_n721), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n728), .A3(new_n1014), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1014), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n727), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  AND4_X1   g0838(.A1(new_n760), .A2(new_n1036), .A3(new_n782), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1029), .A2(new_n1033), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT113), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1029), .A2(new_n1033), .A3(KEYINPUT113), .A4(new_n1039), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1011), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n732), .B(KEYINPUT41), .Z(new_n1045));
  OAI21_X1  g0845(.A(new_n836), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n739), .A2(new_n578), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT109), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n692), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n677), .B2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(KEYINPUT43), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT111), .Z(new_n1052));
  OAI21_X1  g0852(.A(new_n620), .B1(new_n1018), .B2(new_n535), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT110), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n1055), .A2(new_n739), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n719), .A2(new_n721), .A3(new_n1020), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1057), .B1(KEYINPUT42), .B2(new_n1058), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1058), .A2(KEYINPUT42), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1052), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1050), .A2(KEYINPUT43), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT112), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  OR3_X1    g0865(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1064), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n729), .A2(new_n1021), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1046), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n842), .A2(new_n785), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n223), .B2(new_n571), .C1(new_n851), .C2(new_n239), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n838), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n814), .A2(G77), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n207), .B2(new_n808), .C1(new_n885), .C2(new_n792), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n329), .B1(new_n812), .B2(G150), .ZN(new_n1077));
  INV_X1    g0877(.A(G159), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1077), .B1(new_n203), .B2(new_n789), .C1(new_n1078), .C2(new_n797), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1076), .B(new_n1079), .C1(G58), .C2(new_n805), .ZN(new_n1080));
  INV_X1    g0880(.A(G143), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n1081), .B2(new_n822), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT115), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT114), .B1(new_n805), .B2(G116), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT46), .Z(new_n1085));
  INV_X1    g0885(.A(new_n849), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n826), .B2(new_n797), .C1(new_n211), .C2(new_n789), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n811), .A2(new_n831), .B1(new_n808), .B2(new_n830), .ZN(new_n1088));
  INV_X1    g0888(.A(G317), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n813), .A2(new_n210), .B1(new_n792), .B2(new_n1089), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1087), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n893), .B2(new_n822), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1083), .B1(new_n1085), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT47), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1074), .B1(new_n1094), .B2(new_n785), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1050), .A2(new_n859), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1071), .A2(new_n1097), .ZN(G387));
  NOR2_X1   g0898(.A1(new_n1039), .A2(new_n733), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n783), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n837), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n734), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n843), .A2(new_n1103), .B1(new_n211), .B2(new_n731), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n236), .A2(new_n504), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n323), .A2(new_n207), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT50), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n734), .B(new_n504), .C1(new_n203), .C2(new_n260), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n850), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1104), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n839), .B1(new_n1110), .B2(new_n1072), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n785), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n788), .A2(new_n432), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n849), .C1(new_n325), .C2(new_n797), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G97), .A2(new_n814), .B1(new_n793), .B2(G150), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G50), .A2(new_n812), .B1(new_n809), .B2(G68), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(new_n804), .C2(new_n260), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1114), .B(new_n1117), .C1(G159), .C2(new_n823), .ZN(new_n1118));
  INV_X1    g0918(.A(G326), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n813), .A2(new_n628), .B1(new_n792), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G317), .A2(new_n812), .B1(new_n809), .B2(G303), .ZN(new_n1121));
  INV_X1    g0921(.A(G322), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1121), .B1(new_n893), .B2(new_n797), .C1(new_n822), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT48), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n805), .A2(G294), .B1(G283), .B2(new_n788), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n849), .B(new_n1120), .C1(new_n1129), .C2(KEYINPUT49), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1129), .A2(KEYINPUT49), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1118), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1111), .B1(new_n1112), .B2(new_n1132), .C1(new_n719), .C2(new_n859), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1101), .A2(new_n1102), .A3(new_n1133), .ZN(G393));
  OAI221_X1 g0934(.A(new_n1072), .B1(new_n210), .B2(new_n223), .C1(new_n244), .C2(new_n851), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1135), .A2(KEYINPUT116), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(KEYINPUT116), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n838), .A3(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n822), .A2(new_n884), .B1(new_n1078), .B2(new_n811), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT51), .Z(new_n1140));
  NOR2_X1   g0940(.A1(new_n804), .A2(new_n203), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n849), .B1(new_n797), .B2(new_n207), .C1(new_n789), .C2(new_n260), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n897), .B1(new_n1081), .B2(new_n792), .C1(new_n325), .C2(new_n808), .ZN(new_n1143));
  OR3_X1    g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n822), .A2(new_n1089), .B1(new_n893), .B2(new_n811), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT52), .Z(new_n1146));
  OAI22_X1  g0946(.A1(new_n789), .A2(new_n628), .B1(new_n797), .B2(new_n831), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n329), .B1(new_n813), .B2(new_n211), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n808), .A2(new_n826), .B1(new_n792), .B2(new_n1122), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n830), .B2(new_n804), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1140), .A2(new_n1144), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1138), .B1(new_n1152), .B2(new_n785), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n1020), .B2(new_n859), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n836), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1039), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n733), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1156), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(G390));
  INV_X1    g0961(.A(new_n868), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n695), .B2(new_n700), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n950), .B1(new_n1163), .B2(new_n914), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n962), .A2(new_n971), .B1(new_n1164), .B2(new_n973), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n982), .B(new_n739), .C1(new_n756), .C2(new_n757), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n984), .B1(new_n1166), .B2(new_n915), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n973), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n1001), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n781), .A2(new_n950), .A3(G330), .A4(new_n982), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1165), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(G330), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n764), .B2(new_n979), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n985), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n984), .B1(new_n873), .B2(new_n915), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n970), .B1(new_n939), .B2(new_n934), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT39), .B1(new_n968), .B2(new_n938), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1176), .A2(new_n1168), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n914), .B1(new_n753), .B2(new_n982), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n973), .B(new_n969), .C1(new_n1180), .C2(new_n984), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1175), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1172), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n972), .A2(new_n840), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n838), .B1(new_n323), .B2(new_n881), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n804), .A2(new_n884), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1186), .B(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(G125), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n289), .B1(new_n792), .B2(new_n1189), .C1(new_n789), .C2(new_n1078), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n812), .A2(G132), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1191), .B1(new_n207), .B2(new_n813), .C1(new_n808), .C2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1190), .B(new_n1193), .C1(G137), .C2(new_n895), .ZN(new_n1194));
  INV_X1    g0994(.A(G128), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1188), .B(new_n1194), .C1(new_n1195), .C2(new_n822), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n797), .A2(new_n211), .B1(new_n808), .B2(new_n210), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n823), .B2(G283), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT119), .Z(new_n1199));
  AOI22_X1  g0999(.A1(new_n812), .A2(G116), .B1(new_n788), .B2(G77), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT121), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n813), .A2(new_n203), .B1(new_n792), .B2(new_n826), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT120), .Z(new_n1203));
  NAND4_X1  g1003(.A1(new_n806), .A2(new_n1201), .A3(new_n1203), .A4(new_n329), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1196), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1185), .B1(new_n1205), .B2(new_n785), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1183), .A2(new_n837), .B1(new_n1184), .B2(new_n1206), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n652), .A2(new_n538), .A3(new_n710), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n778), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n776), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(G330), .B(new_n982), .C1(new_n1208), .C2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n984), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n1180), .A3(new_n1170), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n781), .A2(G330), .A3(new_n982), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1215), .A2(new_n984), .B1(new_n985), .B2(new_n1174), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1163), .A2(new_n914), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n462), .A2(new_n1174), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1218), .A2(new_n671), .A3(new_n975), .A4(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(KEYINPUT117), .C1(new_n1172), .C2(new_n1182), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1175), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1179), .A2(new_n1181), .A3(new_n1170), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n975), .A2(new_n671), .A3(new_n1219), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1218), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1221), .A2(new_n732), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT117), .B1(new_n1228), .B2(new_n1220), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1207), .B1(new_n1227), .B2(new_n1229), .ZN(G378));
  OAI211_X1 g1030(.A(new_n429), .B(new_n922), .C1(new_n407), .C2(new_n409), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n419), .B1(new_n410), .B2(new_n708), .C1(new_n427), .C2(new_n428), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1004), .B2(G330), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1173), .B(new_n1236), .C1(new_n998), .C2(new_n1003), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n974), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1236), .B1(new_n994), .B2(new_n1173), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n962), .A2(new_n971), .A3(new_n1168), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1242), .A2(new_n951), .A3(new_n952), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1004), .A2(G330), .A3(new_n1237), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1241), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1240), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1236), .A2(new_n840), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n881), .A2(G50), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n812), .A2(G107), .B1(new_n809), .B2(new_n432), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n203), .B2(new_n789), .C1(new_n210), .C2(new_n797), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1086), .A2(new_n498), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n813), .A2(new_n202), .B1(new_n792), .B2(new_n830), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n805), .C2(G77), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT122), .Z(new_n1254));
  AOI211_X1 g1054(.A(new_n1250), .B(new_n1254), .C1(G116), .C2(new_n823), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(G33), .A2(G41), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(G50), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1255), .A2(KEYINPUT58), .B1(new_n1251), .B2(new_n1257), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n811), .A2(new_n1195), .B1(new_n808), .B2(new_n885), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n789), .A2(new_n884), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(G132), .C2(new_n895), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1261), .B1(new_n1189), .B2(new_n822), .C1(new_n804), .C2(new_n1192), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1264));
  INV_X1    g1064(.A(G124), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1256), .B1(new_n792), .B2(new_n1265), .C1(new_n1078), .C2(new_n813), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT123), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1258), .B1(KEYINPUT58), .B2(new_n1255), .C1(new_n1263), .C2(new_n1268), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n839), .B(new_n1248), .C1(new_n1269), .C2(new_n785), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1246), .A2(new_n837), .B1(new_n1247), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1245), .A2(new_n1240), .B1(new_n1226), .B2(new_n1225), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(KEYINPUT57), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n733), .B1(new_n1273), .B2(KEYINPUT57), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1272), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(G375));
  NAND2_X1  g1078(.A1(new_n895), .A2(G116), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1279), .A2(new_n329), .A3(new_n1075), .A4(new_n1113), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(G283), .A2(new_n812), .B1(new_n809), .B2(G107), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n1281), .B1(new_n831), .B2(new_n792), .C1(new_n804), .C2(new_n210), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n1280), .B(new_n1282), .C1(G294), .C2(new_n823), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n849), .B1(new_n797), .B2(new_n1192), .C1(new_n789), .C2(new_n207), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(G137), .A2(new_n812), .B1(new_n814), .B2(G58), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G150), .A2(new_n809), .B1(new_n793), .B2(G128), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1285), .B(new_n1286), .C1(new_n804), .C2(new_n1078), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1284), .B(new_n1287), .C1(G132), .C2(new_n823), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n785), .B1(new_n1283), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n839), .B1(new_n203), .B2(new_n880), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1289), .B(new_n1290), .C1(new_n950), .C2(new_n841), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1218), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(new_n836), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1045), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1220), .A2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1225), .A2(new_n1218), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(KEYINPUT124), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(G381));
  OR4_X1    g1100(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G378), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(KEYINPUT125), .B(new_n1207), .C1(new_n1227), .C2(new_n1229), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1277), .A2(new_n1303), .A3(new_n1304), .ZN(new_n1305));
  OR4_X1    g1105(.A1(G387), .A2(new_n1301), .A3(G381), .A4(new_n1305), .ZN(G407));
  OAI211_X1 g1106(.A(G407), .B(G213), .C1(G343), .C2(new_n1305), .ZN(G409));
  NAND2_X1  g1107(.A1(new_n709), .A2(G213), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1226), .A2(new_n1225), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1246), .A2(new_n1310), .A3(new_n1295), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1271), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1303), .A2(new_n1304), .A3(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1246), .A2(new_n1310), .A3(KEYINPUT57), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n732), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G378), .B(new_n1271), .C1(new_n1315), .C2(new_n1274), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1309), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n975), .A2(new_n671), .A3(new_n1219), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1292), .A2(KEYINPUT60), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT126), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT126), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1292), .A2(new_n1319), .A3(new_n1322), .A4(KEYINPUT60), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1220), .A2(new_n732), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT60), .B1(new_n1292), .B2(new_n1319), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(G384), .B1(new_n1328), .B2(new_n1294), .ZN(new_n1329));
  AOI211_X1 g1129(.A(new_n1293), .B(new_n903), .C1(new_n1324), .C2(new_n1327), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1317), .A2(new_n1318), .A3(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1329), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1330), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1309), .A2(G2897), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1334), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  OAI211_X1 g1137(.A(G2897), .B(new_n1309), .C1(new_n1329), .C2(new_n1330), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1333), .B1(new_n1317), .B2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1318), .B1(new_n1317), .B2(new_n1331), .ZN(new_n1341));
  NOR3_X1   g1141(.A1(new_n1332), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G387), .A2(new_n1160), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(G393), .B(new_n863), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1071), .A2(new_n1097), .A3(G390), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1344), .ZN(new_n1347));
  AOI21_X1  g1147(.A(G390), .B1(new_n1071), .B2(new_n1097), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1097), .ZN(new_n1349));
  AOI211_X1 g1149(.A(new_n1349), .B(new_n1160), .C1(new_n1046), .C2(new_n1070), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1347), .B1(new_n1348), .B2(new_n1350), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1346), .A2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT63), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1308), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1331), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1353), .B1(new_n1355), .B2(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1317), .A2(KEYINPUT63), .A3(new_n1331), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  AND2_X1   g1159(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1355), .A2(new_n1360), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1361), .A2(new_n1346), .A3(new_n1351), .A4(new_n1333), .ZN(new_n1362));
  OAI22_X1  g1162(.A1(new_n1342), .A2(new_n1352), .B1(new_n1359), .B2(new_n1362), .ZN(G405));
  AOI21_X1  g1163(.A(KEYINPUT127), .B1(new_n1346), .B2(new_n1351), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1316), .B1(new_n1277), .B2(new_n1365), .ZN(new_n1366));
  XNOR2_X1  g1166(.A(new_n1366), .B(new_n1331), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1364), .A2(new_n1367), .ZN(new_n1368));
  XNOR2_X1  g1168(.A(new_n1366), .B(new_n1356), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1346), .A2(new_n1351), .A3(KEYINPUT127), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1368), .B1(new_n1371), .B2(new_n1364), .ZN(G402));
endmodule


