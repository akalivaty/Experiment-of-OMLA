

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n373, n374, n375, n376, n377, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773;

  XOR2_X1 U368 ( .A(KEYINPUT124), .B(n658), .Z(n659) );
  XNOR2_X1 U369 ( .A(n647), .B(KEYINPUT123), .ZN(n648) );
  OR2_X1 U370 ( .A1(n571), .A2(n435), .ZN(n357) );
  NOR2_X1 U371 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U372 ( .A1(n554), .A2(n625), .ZN(n555) );
  BUF_X1 U373 ( .A(n615), .Z(n348) );
  NOR2_X1 U374 ( .A1(n556), .A2(n548), .ZN(n549) );
  NOR2_X1 U375 ( .A1(n556), .A2(n542), .ZN(n729) );
  XNOR2_X1 U376 ( .A(n542), .B(KEYINPUT6), .ZN(n615) );
  NOR2_X1 U377 ( .A1(n718), .A2(n719), .ZN(n723) );
  XNOR2_X1 U378 ( .A(n532), .B(n349), .ZN(n658) );
  INV_X1 U379 ( .A(n524), .ZN(n350) );
  BUF_X1 U380 ( .A(G113), .Z(n356) );
  XNOR2_X1 U381 ( .A(n510), .B(n471), .ZN(n414) );
  XNOR2_X1 U382 ( .A(n473), .B(n472), .ZN(n424) );
  XNOR2_X1 U383 ( .A(n476), .B(KEYINPUT4), .ZN(n502) );
  XNOR2_X1 U384 ( .A(n351), .B(G125), .ZN(n479) );
  INV_X1 U385 ( .A(G146), .ZN(n351) );
  NOR2_X1 U386 ( .A1(n432), .A2(n575), .ZN(n366) );
  XNOR2_X2 U387 ( .A(n486), .B(KEYINPUT19), .ZN(n487) );
  XNOR2_X1 U388 ( .A(n438), .B(n437), .ZN(n678) );
  NAND2_X4 U389 ( .A1(n347), .A2(n374), .ZN(n352) );
  AND2_X2 U390 ( .A1(n369), .A2(n373), .ZN(n347) );
  XNOR2_X1 U391 ( .A(n754), .B(n350), .ZN(n349) );
  XNOR2_X2 U392 ( .A(n352), .B(KEYINPUT104), .ZN(n662) );
  NOR2_X1 U393 ( .A1(G953), .A2(G237), .ZN(n504) );
  XNOR2_X1 U394 ( .A(G143), .B(n356), .ZN(n449) );
  XNOR2_X1 U395 ( .A(n757), .B(G146), .ZN(n519) );
  NAND2_X2 U396 ( .A1(n391), .A2(n389), .ZN(n587) );
  NOR2_X1 U397 ( .A1(n717), .A2(n606), .ZN(n607) );
  XNOR2_X2 U398 ( .A(G143), .B(G128), .ZN(n478) );
  NAND2_X1 U399 ( .A1(n662), .A2(n544), .ZN(n545) );
  NOR2_X1 U400 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U401 ( .A1(n564), .A2(n563), .ZN(n603) );
  OR2_X1 U402 ( .A1(n714), .A2(n713), .ZN(n716) );
  NOR2_X1 U403 ( .A1(n371), .A2(n370), .ZN(n369) );
  XNOR2_X1 U404 ( .A(n404), .B(n503), .ZN(n757) );
  XNOR2_X1 U405 ( .A(n502), .B(n501), .ZN(n404) );
  XNOR2_X1 U406 ( .A(n478), .B(G134), .ZN(n503) );
  INV_X1 U407 ( .A(G110), .ZN(n472) );
  XNOR2_X1 U408 ( .A(G107), .B(G104), .ZN(n423) );
  XNOR2_X1 U409 ( .A(KEYINPUT73), .B(G131), .ZN(n501) );
  INV_X1 U410 ( .A(KEYINPUT36), .ZN(n618) );
  AND2_X1 U411 ( .A1(n672), .A2(n431), .ZN(n657) );
  AND2_X1 U412 ( .A1(n431), .A2(G475), .ZN(n666) );
  AND2_X1 U413 ( .A1(n431), .A2(G210), .ZN(n673) );
  AND2_X1 U414 ( .A1(n431), .A2(G472), .ZN(n663) );
  XNOR2_X2 U415 ( .A(n683), .B(n413), .ZN(n674) );
  XNOR2_X2 U416 ( .A(n414), .B(n517), .ZN(n683) );
  XNOR2_X1 U417 ( .A(n483), .B(n482), .ZN(n484) );
  INV_X1 U418 ( .A(n563), .ZN(n368) );
  XOR2_X1 U419 ( .A(KEYINPUT10), .B(n479), .Z(n754) );
  NAND2_X1 U420 ( .A1(n399), .A2(n398), .ZN(n397) );
  INV_X1 U421 ( .A(n592), .ZN(n398) );
  XNOR2_X1 U422 ( .A(n561), .B(n400), .ZN(n399) );
  INV_X1 U423 ( .A(KEYINPUT93), .ZN(n400) );
  INV_X1 U424 ( .A(KEYINPUT103), .ZN(n396) );
  INV_X1 U425 ( .A(KEYINPUT46), .ZN(n385) );
  INV_X1 U426 ( .A(G101), .ZN(n505) );
  XOR2_X1 U427 ( .A(KEYINPUT72), .B(KEYINPUT8), .Z(n463) );
  XNOR2_X1 U428 ( .A(G137), .B(G140), .ZN(n523) );
  NOR2_X1 U429 ( .A1(n429), .A2(n426), .ZN(n425) );
  INV_X1 U430 ( .A(n732), .ZN(n426) );
  NAND2_X1 U431 ( .A1(n722), .A2(n723), .ZN(n556) );
  NAND2_X1 U432 ( .A1(n665), .A2(n534), .ZN(n513) );
  XOR2_X1 U433 ( .A(KEYINPUT99), .B(G122), .Z(n457) );
  XNOR2_X1 U434 ( .A(G116), .B(G107), .ZN(n456) );
  XNOR2_X1 U435 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n458) );
  XOR2_X1 U436 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n459) );
  XNOR2_X1 U437 ( .A(n454), .B(n453), .ZN(n670) );
  XNOR2_X1 U438 ( .A(n754), .B(n447), .ZN(n454) );
  INV_X1 U439 ( .A(KEYINPUT89), .ZN(n514) );
  XNOR2_X1 U440 ( .A(n380), .B(KEYINPUT39), .ZN(n633) );
  NAND2_X1 U441 ( .A1(n381), .A2(n358), .ZN(n380) );
  INV_X1 U442 ( .A(n622), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n467), .B(n466), .ZN(n564) );
  AND2_X1 U444 ( .A1(n395), .A2(n688), .ZN(n568) );
  XNOR2_X1 U445 ( .A(n397), .B(n396), .ZN(n395) );
  XNOR2_X1 U446 ( .A(G122), .B(KEYINPUT12), .ZN(n448) );
  XNOR2_X1 U447 ( .A(KEYINPUT94), .B(KEYINPUT97), .ZN(n406) );
  AND2_X1 U448 ( .A1(n626), .A2(n360), .ZN(n383) );
  XOR2_X1 U449 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n527) );
  XOR2_X1 U450 ( .A(G140), .B(G104), .Z(n450) );
  XNOR2_X1 U451 ( .A(n408), .B(n405), .ZN(n452) );
  XNOR2_X1 U452 ( .A(n407), .B(n406), .ZN(n405) );
  XNOR2_X1 U453 ( .A(n409), .B(n448), .ZN(n408) );
  XNOR2_X1 U454 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n407) );
  INV_X1 U455 ( .A(KEYINPUT71), .ZN(n476) );
  NAND2_X1 U456 ( .A1(G234), .A2(G237), .ZN(n488) );
  INV_X1 U457 ( .A(G237), .ZN(n481) );
  AND2_X1 U458 ( .A1(n542), .A2(n621), .ZN(n543) );
  XNOR2_X1 U459 ( .A(n519), .B(n511), .ZN(n665) );
  INV_X1 U460 ( .A(KEYINPUT45), .ZN(n437) );
  NAND2_X1 U461 ( .A1(n366), .A2(n357), .ZN(n438) );
  NOR2_X1 U462 ( .A1(n735), .A2(n738), .ZN(n605) );
  XNOR2_X1 U463 ( .A(n455), .B(n411), .ZN(n410) );
  OR2_X1 U464 ( .A1(n670), .A2(G902), .ZN(n412) );
  INV_X1 U465 ( .A(G475), .ZN(n411) );
  NAND2_X1 U466 ( .A1(n388), .A2(n387), .ZN(n389) );
  AND2_X1 U467 ( .A1(n430), .A2(n390), .ZN(n387) );
  INV_X1 U468 ( .A(n718), .ZN(n370) );
  XNOR2_X1 U469 ( .A(KEYINPUT16), .B(G122), .ZN(n471) );
  XNOR2_X1 U470 ( .A(G128), .B(G119), .ZN(n530) );
  XNOR2_X1 U471 ( .A(n465), .B(n367), .ZN(n647) );
  XNOR2_X1 U472 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U473 ( .A(n519), .B(n520), .ZN(n653) );
  XNOR2_X1 U474 ( .A(n755), .B(n516), .ZN(n518) );
  XNOR2_X1 U475 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U476 ( .A(n379), .B(n604), .ZN(n768) );
  XNOR2_X1 U477 ( .A(n377), .B(KEYINPUT32), .ZN(n544) );
  INV_X1 U478 ( .A(KEYINPUT60), .ZN(n401) );
  INV_X1 U479 ( .A(KEYINPUT56), .ZN(n419) );
  AND2_X1 U480 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U481 ( .A1(n750), .A2(n761), .ZN(n751) );
  XNOR2_X1 U482 ( .A(KEYINPUT38), .B(n602), .ZN(n358) );
  AND2_X1 U483 ( .A1(n543), .A2(KEYINPUT65), .ZN(n359) );
  AND2_X1 U484 ( .A1(n595), .A2(n594), .ZN(n360) );
  INV_X1 U485 ( .A(n441), .ZN(n429) );
  NAND2_X1 U486 ( .A1(n484), .A2(n442), .ZN(n441) );
  AND2_X1 U487 ( .A1(n541), .A2(n540), .ZN(n361) );
  XOR2_X1 U488 ( .A(n665), .B(n664), .Z(n362) );
  XOR2_X1 U489 ( .A(n674), .B(n676), .Z(n363) );
  XOR2_X1 U490 ( .A(n670), .B(n669), .Z(n364) );
  NOR2_X1 U491 ( .A1(n761), .A2(G952), .ZN(n677) );
  XOR2_X1 U492 ( .A(KEYINPUT115), .B(KEYINPUT63), .Z(n365) );
  XNOR2_X1 U493 ( .A(n418), .B(n362), .ZN(n417) );
  INV_X1 U494 ( .A(n393), .ZN(n388) );
  NAND2_X1 U495 ( .A1(n427), .A2(n425), .ZN(n393) );
  XNOR2_X1 U496 ( .A(n464), .B(n503), .ZN(n367) );
  INV_X1 U497 ( .A(n564), .ZN(n553) );
  NAND2_X1 U498 ( .A1(n368), .A2(n564), .ZN(n735) );
  NAND2_X1 U499 ( .A1(n666), .A2(n672), .ZN(n403) );
  XNOR2_X2 U500 ( .A(n585), .B(KEYINPUT1), .ZN(n722) );
  NAND2_X1 U501 ( .A1(n663), .A2(n672), .ZN(n418) );
  NOR2_X1 U502 ( .A1(n543), .A2(KEYINPUT65), .ZN(n371) );
  NAND2_X1 U503 ( .A1(n565), .A2(n359), .ZN(n373) );
  NAND2_X1 U504 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U505 ( .A(KEYINPUT65), .ZN(n375) );
  INV_X1 U506 ( .A(n565), .ZN(n376) );
  XNOR2_X2 U507 ( .A(n500), .B(n499), .ZN(n565) );
  NAND2_X1 U508 ( .A1(n565), .A2(n361), .ZN(n377) );
  NAND2_X1 U509 ( .A1(n633), .A2(n612), .ZN(n379) );
  XNOR2_X1 U510 ( .A(n382), .B(n627), .ZN(n637) );
  NAND2_X1 U511 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U512 ( .A(n611), .B(n385), .ZN(n384) );
  INV_X1 U513 ( .A(n430), .ZN(n392) );
  NAND2_X1 U514 ( .A1(n386), .A2(n487), .ZN(n391) );
  NAND2_X1 U515 ( .A1(n388), .A2(n430), .ZN(n386) );
  OR2_X1 U516 ( .A1(n392), .A2(n393), .ZN(n616) );
  INV_X1 U517 ( .A(n487), .ZN(n390) );
  NAND2_X1 U518 ( .A1(n587), .A2(n493), .ZN(n495) );
  NAND2_X1 U519 ( .A1(n417), .A2(n671), .ZN(n416) );
  XNOR2_X1 U520 ( .A(n403), .B(n364), .ZN(n394) );
  NAND2_X1 U521 ( .A1(n394), .A2(n671), .ZN(n402) );
  AND2_X2 U522 ( .A1(n715), .A2(n646), .ZN(n672) );
  XNOR2_X1 U523 ( .A(n402), .B(n401), .ZN(G60) );
  NAND2_X1 U524 ( .A1(n729), .A2(n560), .ZN(n558) );
  NAND2_X1 U525 ( .A1(n504), .A2(G214), .ZN(n409) );
  XNOR2_X1 U526 ( .A(n420), .B(n419), .ZN(G51) );
  XNOR2_X2 U527 ( .A(n412), .B(n410), .ZN(n563) );
  NAND2_X1 U528 ( .A1(n674), .A2(n484), .ZN(n427) );
  XNOR2_X1 U529 ( .A(n415), .B(n480), .ZN(n413) );
  XNOR2_X2 U530 ( .A(n424), .B(n423), .ZN(n517) );
  XNOR2_X1 U531 ( .A(n477), .B(n502), .ZN(n415) );
  XNOR2_X1 U532 ( .A(n416), .B(n365), .ZN(G57) );
  NAND2_X2 U533 ( .A1(n643), .A2(n642), .ZN(n431) );
  INV_X4 U534 ( .A(G953), .ZN(n761) );
  NAND2_X1 U535 ( .A1(n428), .A2(n430), .ZN(n602) );
  XNOR2_X1 U536 ( .A(n422), .B(n363), .ZN(n421) );
  NAND2_X1 U537 ( .A1(n421), .A2(n671), .ZN(n420) );
  NAND2_X1 U538 ( .A1(n436), .A2(KEYINPUT81), .ZN(n435) );
  NAND2_X1 U539 ( .A1(n673), .A2(n672), .ZN(n422) );
  AND2_X1 U540 ( .A1(n427), .A2(n441), .ZN(n428) );
  OR2_X2 U541 ( .A1(n674), .A2(n440), .ZN(n430) );
  NAND2_X1 U542 ( .A1(n434), .A2(n433), .ZN(n432) );
  NAND2_X1 U543 ( .A1(n570), .A2(n439), .ZN(n433) );
  NAND2_X1 U544 ( .A1(n571), .A2(n439), .ZN(n434) );
  INV_X1 U545 ( .A(n570), .ZN(n436) );
  INV_X1 U546 ( .A(KEYINPUT81), .ZN(n439) );
  OR2_X1 U547 ( .A1(n484), .A2(n442), .ZN(n440) );
  INV_X1 U548 ( .A(n638), .ZN(n442) );
  XNOR2_X2 U549 ( .A(n444), .B(n443), .ZN(n510) );
  XNOR2_X2 U550 ( .A(G119), .B(KEYINPUT3), .ZN(n443) );
  XNOR2_X2 U551 ( .A(G116), .B(G113), .ZN(n444) );
  NOR2_X2 U552 ( .A1(n678), .A2(n759), .ZN(n712) );
  XNOR2_X1 U553 ( .A(n446), .B(KEYINPUT11), .ZN(n447) );
  XNOR2_X1 U554 ( .A(KEYINPUT74), .B(KEYINPUT48), .ZN(n627) );
  XNOR2_X1 U555 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U556 ( .A(n531), .B(n530), .ZN(n532) );
  OR2_X1 U557 ( .A1(n712), .A2(n711), .ZN(n714) );
  INV_X1 U558 ( .A(KEYINPUT34), .ZN(n551) );
  INV_X1 U559 ( .A(KEYINPUT0), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n552), .B(n551), .ZN(n554) );
  INV_X1 U561 ( .A(n677), .ZN(n671) );
  XOR2_X1 U562 ( .A(KEYINPUT35), .B(n555), .Z(n770) );
  INV_X1 U563 ( .A(n501), .ZN(n446) );
  XNOR2_X1 U564 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U565 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n455) );
  XNOR2_X1 U566 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U567 ( .A(n461), .B(n460), .Z(n465) );
  NAND2_X1 U568 ( .A1(G234), .A2(n761), .ZN(n462) );
  XNOR2_X1 U569 ( .A(n463), .B(n462), .ZN(n525) );
  NAND2_X1 U570 ( .A1(G217), .A2(n525), .ZN(n464) );
  INV_X1 U571 ( .A(G902), .ZN(n534) );
  NAND2_X1 U572 ( .A1(n647), .A2(n534), .ZN(n467) );
  INV_X1 U573 ( .A(G478), .ZN(n466) );
  XNOR2_X1 U574 ( .A(KEYINPUT15), .B(G902), .ZN(n638) );
  NAND2_X1 U575 ( .A1(n638), .A2(G234), .ZN(n468) );
  XNOR2_X1 U576 ( .A(n468), .B(KEYINPUT20), .ZN(n535) );
  AND2_X1 U577 ( .A1(n535), .A2(G221), .ZN(n470) );
  INV_X1 U578 ( .A(KEYINPUT21), .ZN(n469) );
  XNOR2_X1 U579 ( .A(n470), .B(n469), .ZN(n719) );
  NOR2_X1 U580 ( .A1(n735), .A2(n719), .ZN(n496) );
  XNOR2_X2 U581 ( .A(G101), .B(KEYINPUT84), .ZN(n473) );
  XNOR2_X1 U582 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n475) );
  NAND2_X1 U583 ( .A1(n761), .A2(G224), .ZN(n474) );
  XNOR2_X1 U584 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X1 U585 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U586 ( .A1(n534), .A2(n481), .ZN(n485) );
  NAND2_X1 U587 ( .A1(n485), .A2(G210), .ZN(n483) );
  INV_X1 U588 ( .A(KEYINPUT85), .ZN(n482) );
  NAND2_X1 U589 ( .A1(n485), .A2(G214), .ZN(n732) );
  INV_X1 U590 ( .A(KEYINPUT69), .ZN(n486) );
  XNOR2_X1 U591 ( .A(n488), .B(KEYINPUT86), .ZN(n489) );
  XNOR2_X1 U592 ( .A(KEYINPUT14), .B(n489), .ZN(n491) );
  AND2_X1 U593 ( .A1(n491), .A2(G902), .ZN(n576) );
  NOR2_X1 U594 ( .A1(G898), .A2(n761), .ZN(n684) );
  NAND2_X1 U595 ( .A1(n576), .A2(n684), .ZN(n490) );
  XNOR2_X1 U596 ( .A(n490), .B(KEYINPUT87), .ZN(n492) );
  NAND2_X1 U597 ( .A1(G952), .A2(n491), .ZN(n746) );
  NOR2_X1 U598 ( .A1(n746), .A2(G953), .ZN(n579) );
  OR2_X1 U599 ( .A1(n492), .A2(n579), .ZN(n493) );
  XNOR2_X2 U600 ( .A(n495), .B(n494), .ZN(n560) );
  NAND2_X1 U601 ( .A1(n496), .A2(n560), .ZN(n500) );
  XNOR2_X1 U602 ( .A(KEYINPUT76), .B(KEYINPUT22), .ZN(n498) );
  INV_X1 U603 ( .A(KEYINPUT66), .ZN(n497) );
  XNOR2_X1 U604 ( .A(n498), .B(n497), .ZN(n499) );
  NAND2_X1 U605 ( .A1(n504), .A2(G210), .ZN(n506) );
  XNOR2_X1 U606 ( .A(n506), .B(n505), .ZN(n508) );
  XOR2_X1 U607 ( .A(G137), .B(KEYINPUT5), .Z(n507) );
  XNOR2_X1 U608 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U609 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U610 ( .A(G472), .ZN(n512) );
  XNOR2_X2 U611 ( .A(n513), .B(n512), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n615), .B(KEYINPUT77), .ZN(n541) );
  XNOR2_X1 U613 ( .A(KEYINPUT88), .B(n523), .ZN(n755) );
  NAND2_X1 U614 ( .A1(G227), .A2(n761), .ZN(n515) );
  XNOR2_X1 U615 ( .A(n518), .B(n517), .ZN(n520) );
  NAND2_X1 U616 ( .A1(n653), .A2(n534), .ZN(n522) );
  XOR2_X1 U617 ( .A(KEYINPUT75), .B(G469), .Z(n521) );
  XNOR2_X2 U618 ( .A(n522), .B(n521), .ZN(n585) );
  INV_X1 U619 ( .A(n523), .ZN(n524) );
  NAND2_X1 U620 ( .A1(n525), .A2(G221), .ZN(n529) );
  XNOR2_X1 U621 ( .A(G110), .B(KEYINPUT90), .ZN(n526) );
  XNOR2_X1 U622 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U623 ( .A(n529), .B(n528), .ZN(n531) );
  NAND2_X1 U624 ( .A1(n658), .A2(n534), .ZN(n539) );
  XOR2_X1 U625 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n537) );
  NAND2_X1 U626 ( .A1(n535), .A2(G217), .ZN(n536) );
  XNOR2_X1 U627 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X2 U628 ( .A(n539), .B(n538), .ZN(n718) );
  AND2_X1 U629 ( .A1(n722), .A2(n718), .ZN(n540) );
  XNOR2_X1 U630 ( .A(n544), .B(G119), .ZN(G21) );
  INV_X1 U631 ( .A(n722), .ZN(n621) );
  XNOR2_X2 U632 ( .A(n545), .B(KEYINPUT82), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n572), .A2(KEYINPUT44), .ZN(n547) );
  INV_X1 U634 ( .A(KEYINPUT64), .ZN(n546) );
  XNOR2_X1 U635 ( .A(n547), .B(n546), .ZN(n571) );
  INV_X1 U636 ( .A(n615), .ZN(n548) );
  XNOR2_X1 U637 ( .A(n549), .B(KEYINPUT33), .ZN(n747) );
  INV_X1 U638 ( .A(n560), .ZN(n550) );
  NOR2_X1 U639 ( .A1(n747), .A2(n550), .ZN(n552) );
  NAND2_X1 U640 ( .A1(n553), .A2(n563), .ZN(n625) );
  NAND2_X1 U641 ( .A1(n770), .A2(KEYINPUT44), .ZN(n569) );
  XOR2_X1 U642 ( .A(KEYINPUT31), .B(KEYINPUT92), .Z(n557) );
  XNOR2_X2 U643 ( .A(n558), .B(n557), .ZN(n705) );
  NAND2_X1 U644 ( .A1(n585), .A2(n723), .ZN(n598) );
  NOR2_X1 U645 ( .A1(n581), .A2(n598), .ZN(n559) );
  NAND2_X1 U646 ( .A1(n560), .A2(n559), .ZN(n690) );
  NAND2_X1 U647 ( .A1(n705), .A2(n690), .ZN(n561) );
  NOR2_X1 U648 ( .A1(n564), .A2(n563), .ZN(n562) );
  XNOR2_X1 U649 ( .A(KEYINPUT102), .B(n562), .ZN(n694) );
  INV_X1 U650 ( .A(n694), .ZN(n706) );
  NAND2_X1 U651 ( .A1(n706), .A2(n603), .ZN(n589) );
  INV_X1 U652 ( .A(n589), .ZN(n737) );
  XNOR2_X1 U653 ( .A(KEYINPUT80), .B(n737), .ZN(n592) );
  AND2_X1 U654 ( .A1(n565), .A2(n621), .ZN(n567) );
  NOR2_X1 U655 ( .A1(n348), .A2(n718), .ZN(n566) );
  NAND2_X1 U656 ( .A1(n567), .A2(n566), .ZN(n688) );
  NAND2_X1 U657 ( .A1(n569), .A2(n568), .ZN(n570) );
  OR2_X1 U658 ( .A1(n770), .A2(KEYINPUT44), .ZN(n574) );
  BUF_X1 U659 ( .A(n572), .Z(n573) );
  NAND2_X1 U660 ( .A1(G953), .A2(n576), .ZN(n577) );
  NOR2_X1 U661 ( .A1(G900), .A2(n577), .ZN(n578) );
  NOR2_X1 U662 ( .A1(n579), .A2(n578), .ZN(n599) );
  NOR2_X1 U663 ( .A1(n719), .A2(n599), .ZN(n580) );
  NAND2_X1 U664 ( .A1(n718), .A2(n580), .ZN(n613) );
  INV_X1 U665 ( .A(n613), .ZN(n582) );
  INV_X1 U666 ( .A(n542), .ZN(n581) );
  NAND2_X1 U667 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U668 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n583) );
  XNOR2_X1 U669 ( .A(n584), .B(n583), .ZN(n586) );
  NAND2_X1 U670 ( .A1(n586), .A2(n585), .ZN(n606) );
  INV_X1 U671 ( .A(n587), .ZN(n588) );
  NOR2_X1 U672 ( .A1(n606), .A2(n588), .ZN(n701) );
  NAND2_X1 U673 ( .A1(n701), .A2(n589), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n590), .A2(KEYINPUT47), .ZN(n595) );
  XNOR2_X1 U675 ( .A(KEYINPUT70), .B(KEYINPUT47), .ZN(n591) );
  NOR2_X1 U676 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n593), .A2(n701), .ZN(n594) );
  XOR2_X1 U678 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n604) );
  NAND2_X1 U679 ( .A1(n581), .A2(n732), .ZN(n597) );
  XNOR2_X1 U680 ( .A(KEYINPUT30), .B(KEYINPUT107), .ZN(n596) );
  XNOR2_X1 U681 ( .A(n597), .B(n596), .ZN(n601) );
  NOR2_X1 U682 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U683 ( .A1(n601), .A2(n600), .ZN(n622) );
  INV_X1 U684 ( .A(n603), .ZN(n612) );
  INV_X1 U685 ( .A(n768), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n358), .A2(n732), .ZN(n738) );
  XNOR2_X1 U687 ( .A(KEYINPUT41), .B(n605), .ZN(n717) );
  XOR2_X1 U688 ( .A(KEYINPUT42), .B(n607), .Z(n608) );
  XNOR2_X1 U689 ( .A(KEYINPUT111), .B(n608), .ZN(n772) );
  INV_X1 U690 ( .A(n772), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U692 ( .A(KEYINPUT105), .B(n612), .Z(n700) );
  INV_X1 U693 ( .A(n700), .ZN(n703) );
  NOR2_X1 U694 ( .A1(n703), .A2(n613), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n348), .A2(n614), .ZN(n628) );
  XNOR2_X1 U696 ( .A(KEYINPUT112), .B(n628), .ZN(n617) );
  XNOR2_X1 U697 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n708) );
  NOR2_X1 U699 ( .A1(n622), .A2(n602), .ZN(n623) );
  XOR2_X1 U700 ( .A(KEYINPUT108), .B(n623), .Z(n624) );
  NOR2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n698) );
  NOR2_X1 U702 ( .A1(n708), .A2(n698), .ZN(n626) );
  NOR2_X1 U703 ( .A1(n722), .A2(n628), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n629), .A2(n732), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT43), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n631), .A2(n602), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n632), .B(KEYINPUT106), .ZN(n773) );
  NAND2_X1 U708 ( .A1(n633), .A2(n694), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(KEYINPUT113), .ZN(n771) );
  INV_X1 U710 ( .A(n771), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n773), .A2(n635), .ZN(n636) );
  OR2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n759) );
  INV_X1 U713 ( .A(n712), .ZN(n643) );
  NAND2_X1 U714 ( .A1(KEYINPUT2), .A2(KEYINPUT68), .ZN(n641) );
  NAND2_X1 U715 ( .A1(n442), .A2(KEYINPUT2), .ZN(n640) );
  INV_X1 U716 ( .A(KEYINPUT68), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n644) );
  AND2_X1 U718 ( .A1(n641), .A2(n644), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n712), .A2(KEYINPUT2), .ZN(n715) );
  INV_X1 U720 ( .A(n644), .ZN(n645) );
  OR2_X1 U721 ( .A1(n645), .A2(n442), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n657), .A2(G478), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X1 U724 ( .A1(n650), .A2(n677), .ZN(G63) );
  NAND2_X1 U725 ( .A1(n657), .A2(G469), .ZN(n655) );
  XOR2_X1 U726 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n651) );
  XNOR2_X1 U727 ( .A(n651), .B(KEYINPUT58), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X1 U730 ( .A1(n656), .A2(n677), .ZN(G54) );
  NAND2_X1 U731 ( .A1(n657), .A2(G217), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U733 ( .A1(n661), .A2(n677), .ZN(G66) );
  XNOR2_X1 U734 ( .A(n662), .B(G110), .ZN(G12) );
  XOR2_X1 U735 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n664) );
  XOR2_X1 U736 ( .A(KEYINPUT67), .B(KEYINPUT83), .Z(n668) );
  XNOR2_X1 U737 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U739 ( .A(KEYINPUT78), .B(KEYINPUT54), .ZN(n675) );
  XOR2_X1 U740 ( .A(n675), .B(KEYINPUT55), .Z(n676) );
  OR2_X1 U741 ( .A1(n678), .A2(G953), .ZN(n682) );
  NAND2_X1 U742 ( .A1(G953), .A2(G224), .ZN(n679) );
  XNOR2_X1 U743 ( .A(n679), .B(KEYINPUT61), .ZN(n680) );
  NAND2_X1 U744 ( .A1(n680), .A2(G898), .ZN(n681) );
  NAND2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n687) );
  INV_X1 U746 ( .A(n683), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U748 ( .A(n687), .B(n686), .ZN(G69) );
  XNOR2_X1 U749 ( .A(G101), .B(n688), .ZN(G3) );
  NOR2_X1 U750 ( .A1(n703), .A2(n690), .ZN(n689) );
  XOR2_X1 U751 ( .A(G104), .B(n689), .Z(G6) );
  NOR2_X1 U752 ( .A1(n706), .A2(n690), .ZN(n692) );
  XNOR2_X1 U753 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n691) );
  XNOR2_X1 U754 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U755 ( .A(G107), .B(n693), .ZN(G9) );
  XOR2_X1 U756 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n696) );
  NAND2_X1 U757 ( .A1(n701), .A2(n694), .ZN(n695) );
  XNOR2_X1 U758 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U759 ( .A(G128), .B(n697), .ZN(G30) );
  XNOR2_X1 U760 ( .A(G143), .B(n698), .ZN(n699) );
  XNOR2_X1 U761 ( .A(n699), .B(KEYINPUT117), .ZN(G45) );
  NAND2_X1 U762 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U763 ( .A(n702), .B(G146), .ZN(G48) );
  NOR2_X1 U764 ( .A1(n705), .A2(n703), .ZN(n704) );
  XOR2_X1 U765 ( .A(n356), .B(n704), .Z(G15) );
  NOR2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U767 ( .A(G116), .B(n707), .Z(G18) );
  XNOR2_X1 U768 ( .A(G125), .B(n708), .ZN(n709) );
  XNOR2_X1 U769 ( .A(n709), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U770 ( .A(KEYINPUT2), .ZN(n710) );
  AND2_X1 U771 ( .A1(n710), .A2(KEYINPUT79), .ZN(n711) );
  NOR2_X1 U772 ( .A1(n710), .A2(KEYINPUT79), .ZN(n713) );
  NAND2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n752) );
  NAND2_X1 U774 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U775 ( .A(KEYINPUT49), .B(n720), .Z(n721) );
  NAND2_X1 U776 ( .A1(n542), .A2(n721), .ZN(n726) );
  NOR2_X1 U777 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U778 ( .A(n724), .B(KEYINPUT50), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n727), .B(KEYINPUT118), .ZN(n728) );
  NOR2_X1 U781 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U782 ( .A(KEYINPUT51), .B(n730), .Z(n731) );
  NOR2_X1 U783 ( .A1(n717), .A2(n731), .ZN(n743) );
  NOR2_X1 U784 ( .A1(n358), .A2(n732), .ZN(n733) );
  XOR2_X1 U785 ( .A(KEYINPUT119), .B(n733), .Z(n734) );
  NOR2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U787 ( .A(n736), .B(KEYINPUT120), .ZN(n740) );
  NOR2_X1 U788 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U789 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U790 ( .A1(n741), .A2(n747), .ZN(n742) );
  NOR2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U792 ( .A(n744), .B(KEYINPUT52), .ZN(n745) );
  NOR2_X1 U793 ( .A1(n746), .A2(n745), .ZN(n749) );
  NOR2_X1 U794 ( .A1(n747), .A2(n717), .ZN(n748) );
  NOR2_X1 U795 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U796 ( .A(n753), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U797 ( .A(n755), .B(n754), .Z(n756) );
  XOR2_X1 U798 ( .A(n757), .B(n756), .Z(n763) );
  XOR2_X1 U799 ( .A(n763), .B(KEYINPUT125), .Z(n758) );
  XNOR2_X1 U800 ( .A(n759), .B(n758), .ZN(n760) );
  NAND2_X1 U801 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U802 ( .A(n762), .B(KEYINPUT126), .ZN(n767) );
  XNOR2_X1 U803 ( .A(G227), .B(n763), .ZN(n764) );
  NAND2_X1 U804 ( .A1(n764), .A2(G900), .ZN(n765) );
  NAND2_X1 U805 ( .A1(G953), .A2(n765), .ZN(n766) );
  NAND2_X1 U806 ( .A1(n767), .A2(n766), .ZN(G72) );
  XNOR2_X1 U807 ( .A(G131), .B(n768), .ZN(n769) );
  XNOR2_X1 U808 ( .A(n769), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U809 ( .A(n770), .B(G122), .Z(G24) );
  XOR2_X1 U810 ( .A(G134), .B(n771), .Z(G36) );
  XOR2_X1 U811 ( .A(G137), .B(n772), .Z(G39) );
  XNOR2_X1 U812 ( .A(G140), .B(n773), .ZN(G42) );
endmodule

