

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762;

  XNOR2_X1 U380 ( .A(G104), .B(G110), .ZN(n473) );
  XOR2_X1 U381 ( .A(G113), .B(G104), .Z(n422) );
  INV_X1 U382 ( .A(G146), .ZN(n455) );
  XNOR2_X1 U383 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n436) );
  XOR2_X1 U384 ( .A(KEYINPUT16), .B(G110), .Z(n402) );
  INV_X2 U385 ( .A(G128), .ZN(n391) );
  XNOR2_X1 U386 ( .A(G137), .B(G113), .ZN(n462) );
  XNOR2_X1 U387 ( .A(G110), .B(KEYINPUT96), .ZN(n481) );
  INV_X1 U388 ( .A(G902), .ZN(n468) );
  XNOR2_X1 U389 ( .A(G119), .B(KEYINPUT69), .ZN(n403) );
  XOR2_X1 U390 ( .A(G116), .B(KEYINPUT3), .Z(n404) );
  BUF_X1 U391 ( .A(G122), .Z(n760) );
  BUF_X1 U392 ( .A(G143), .Z(n705) );
  NOR2_X2 U393 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X2 U394 ( .A1(n367), .A2(n377), .ZN(n693) );
  AND2_X2 U395 ( .A1(n386), .A2(n382), .ZN(n367) );
  INV_X1 U396 ( .A(n709), .ZN(n707) );
  NOR2_X2 U397 ( .A1(n609), .A2(n707), .ZN(n626) );
  XNOR2_X1 U398 ( .A(n520), .B(KEYINPUT102), .ZN(n709) );
  INV_X1 U399 ( .A(KEYINPUT53), .ZN(n356) );
  XNOR2_X1 U400 ( .A(n660), .B(n356), .ZN(G75) );
  AND2_X1 U401 ( .A1(n523), .A2(n362), .ZN(n526) );
  NAND2_X1 U402 ( .A1(n384), .A2(n383), .ZN(n377) );
  NOR2_X1 U403 ( .A1(n637), .A2(n553), .ZN(n714) );
  XNOR2_X1 U404 ( .A(n506), .B(KEYINPUT33), .ZN(n630) );
  NOR2_X1 U405 ( .A1(n709), .A2(n548), .ZN(n599) );
  NOR2_X1 U406 ( .A1(n477), .A2(n387), .ZN(n383) );
  NOR2_X1 U407 ( .A1(n559), .A2(n558), .ZN(n584) );
  BUF_X1 U408 ( .A(n502), .Z(n637) );
  XNOR2_X1 U409 ( .A(n566), .B(KEYINPUT1), .ZN(n502) );
  XNOR2_X1 U410 ( .A(KEYINPUT75), .B(KEYINPUT93), .ZN(n395) );
  XNOR2_X2 U411 ( .A(G902), .B(KEYINPUT15), .ZN(n664) );
  XOR2_X2 U412 ( .A(G137), .B(G140), .Z(n479) );
  INV_X4 U413 ( .A(G953), .ZN(n750) );
  XNOR2_X2 U414 ( .A(G128), .B(G119), .ZN(n480) );
  NAND2_X1 U415 ( .A1(n718), .A2(G210), .ZN(n689) );
  NOR2_X2 U416 ( .A1(n666), .A2(n667), .ZN(n718) );
  BUF_X1 U417 ( .A(n560), .Z(n604) );
  XNOR2_X2 U418 ( .A(n514), .B(n371), .ZN(n516) );
  INV_X1 U419 ( .A(G237), .ZN(n407) );
  NOR2_X1 U420 ( .A1(G953), .A2(G237), .ZN(n458) );
  INV_X1 U421 ( .A(KEYINPUT65), .ZN(n387) );
  XNOR2_X1 U422 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n396) );
  INV_X1 U423 ( .A(KEYINPUT46), .ZN(n594) );
  XOR2_X1 U424 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n460) );
  INV_X1 U425 ( .A(n620), .ZN(n374) );
  INV_X1 U426 ( .A(KEYINPUT30), .ZN(n554) );
  AND2_X1 U427 ( .A1(n385), .A2(n495), .ZN(n382) );
  XNOR2_X1 U428 ( .A(n435), .B(n434), .ZN(n518) );
  INV_X1 U429 ( .A(KEYINPUT95), .ZN(n371) );
  INV_X1 U430 ( .A(n369), .ZN(n636) );
  XNOR2_X1 U431 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U432 ( .A(n685), .B(n687), .ZN(n688) );
  XNOR2_X1 U433 ( .A(n673), .B(KEYINPUT92), .ZN(n717) );
  NAND2_X1 U434 ( .A1(n498), .A2(KEYINPUT32), .ZN(n381) );
  NAND2_X1 U435 ( .A1(n380), .A2(n379), .ZN(n375) );
  NOR2_X1 U436 ( .A1(n498), .A2(KEYINPUT32), .ZN(n379) );
  XNOR2_X1 U437 ( .A(G107), .B(G122), .ZN(n440) );
  XNOR2_X1 U438 ( .A(n409), .B(n408), .ZN(n560) );
  NOR2_X1 U439 ( .A1(n560), .A2(n374), .ZN(n373) );
  NAND2_X1 U440 ( .A1(n364), .A2(n665), .ZN(n357) );
  NAND2_X1 U441 ( .A1(n364), .A2(n665), .ZN(n666) );
  NAND2_X1 U442 ( .A1(n406), .A2(n739), .ZN(n360) );
  NAND2_X1 U443 ( .A1(n358), .A2(n359), .ZN(n361) );
  NAND2_X1 U444 ( .A1(n360), .A2(n361), .ZN(n684) );
  INV_X1 U445 ( .A(n406), .ZN(n358) );
  INV_X1 U446 ( .A(n739), .ZN(n359) );
  XOR2_X2 U447 ( .A(n405), .B(n466), .Z(n739) );
  XNOR2_X1 U448 ( .A(n373), .B(KEYINPUT89), .ZN(n549) );
  AND2_X1 U449 ( .A1(n522), .A2(n695), .ZN(n362) );
  XNOR2_X2 U450 ( .A(n372), .B(KEYINPUT22), .ZN(n366) );
  BUF_X1 U451 ( .A(n443), .Z(n444) );
  NOR2_X1 U452 ( .A1(n667), .A2(n357), .ZN(n363) );
  OR2_X2 U453 ( .A1(n662), .A2(n613), .ZN(n364) );
  XNOR2_X1 U454 ( .A(n372), .B(KEYINPUT22), .ZN(n365) );
  NAND2_X2 U455 ( .A1(n501), .A2(n453), .ZN(n372) );
  XNOR2_X2 U456 ( .A(n503), .B(KEYINPUT71), .ZN(n513) );
  NOR2_X2 U457 ( .A1(n502), .A2(n638), .ZN(n503) );
  NAND2_X1 U458 ( .A1(n376), .A2(n375), .ZN(n368) );
  NAND2_X1 U459 ( .A1(n376), .A2(n375), .ZN(n762) );
  AND2_X2 U460 ( .A1(n378), .A2(n381), .ZN(n376) );
  XNOR2_X2 U461 ( .A(n469), .B(G472), .ZN(n369) );
  NOR2_X2 U462 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U463 ( .A(n595), .B(n594), .ZN(n596) );
  BUF_X1 U464 ( .A(n630), .Z(n370) );
  NAND2_X1 U465 ( .A1(n693), .A2(n762), .ZN(n499) );
  NAND2_X1 U466 ( .A1(n366), .A2(KEYINPUT32), .ZN(n378) );
  INV_X1 U467 ( .A(n366), .ZN(n380) );
  INV_X1 U468 ( .A(n365), .ZN(n384) );
  NAND2_X1 U469 ( .A1(n477), .A2(n387), .ZN(n385) );
  NAND2_X1 U470 ( .A1(n366), .A2(n387), .ZN(n386) );
  NOR2_X1 U471 ( .A1(n663), .A2(KEYINPUT2), .ZN(n667) );
  BUF_X1 U472 ( .A(n662), .Z(n733) );
  XOR2_X1 U473 ( .A(KEYINPUT40), .B(KEYINPUT114), .Z(n388) );
  XOR2_X1 U474 ( .A(n473), .B(n472), .Z(n389) );
  XOR2_X1 U475 ( .A(G113), .B(G104), .Z(n390) );
  INV_X1 U476 ( .A(KEYINPUT72), .ZN(n461) );
  XNOR2_X1 U477 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U478 ( .A(n454), .B(n399), .ZN(n406) );
  XNOR2_X1 U479 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U480 ( .A(n661), .ZN(n607) );
  BUF_X1 U481 ( .A(n744), .Z(n746) );
  XNOR2_X1 U482 ( .A(n587), .B(n388), .ZN(n588) );
  XNOR2_X1 U483 ( .A(n586), .B(n585), .ZN(n610) );
  XNOR2_X2 U484 ( .A(G143), .B(KEYINPUT78), .ZN(n392) );
  XNOR2_X2 U485 ( .A(n392), .B(n391), .ZN(n443) );
  XNOR2_X2 U486 ( .A(n443), .B(KEYINPUT4), .ZN(n744) );
  XNOR2_X2 U487 ( .A(n744), .B(G101), .ZN(n454) );
  XNOR2_X1 U488 ( .A(G125), .B(G146), .ZN(n421) );
  NAND2_X1 U489 ( .A1(n750), .A2(G224), .ZN(n393) );
  XNOR2_X1 U490 ( .A(n393), .B(KEYINPUT94), .ZN(n394) );
  XNOR2_X1 U491 ( .A(n421), .B(n394), .ZN(n398) );
  XNOR2_X1 U492 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U493 ( .A(n398), .B(n397), .ZN(n399) );
  INV_X1 U494 ( .A(n440), .ZN(n400) );
  XNOR2_X1 U495 ( .A(n390), .B(n400), .ZN(n401) );
  XNOR2_X1 U496 ( .A(n402), .B(n401), .ZN(n405) );
  XNOR2_X1 U497 ( .A(n404), .B(n403), .ZN(n466) );
  NAND2_X1 U498 ( .A1(n684), .A2(n664), .ZN(n409) );
  NAND2_X1 U499 ( .A1(n468), .A2(n407), .ZN(n410) );
  NAND2_X1 U500 ( .A1(n410), .A2(G210), .ZN(n408) );
  NAND2_X1 U501 ( .A1(n410), .A2(G214), .ZN(n620) );
  XNOR2_X1 U502 ( .A(KEYINPUT73), .B(KEYINPUT19), .ZN(n411) );
  XNOR2_X1 U503 ( .A(n549), .B(n411), .ZN(n572) );
  NOR2_X1 U504 ( .A1(G898), .A2(n750), .ZN(n741) );
  NAND2_X1 U505 ( .A1(n741), .A2(G902), .ZN(n412) );
  NAND2_X1 U506 ( .A1(n750), .A2(G952), .ZN(n541) );
  NAND2_X1 U507 ( .A1(n412), .A2(n541), .ZN(n416) );
  NAND2_X1 U508 ( .A1(G237), .A2(G234), .ZN(n414) );
  INV_X1 U509 ( .A(KEYINPUT14), .ZN(n413) );
  XNOR2_X1 U510 ( .A(n414), .B(n413), .ZN(n653) );
  INV_X1 U511 ( .A(n653), .ZN(n415) );
  NAND2_X1 U512 ( .A1(n416), .A2(n415), .ZN(n417) );
  OR2_X2 U513 ( .A1(n572), .A2(n417), .ZN(n420) );
  INV_X1 U514 ( .A(KEYINPUT66), .ZN(n418) );
  XNOR2_X1 U515 ( .A(n418), .B(KEYINPUT0), .ZN(n419) );
  XNOR2_X2 U516 ( .A(n420), .B(n419), .ZN(n501) );
  XNOR2_X1 U517 ( .A(KEYINPUT13), .B(G475), .ZN(n435) );
  XOR2_X1 U518 ( .A(KEYINPUT10), .B(n421), .Z(n478) );
  INV_X1 U519 ( .A(n478), .ZN(n423) );
  XOR2_X1 U520 ( .A(n423), .B(n422), .Z(n425) );
  XNOR2_X1 U521 ( .A(n705), .B(G131), .ZN(n424) );
  XNOR2_X1 U522 ( .A(n425), .B(n424), .ZN(n433) );
  XOR2_X1 U523 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n427) );
  XNOR2_X1 U524 ( .A(n760), .B(G140), .ZN(n426) );
  XNOR2_X1 U525 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U526 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n429) );
  NAND2_X1 U527 ( .A1(G214), .A2(n458), .ZN(n428) );
  XNOR2_X1 U528 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U529 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U530 ( .A(n433), .B(n432), .ZN(n669) );
  NOR2_X1 U531 ( .A1(G902), .A2(n669), .ZN(n434) );
  XOR2_X1 U532 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n439) );
  NAND2_X1 U533 ( .A1(n750), .A2(G234), .ZN(n437) );
  XNOR2_X1 U534 ( .A(n437), .B(n436), .ZN(n485) );
  NAND2_X1 U535 ( .A1(G217), .A2(n485), .ZN(n438) );
  XNOR2_X1 U536 ( .A(n439), .B(n438), .ZN(n442) );
  XOR2_X1 U537 ( .A(n400), .B(G116), .Z(n441) );
  XNOR2_X1 U538 ( .A(n442), .B(n441), .ZN(n446) );
  XNOR2_X1 U539 ( .A(n444), .B(G134), .ZN(n445) );
  XNOR2_X1 U540 ( .A(n446), .B(n445), .ZN(n725) );
  NOR2_X1 U541 ( .A1(G902), .A2(n725), .ZN(n447) );
  XNOR2_X1 U542 ( .A(G478), .B(n447), .ZN(n519) );
  INV_X1 U543 ( .A(n519), .ZN(n509) );
  NOR2_X1 U544 ( .A1(n518), .A2(n509), .ZN(n448) );
  XNOR2_X1 U545 ( .A(n448), .B(KEYINPUT105), .ZN(n623) );
  NAND2_X1 U546 ( .A1(G234), .A2(n664), .ZN(n449) );
  XNOR2_X1 U547 ( .A(KEYINPUT20), .B(n449), .ZN(n489) );
  AND2_X1 U548 ( .A1(n489), .A2(G221), .ZN(n451) );
  XNOR2_X1 U549 ( .A(KEYINPUT98), .B(KEYINPUT21), .ZN(n450) );
  XNOR2_X1 U550 ( .A(n451), .B(n450), .ZN(n633) );
  INV_X1 U551 ( .A(n633), .ZN(n452) );
  NOR2_X1 U552 ( .A1(n623), .A2(n452), .ZN(n453) );
  BUF_X2 U553 ( .A(n454), .Z(n457) );
  XNOR2_X1 U554 ( .A(G131), .B(G134), .ZN(n745) );
  XNOR2_X1 U555 ( .A(n745), .B(n455), .ZN(n456) );
  XNOR2_X2 U556 ( .A(n457), .B(n456), .ZN(n474) );
  NAND2_X1 U557 ( .A1(n458), .A2(G210), .ZN(n459) );
  XNOR2_X1 U558 ( .A(n460), .B(n459), .ZN(n464) );
  XNOR2_X1 U559 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U560 ( .A(n474), .B(n467), .ZN(n679) );
  NAND2_X1 U561 ( .A1(n679), .A2(n468), .ZN(n469) );
  XOR2_X1 U562 ( .A(G107), .B(n479), .Z(n471) );
  NAND2_X1 U563 ( .A1(G227), .A2(n750), .ZN(n470) );
  XNOR2_X1 U564 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U565 ( .A(n474), .B(n389), .ZN(n719) );
  NOR2_X1 U566 ( .A1(G902), .A2(n719), .ZN(n476) );
  XNOR2_X1 U567 ( .A(KEYINPUT68), .B(G469), .ZN(n475) );
  XNOR2_X2 U568 ( .A(n476), .B(n475), .ZN(n566) );
  INV_X1 U569 ( .A(n637), .ZN(n601) );
  OR2_X1 U570 ( .A1(n369), .A2(n601), .ZN(n477) );
  XNOR2_X1 U571 ( .A(n479), .B(n478), .ZN(n748) );
  XNOR2_X1 U572 ( .A(n480), .B(KEYINPUT23), .ZN(n484) );
  XOR2_X1 U573 ( .A(KEYINPUT24), .B(KEYINPUT82), .Z(n482) );
  XNOR2_X1 U574 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U575 ( .A(n484), .B(n483), .Z(n487) );
  NAND2_X1 U576 ( .A1(G221), .A2(n485), .ZN(n486) );
  XNOR2_X1 U577 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U578 ( .A(n748), .B(n488), .ZN(n728) );
  NOR2_X1 U579 ( .A1(n728), .A2(G902), .ZN(n494) );
  XOR2_X1 U580 ( .A(KEYINPUT74), .B(KEYINPUT97), .Z(n491) );
  NAND2_X1 U581 ( .A1(G217), .A2(n489), .ZN(n490) );
  XNOR2_X1 U582 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U583 ( .A(n492), .B(KEYINPUT25), .ZN(n493) );
  XNOR2_X1 U584 ( .A(n494), .B(n493), .ZN(n544) );
  INV_X1 U585 ( .A(n544), .ZN(n495) );
  XNOR2_X1 U586 ( .A(n544), .B(KEYINPUT106), .ZN(n632) );
  XNOR2_X1 U587 ( .A(n369), .B(KEYINPUT6), .ZN(n496) );
  XNOR2_X1 U588 ( .A(n496), .B(KEYINPUT104), .ZN(n546) );
  INV_X1 U589 ( .A(n546), .ZN(n504) );
  NOR2_X1 U590 ( .A1(n632), .A2(n504), .ZN(n497) );
  NAND2_X1 U591 ( .A1(n601), .A2(n497), .ZN(n498) );
  XNOR2_X1 U592 ( .A(n499), .B(KEYINPUT88), .ZN(n529) );
  NAND2_X1 U593 ( .A1(n529), .A2(KEYINPUT44), .ZN(n500) );
  XNOR2_X1 U594 ( .A(n500), .B(KEYINPUT64), .ZN(n527) );
  BUF_X2 U595 ( .A(n501), .Z(n514) );
  NAND2_X1 U596 ( .A1(n544), .A2(n633), .ZN(n638) );
  XNOR2_X1 U597 ( .A(n513), .B(KEYINPUT107), .ZN(n505) );
  NAND2_X1 U598 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U599 ( .A1(n516), .A2(n630), .ZN(n508) );
  XOR2_X1 U600 ( .A(KEYINPUT34), .B(KEYINPUT76), .Z(n507) );
  XNOR2_X1 U601 ( .A(n508), .B(n507), .ZN(n511) );
  NAND2_X1 U602 ( .A1(n518), .A2(n509), .ZN(n561) );
  INV_X1 U603 ( .A(n561), .ZN(n510) );
  NAND2_X1 U604 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X2 U605 ( .A(n512), .B(KEYINPUT35), .ZN(n761) );
  NAND2_X1 U606 ( .A1(n761), .A2(KEYINPUT44), .ZN(n523) );
  NOR2_X1 U607 ( .A1(n636), .A2(n513), .ZN(n643) );
  NAND2_X1 U608 ( .A1(n643), .A2(n514), .ZN(n515) );
  XOR2_X1 U609 ( .A(KEYINPUT31), .B(n515), .Z(n711) );
  NOR2_X1 U610 ( .A1(n566), .A2(n638), .ZN(n556) );
  AND2_X1 U611 ( .A1(n516), .A2(n636), .ZN(n517) );
  NAND2_X1 U612 ( .A1(n556), .A2(n517), .ZN(n697) );
  NAND2_X1 U613 ( .A1(n711), .A2(n697), .ZN(n521) );
  NOR2_X1 U614 ( .A1(n518), .A2(n519), .ZN(n701) );
  XOR2_X1 U615 ( .A(KEYINPUT103), .B(n701), .Z(n609) );
  NAND2_X1 U616 ( .A1(n519), .A2(n518), .ZN(n520) );
  INV_X1 U617 ( .A(n626), .ZN(n578) );
  NAND2_X1 U618 ( .A1(n521), .A2(n578), .ZN(n522) );
  NOR2_X1 U619 ( .A1(n365), .A2(n601), .ZN(n525) );
  AND2_X1 U620 ( .A1(n546), .A2(n632), .ZN(n524) );
  NAND2_X1 U621 ( .A1(n525), .A2(n524), .ZN(n695) );
  NAND2_X1 U622 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U623 ( .A(n528), .B(KEYINPUT87), .ZN(n535) );
  BUF_X1 U624 ( .A(n529), .Z(n530) );
  INV_X1 U625 ( .A(n530), .ZN(n532) );
  NOR2_X1 U626 ( .A1(n761), .A2(KEYINPUT44), .ZN(n531) );
  NAND2_X1 U627 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U628 ( .A(n533), .B(KEYINPUT70), .ZN(n534) );
  NAND2_X1 U629 ( .A1(n535), .A2(n534), .ZN(n537) );
  XOR2_X1 U630 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n536) );
  XNOR2_X2 U631 ( .A(n537), .B(n536), .ZN(n662) );
  NAND2_X1 U632 ( .A1(G953), .A2(G902), .ZN(n538) );
  NOR2_X1 U633 ( .A1(n653), .A2(n538), .ZN(n539) );
  XOR2_X1 U634 ( .A(KEYINPUT108), .B(n539), .Z(n540) );
  NOR2_X1 U635 ( .A1(G900), .A2(n540), .ZN(n543) );
  NOR2_X1 U636 ( .A1(n653), .A2(n541), .ZN(n542) );
  NOR2_X1 U637 ( .A1(n543), .A2(n542), .ZN(n559) );
  NOR2_X1 U638 ( .A1(n544), .A2(n559), .ZN(n545) );
  NAND2_X1 U639 ( .A1(n633), .A2(n545), .ZN(n567) );
  NOR2_X1 U640 ( .A1(n546), .A2(n567), .ZN(n547) );
  XNOR2_X1 U641 ( .A(n547), .B(KEYINPUT109), .ZN(n548) );
  INV_X1 U642 ( .A(n599), .ZN(n551) );
  BUF_X1 U643 ( .A(n549), .Z(n550) );
  XOR2_X1 U644 ( .A(KEYINPUT36), .B(n552), .Z(n553) );
  XNOR2_X1 U645 ( .A(KEYINPUT85), .B(n714), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n369), .A2(n620), .ZN(n555) );
  XNOR2_X1 U647 ( .A(n555), .B(n554), .ZN(n557) );
  NAND2_X1 U648 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U649 ( .A1(n604), .A2(n561), .ZN(n562) );
  AND2_X1 U650 ( .A1(n584), .A2(n562), .ZN(n704) );
  NAND2_X1 U651 ( .A1(n626), .A2(KEYINPUT47), .ZN(n563) );
  XNOR2_X1 U652 ( .A(KEYINPUT81), .B(n563), .ZN(n564) );
  NOR2_X1 U653 ( .A1(n704), .A2(n564), .ZN(n565) );
  XNOR2_X1 U654 ( .A(n565), .B(KEYINPUT80), .ZN(n577) );
  XNOR2_X1 U655 ( .A(n566), .B(KEYINPUT111), .ZN(n571) );
  NOR2_X1 U656 ( .A1(n636), .A2(n567), .ZN(n569) );
  XNOR2_X1 U657 ( .A(KEYINPUT112), .B(KEYINPUT28), .ZN(n568) );
  XNOR2_X1 U658 ( .A(n569), .B(n568), .ZN(n570) );
  AND2_X1 U659 ( .A1(n571), .A2(n570), .ZN(n591) );
  INV_X1 U660 ( .A(n591), .ZN(n573) );
  OR2_X1 U661 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U662 ( .A(n574), .B(KEYINPUT77), .ZN(n706) );
  INV_X1 U663 ( .A(n706), .ZN(n575) );
  NAND2_X1 U664 ( .A1(KEYINPUT47), .A2(n575), .ZN(n576) );
  NAND2_X1 U665 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U666 ( .A1(n706), .A2(n578), .ZN(n579) );
  NOR2_X1 U667 ( .A1(KEYINPUT47), .A2(n579), .ZN(n580) );
  NOR2_X1 U668 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U669 ( .A1(n583), .A2(n582), .ZN(n597) );
  XNOR2_X1 U670 ( .A(n604), .B(KEYINPUT38), .ZN(n621) );
  NAND2_X1 U671 ( .A1(n584), .A2(n621), .ZN(n586) );
  XNOR2_X1 U672 ( .A(KEYINPUT86), .B(KEYINPUT39), .ZN(n585) );
  NAND2_X1 U673 ( .A1(n610), .A2(n707), .ZN(n587) );
  XOR2_X1 U674 ( .A(KEYINPUT113), .B(n588), .Z(n758) );
  NAND2_X1 U675 ( .A1(n621), .A2(n620), .ZN(n625) );
  NOR2_X1 U676 ( .A1(n623), .A2(n625), .ZN(n590) );
  XNOR2_X1 U677 ( .A(KEYINPUT41), .B(KEYINPUT115), .ZN(n589) );
  XNOR2_X1 U678 ( .A(n590), .B(n589), .ZN(n645) );
  NAND2_X1 U679 ( .A1(n645), .A2(n591), .ZN(n592) );
  XOR2_X1 U680 ( .A(KEYINPUT42), .B(n592), .Z(n593) );
  XNOR2_X1 U681 ( .A(KEYINPUT116), .B(n593), .ZN(n757) );
  NOR2_X1 U682 ( .A1(n758), .A2(n757), .ZN(n595) );
  XNOR2_X1 U683 ( .A(n598), .B(KEYINPUT48), .ZN(n608) );
  XNOR2_X1 U684 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n603) );
  NAND2_X1 U685 ( .A1(n599), .A2(n620), .ZN(n600) );
  NOR2_X1 U686 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U687 ( .A(n603), .B(n602), .ZN(n606) );
  INV_X1 U688 ( .A(n604), .ZN(n605) );
  NOR2_X1 U689 ( .A1(n606), .A2(n605), .ZN(n661) );
  AND2_X2 U690 ( .A1(n608), .A2(n607), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n716) );
  NAND2_X1 U692 ( .A1(n716), .A2(KEYINPUT2), .ZN(n611) );
  XNOR2_X1 U693 ( .A(n611), .B(KEYINPUT79), .ZN(n612) );
  NAND2_X1 U694 ( .A1(n614), .A2(n612), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n614), .A2(n716), .ZN(n749) );
  INV_X1 U696 ( .A(KEYINPUT2), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n749), .A2(n616), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n364), .A2(n615), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n733), .A2(n616), .ZN(n617) );
  XNOR2_X1 U700 ( .A(n617), .B(KEYINPUT83), .ZN(n618) );
  NOR2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n658) );
  NAND2_X1 U702 ( .A1(n370), .A2(n645), .ZN(n656) );
  NOR2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U705 ( .A(KEYINPUT119), .B(n624), .Z(n628) );
  NOR2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U708 ( .A(KEYINPUT120), .B(n629), .Z(n631) );
  NAND2_X1 U709 ( .A1(n631), .A2(n370), .ZN(n649) );
  NOR2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n634), .B(KEYINPUT49), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n641) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U714 ( .A(KEYINPUT50), .B(n639), .Z(n640) );
  NOR2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U717 ( .A(KEYINPUT51), .B(n644), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U719 ( .A(KEYINPUT118), .B(n647), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(KEYINPUT121), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n651), .B(KEYINPUT52), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n654), .A2(G952), .ZN(n655) );
  NAND2_X1 U725 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U727 ( .A1(n750), .A2(n659), .ZN(n660) );
  XOR2_X1 U728 ( .A(G140), .B(n661), .Z(G42) );
  NOR2_X1 U729 ( .A1(n662), .A2(n749), .ZN(n663) );
  INV_X1 U730 ( .A(n664), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n718), .A2(G475), .ZN(n671) );
  XNOR2_X1 U732 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n671), .B(n670), .ZN(n674) );
  INV_X1 U734 ( .A(G952), .ZN(n672) );
  NAND2_X1 U735 ( .A1(n672), .A2(G953), .ZN(n673) );
  NAND2_X1 U736 ( .A1(n674), .A2(n717), .ZN(n676) );
  XNOR2_X1 U737 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n675) );
  XNOR2_X1 U738 ( .A(n676), .B(n675), .ZN(G60) );
  NAND2_X1 U739 ( .A1(n718), .A2(G472), .ZN(n681) );
  XNOR2_X1 U740 ( .A(KEYINPUT91), .B(KEYINPUT117), .ZN(n677) );
  XNOR2_X1 U741 ( .A(n677), .B(KEYINPUT62), .ZN(n678) );
  XNOR2_X1 U742 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U743 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U744 ( .A1(n682), .A2(n717), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n683), .B(KEYINPUT63), .ZN(G57) );
  BUF_X1 U746 ( .A(n684), .Z(n685) );
  XNOR2_X1 U747 ( .A(KEYINPUT90), .B(KEYINPUT54), .ZN(n686) );
  XOR2_X1 U748 ( .A(n686), .B(KEYINPUT55), .Z(n687) );
  XNOR2_X1 U749 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U750 ( .A1(n690), .A2(n717), .ZN(n692) );
  XOR2_X1 U751 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n691) );
  XNOR2_X1 U752 ( .A(n692), .B(n691), .ZN(G51) );
  BUF_X1 U753 ( .A(n693), .Z(n694) );
  XNOR2_X1 U754 ( .A(n694), .B(G110), .ZN(G12) );
  XNOR2_X1 U755 ( .A(G101), .B(n695), .ZN(G3) );
  NOR2_X1 U756 ( .A1(n709), .A2(n697), .ZN(n696) );
  XOR2_X1 U757 ( .A(G104), .B(n696), .Z(G6) );
  INV_X1 U758 ( .A(n701), .ZN(n712) );
  NOR2_X1 U759 ( .A1(n712), .A2(n697), .ZN(n699) );
  XNOR2_X1 U760 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U762 ( .A(G107), .B(n700), .ZN(G9) );
  XOR2_X1 U763 ( .A(G128), .B(KEYINPUT29), .Z(n703) );
  NAND2_X1 U764 ( .A1(n706), .A2(n701), .ZN(n702) );
  XNOR2_X1 U765 ( .A(n703), .B(n702), .ZN(G30) );
  XOR2_X1 U766 ( .A(n705), .B(n704), .Z(G45) );
  NAND2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U768 ( .A(n708), .B(G146), .ZN(G48) );
  NOR2_X1 U769 ( .A1(n709), .A2(n711), .ZN(n710) );
  XOR2_X1 U770 ( .A(G113), .B(n710), .Z(G15) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U772 ( .A(G116), .B(n713), .Z(G18) );
  XNOR2_X1 U773 ( .A(G125), .B(n714), .ZN(n715) );
  XNOR2_X1 U774 ( .A(n715), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U775 ( .A(G134), .B(n716), .ZN(G36) );
  INV_X1 U776 ( .A(n717), .ZN(n731) );
  NAND2_X1 U777 ( .A1(n363), .A2(G469), .ZN(n723) );
  XNOR2_X1 U778 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n721) );
  XNOR2_X1 U779 ( .A(n719), .B(KEYINPUT57), .ZN(n720) );
  XNOR2_X1 U780 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U781 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U782 ( .A1(n731), .A2(n724), .ZN(G54) );
  NAND2_X1 U783 ( .A1(n363), .A2(G478), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U785 ( .A1(n731), .A2(n727), .ZN(G63) );
  NAND2_X1 U786 ( .A1(n363), .A2(G217), .ZN(n730) );
  XNOR2_X1 U787 ( .A(n728), .B(KEYINPUT126), .ZN(n729) );
  XNOR2_X1 U788 ( .A(n730), .B(n729), .ZN(n732) );
  NOR2_X1 U789 ( .A1(n732), .A2(n731), .ZN(G66) );
  INV_X1 U790 ( .A(n733), .ZN(n734) );
  NAND2_X1 U791 ( .A1(n734), .A2(n750), .ZN(n738) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n735) );
  XNOR2_X1 U793 ( .A(KEYINPUT61), .B(n735), .ZN(n736) );
  NAND2_X1 U794 ( .A1(n736), .A2(G898), .ZN(n737) );
  NAND2_X1 U795 ( .A1(n738), .A2(n737), .ZN(n743) );
  XNOR2_X1 U796 ( .A(n739), .B(G101), .ZN(n740) );
  NOR2_X1 U797 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U798 ( .A(n743), .B(n742), .ZN(G69) );
  XNOR2_X1 U799 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U800 ( .A(n748), .B(n747), .ZN(n752) );
  XNOR2_X1 U801 ( .A(n752), .B(n749), .ZN(n751) );
  NAND2_X1 U802 ( .A1(n751), .A2(n750), .ZN(n756) );
  XNOR2_X1 U803 ( .A(G227), .B(n752), .ZN(n753) );
  NAND2_X1 U804 ( .A1(n753), .A2(G900), .ZN(n754) );
  NAND2_X1 U805 ( .A1(G953), .A2(n754), .ZN(n755) );
  NAND2_X1 U806 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U807 ( .A(G137), .B(n757), .Z(G39) );
  XNOR2_X1 U808 ( .A(G131), .B(n758), .ZN(n759) );
  XNOR2_X1 U809 ( .A(n759), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U810 ( .A(n761), .B(n760), .Z(G24) );
  XNOR2_X1 U811 ( .A(G119), .B(n368), .ZN(G21) );
endmodule

