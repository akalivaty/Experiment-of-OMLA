//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G101), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  INV_X1    g014(.A(G116), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G119), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G116), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n200), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT2), .B(G113), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(G116), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n201), .A2(G119), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT68), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n206), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n202), .A2(new_n204), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n198), .A2(new_n199), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n197), .A2(KEYINPUT74), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n191), .A2(new_n194), .A3(new_n216), .A4(new_n195), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n196), .A2(new_n219), .A3(G101), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n215), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n206), .A2(new_n202), .A3(new_n204), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT68), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT68), .B1(new_n207), .B2(new_n208), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT5), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G113), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT5), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(new_n202), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n222), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n190), .A2(G107), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n193), .A2(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n217), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n214), .A2(new_n221), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n189), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n225), .A2(new_n228), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n213), .A3(new_n233), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n215), .A2(new_n218), .A3(new_n220), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n210), .A2(new_n213), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n196), .A2(G101), .A3(new_n199), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n238), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n235), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G143), .ZN(new_n248));
  INV_X1    g062(.A(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G146), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n248), .A2(new_n250), .A3(new_n251), .A4(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n249), .A2(G146), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n247), .B2(G143), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n249), .A2(KEYINPUT64), .A3(G146), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n248), .B2(KEYINPUT1), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n252), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  OR2_X1    g074(.A1(new_n260), .A2(G125), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT0), .B(G128), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n248), .A2(new_n250), .ZN(new_n264));
  OAI22_X1  g078(.A1(new_n257), .A2(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G125), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G224), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT79), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n214), .A2(new_n221), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n235), .B1(new_n272), .B2(new_n238), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n271), .B1(new_n273), .B2(new_n189), .ZN(new_n274));
  NOR4_X1   g088(.A1(new_n234), .A2(KEYINPUT79), .A3(KEYINPUT6), .A4(new_n235), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n246), .B(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n243), .A2(new_n189), .A3(new_n244), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT79), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n271), .A3(new_n189), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n282), .A2(KEYINPUT80), .A3(new_n246), .A4(new_n270), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n234), .A2(new_n235), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n235), .B(KEYINPUT81), .ZN(new_n286));
  XOR2_X1   g100(.A(new_n286), .B(KEYINPUT8), .Z(new_n287));
  INV_X1    g101(.A(new_n233), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n229), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n212), .A2(KEYINPUT5), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n222), .B1(new_n228), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n287), .B(new_n289), .C1(new_n288), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n269), .A2(KEYINPUT7), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT82), .A2(KEYINPUT7), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n267), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n267), .B2(new_n294), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n285), .B(new_n292), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n284), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n284), .A2(new_n302), .A3(new_n300), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n188), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT83), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT18), .A2(G131), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(G237), .A2(G953), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n311), .A2(G143), .A3(G214), .ZN(new_n312));
  AOI21_X1  g126(.A(G143), .B1(new_n311), .B2(G214), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(G214), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n249), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n311), .A2(G143), .A3(G214), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n309), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G125), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G140), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n247), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n323), .A3(new_n247), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT72), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n321), .A2(new_n323), .A3(new_n327), .A4(new_n247), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n324), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT84), .B1(new_n319), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n324), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n327), .B1(new_n332), .B2(new_n247), .ZN(new_n333));
  AND4_X1   g147(.A1(new_n327), .A2(new_n321), .A3(new_n323), .A4(new_n247), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n318), .A4(new_n314), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT16), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G146), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(G146), .B1(new_n339), .B2(new_n340), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G131), .B1(new_n312), .B2(new_n313), .ZN(new_n345));
  INV_X1    g159(.A(G131), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n316), .A2(new_n346), .A3(new_n317), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT17), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n344), .B(new_n349), .C1(new_n348), .C2(new_n345), .ZN(new_n350));
  XNOR2_X1  g164(.A(G113), .B(G122), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(new_n190), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n338), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n332), .A2(KEYINPUT19), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n332), .A2(KEYINPUT19), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n247), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n341), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(new_n345), .B2(new_n347), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n345), .A2(new_n347), .A3(new_n358), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n360), .A2(new_n361), .B1(new_n330), .B2(new_n337), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n353), .B1(new_n362), .B2(new_n352), .ZN(new_n363));
  NOR3_X1   g177(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT86), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n338), .A2(new_n352), .A3(new_n350), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n345), .A2(new_n347), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT85), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n369), .A2(new_n341), .A3(new_n361), .A4(new_n356), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n352), .B1(new_n338), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n366), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(G475), .A2(G902), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n353), .B(KEYINPUT86), .C1(new_n362), .C2(new_n352), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n365), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G475), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n352), .B1(new_n338), .B2(new_n350), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n367), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n379), .B1(new_n381), .B2(new_n298), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  INV_X1    g199(.A(G217), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n385), .A2(new_n386), .A3(G953), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n249), .A2(G128), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n258), .A2(G143), .ZN(new_n390));
  INV_X1    g204(.A(G134), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G116), .B(G122), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(new_n193), .ZN(new_n394));
  INV_X1    g208(.A(G122), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G116), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n201), .A2(G122), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n396), .A2(new_n397), .A3(new_n193), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n392), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT13), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT87), .B1(new_n389), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT87), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n402), .A2(new_n249), .A3(KEYINPUT13), .A4(G128), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n389), .A2(new_n400), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n401), .A2(new_n403), .A3(new_n390), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n399), .B1(G134), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n393), .A2(new_n193), .ZN(new_n407));
  INV_X1    g221(.A(new_n392), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n391), .B1(new_n389), .B2(new_n390), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n411));
  OAI21_X1  g225(.A(G107), .B1(new_n397), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n411), .B2(new_n393), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n388), .B1(new_n406), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n405), .A2(G134), .ZN(new_n416));
  OAI221_X1 g230(.A(new_n387), .B1(new_n413), .B2(new_n410), .C1(new_n416), .C2(new_n399), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT88), .B(new_n388), .C1(new_n406), .C2(new_n414), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n298), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G478), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(KEYINPUT15), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n423), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n419), .A2(new_n298), .A3(new_n420), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT89), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n424), .A2(KEYINPUT89), .A3(new_n426), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n268), .A2(G952), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(G234), .B2(G237), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n298), .B(new_n268), .C1(G234), .C2(G237), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(G898), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(new_n430), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n384), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  INV_X1    g254(.A(G227), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G953), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n440), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n233), .A2(new_n260), .A3(KEYINPUT10), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n233), .A2(new_n260), .A3(KEYINPUT76), .A4(KEYINPUT10), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n196), .A2(G101), .A3(new_n199), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(new_n265), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT10), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n248), .A2(KEYINPUT1), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n453), .A2(G128), .B1(new_n248), .B2(new_n250), .ZN(new_n454));
  INV_X1    g268(.A(new_n252), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n217), .B(new_n232), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n221), .A2(new_n451), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G137), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT65), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G137), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT11), .A4(G134), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT66), .B1(new_n459), .B2(G134), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n391), .A3(G137), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n459), .A2(G134), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT11), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G131), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n463), .A2(new_n467), .A3(new_n346), .A4(new_n470), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n458), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT78), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT78), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n458), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n474), .B(KEYINPUT77), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n458), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n444), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n458), .A2(new_n480), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n456), .B1(new_n260), .B2(new_n233), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n484), .A2(KEYINPUT12), .A3(new_n474), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT12), .B1(new_n484), .B2(new_n474), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n483), .A2(new_n487), .A3(new_n443), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n439), .B(new_n298), .C1(new_n482), .C2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n477), .B1(new_n458), .B2(new_n474), .ZN(new_n490));
  INV_X1    g304(.A(new_n474), .ZN(new_n491));
  AOI211_X1 g305(.A(KEYINPUT78), .B(new_n491), .C1(new_n449), .C2(new_n457), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n481), .B(new_n444), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n443), .B1(new_n483), .B2(new_n487), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(G469), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n439), .A2(new_n298), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n489), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G221), .B1(new_n385), .B2(G902), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n438), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n326), .A2(new_n328), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n203), .A2(G128), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT23), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT71), .B1(new_n258), .B2(G119), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(G110), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT24), .B(G110), .Z(new_n507));
  NAND2_X1  g321(.A1(new_n258), .A2(G119), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n502), .A2(new_n508), .A3(KEYINPUT70), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n341), .B(new_n501), .C1(new_n506), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n505), .A2(G110), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(new_n512), .A3(new_n507), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n515), .B(new_n516), .C1(new_n343), .C2(new_n342), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n517), .A3(new_n521), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n298), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n523), .A2(KEYINPUT25), .A3(new_n298), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n386), .B1(G234), .B2(new_n298), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n524), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n530), .A2(G902), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT73), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT32), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n311), .A2(G210), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT27), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT69), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n265), .B1(new_n472), .B2(new_n473), .ZN(new_n548));
  AOI21_X1  g362(.A(G134), .B1(new_n460), .B2(new_n462), .ZN(new_n549));
  INV_X1    g363(.A(new_n468), .ZN(new_n550));
  OAI21_X1  g364(.A(G131), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n260), .A2(new_n473), .A3(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n548), .A2(new_n552), .A3(new_n240), .ZN(new_n553));
  INV_X1    g367(.A(new_n240), .ZN(new_n554));
  INV_X1    g368(.A(new_n265), .ZN(new_n555));
  INV_X1    g369(.A(new_n473), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n464), .A2(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n346), .B1(new_n557), .B2(new_n463), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n555), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n260), .A2(new_n473), .A3(new_n551), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT28), .B1(new_n553), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n554), .A3(new_n560), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT28), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n547), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT30), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n567), .A2(KEYINPUT67), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(KEYINPUT67), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n569), .C1(new_n548), .C2(new_n552), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n559), .A2(KEYINPUT67), .A3(new_n567), .A4(new_n560), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n240), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n563), .A3(new_n545), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n566), .B1(new_n574), .B2(KEYINPUT31), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n553), .B1(new_n572), .B2(new_n240), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT31), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n577), .A3(new_n545), .ZN(new_n578));
  AOI211_X1 g392(.A(new_n539), .B(new_n541), .C1(new_n575), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(KEYINPUT31), .ZN(new_n580));
  INV_X1    g394(.A(new_n566), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT32), .B1(new_n582), .B2(new_n540), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n576), .A2(new_n545), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT29), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n562), .A2(new_n565), .ZN(new_n587));
  INV_X1    g401(.A(new_n547), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n562), .A2(new_n565), .A3(KEYINPUT29), .A4(new_n545), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n585), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G472), .B1(new_n591), .B2(G902), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n538), .B1(new_n584), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n302), .B1(new_n284), .B2(new_n300), .ZN(new_n594));
  AOI211_X1 g408(.A(new_n303), .B(new_n299), .C1(new_n278), .C2(new_n283), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n187), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT83), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n308), .A2(new_n500), .A3(new_n593), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT90), .B(G101), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G3));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n582), .B2(new_n298), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT91), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT91), .B1(new_n582), .B2(new_n540), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n604), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n498), .A2(new_n499), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n606), .A2(new_n607), .A3(new_n538), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n419), .A2(new_n609), .A3(new_n420), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n415), .A2(new_n417), .A3(KEYINPUT33), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(G478), .A3(new_n298), .A4(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n421), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(G478), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n375), .A2(KEYINPUT20), .B1(new_n363), .B2(new_n364), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n436), .B(new_n614), .C1(new_n615), .C2(new_n382), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n596), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n608), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  AOI21_X1  g434(.A(new_n382), .B1(new_n429), .B2(new_n430), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n375), .A2(KEYINPUT92), .A3(KEYINPUT20), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT92), .B1(new_n375), .B2(KEYINPUT20), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n372), .A2(new_n374), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT93), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n625), .A2(new_n626), .A3(new_n377), .A4(new_n373), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT93), .B1(new_n375), .B2(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n436), .B(new_n621), .C1(new_n624), .C2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT94), .B1(new_n631), .B2(new_n306), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT94), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n596), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n608), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  NOR2_X1   g451(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n518), .B(new_n638), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n529), .A2(new_n530), .B1(new_n536), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n604), .B(new_n641), .C1(new_n602), .C2(new_n605), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n643), .A2(new_n308), .A3(new_n500), .A4(new_n597), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  AOI21_X1  g460(.A(new_n640), .B1(new_n584), .B2(new_n592), .ZN(new_n647));
  INV_X1    g461(.A(new_n607), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n628), .B(new_n627), .C1(new_n622), .C2(new_n623), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n433), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n432), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n649), .A2(new_n621), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n647), .A2(new_n648), .A3(new_n655), .A4(new_n306), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  XNOR2_X1  g471(.A(new_n653), .B(KEYINPUT39), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n594), .A2(new_n595), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT38), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n378), .A2(new_n383), .B1(new_n429), .B2(new_n430), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n664), .A2(new_n187), .A3(new_n640), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n577), .B1(new_n576), .B2(new_n545), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n554), .B1(new_n570), .B2(new_n571), .ZN(new_n667));
  INV_X1    g481(.A(new_n545), .ZN(new_n668));
  NOR4_X1   g482(.A1(new_n667), .A2(KEYINPUT31), .A3(new_n553), .A4(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n666), .A2(new_n669), .A3(new_n566), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n539), .B1(new_n670), .B2(new_n541), .ZN(new_n671));
  INV_X1    g485(.A(new_n574), .ZN(new_n672));
  INV_X1    g486(.A(new_n561), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n547), .B1(new_n563), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n298), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G472), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n582), .A2(KEYINPUT32), .A3(new_n540), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n671), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n665), .A2(new_n678), .ZN(new_n679));
  OR3_X1    g493(.A1(new_n663), .A2(KEYINPUT95), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT95), .B1(new_n663), .B2(new_n679), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n661), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NAND3_X1  g497(.A1(new_n384), .A2(new_n614), .A3(new_n653), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n647), .A2(new_n648), .A3(new_n306), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  OAI21_X1  g501(.A(new_n481), .B1(new_n490), .B2(new_n492), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n488), .B1(new_n688), .B2(new_n443), .ZN(new_n689));
  OAI21_X1  g503(.A(G469), .B1(new_n689), .B2(G902), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n489), .A2(new_n690), .A3(new_n499), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n617), .A2(new_n593), .A3(KEYINPUT96), .A4(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT96), .ZN(new_n693));
  INV_X1    g507(.A(new_n538), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n671), .A2(new_n592), .A3(new_n677), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n616), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n697), .B(new_n187), .C1(new_n594), .C2(new_n595), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n693), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n692), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  INV_X1    g516(.A(new_n696), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n703), .B1(new_n632), .B2(new_n634), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  AND3_X1   g519(.A1(new_n695), .A2(new_n438), .A3(new_n641), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n489), .A2(new_n690), .A3(new_n499), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n596), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  OAI211_X1 g524(.A(new_n664), .B(new_n187), .C1(new_n594), .C2(new_n595), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n489), .A2(new_n690), .A3(new_n436), .A4(new_n499), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n580), .A2(new_n581), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(KEYINPUT97), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n669), .B1(new_n714), .B2(KEYINPUT97), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n541), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n717), .A2(new_n538), .A3(new_n602), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NOR3_X1   g534(.A1(new_n717), .A2(new_n602), .A3(new_n640), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n708), .A3(new_n685), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  INV_X1    g538(.A(new_n499), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n689), .A2(G902), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n496), .B1(new_n726), .B2(new_n439), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT98), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n493), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n493), .A2(new_n728), .ZN(new_n730));
  OAI211_X1 g544(.A(G469), .B(new_n494), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n725), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n594), .A2(new_n595), .A3(new_n188), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n593), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n724), .B1(new_n734), .B2(new_n684), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n593), .A4(new_n685), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT99), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n735), .A2(new_n737), .A3(KEYINPUT99), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT100), .B(G131), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G33));
  NAND3_X1  g558(.A1(new_n736), .A2(new_n593), .A3(new_n655), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  NOR2_X1   g560(.A1(new_n615), .A2(new_n382), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n747), .A2(new_n748), .A3(new_n614), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n747), .B2(new_n614), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n749), .A2(new_n750), .A3(new_n640), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(KEYINPUT44), .A3(new_n606), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT101), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n733), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT44), .B1(new_n751), .B2(new_n606), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n755), .B1(new_n756), .B2(KEYINPUT102), .ZN(new_n757));
  OAI211_X1 g571(.A(KEYINPUT45), .B(new_n494), .C1(new_n729), .C2(new_n730), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT45), .B1(new_n493), .B2(new_n494), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n439), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n496), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n489), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n499), .B(new_n658), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n756), .A2(KEYINPUT102), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n754), .A2(new_n757), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  NOR4_X1   g582(.A1(new_n755), .A2(new_n694), .A3(new_n695), .A4(new_n684), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT103), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n499), .B1(new_n762), .B2(new_n763), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT47), .B(new_n499), .C1(new_n762), .C2(new_n763), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  NAND3_X1  g591(.A1(new_n663), .A2(new_n188), .A3(new_n691), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n749), .A2(new_n750), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n718), .A2(new_n432), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT113), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n755), .A2(new_n784), .A3(new_n707), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT114), .B1(new_n733), .B2(new_n691), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n785), .A2(new_n652), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n678), .A2(new_n538), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n384), .A2(new_n614), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n721), .A3(new_n779), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT113), .B(KEYINPUT50), .C1(new_n778), .C2(new_n780), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n783), .A2(new_n790), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n489), .A2(new_n690), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT104), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n489), .A2(new_n690), .A3(KEYINPUT104), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n725), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n773), .A2(new_n774), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n780), .A2(new_n755), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n795), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n780), .A2(new_n596), .A3(new_n707), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n431), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n787), .A2(new_n788), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n384), .A2(new_n614), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT116), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n787), .A2(new_n593), .A3(new_n779), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT48), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT48), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n787), .A2(new_n816), .A3(new_n593), .A4(new_n779), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n813), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n801), .A2(new_n805), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n794), .B1(new_n793), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n807), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n807), .A2(new_n821), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n713), .A2(new_n718), .B1(new_n706), .B2(new_n708), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n700), .A2(new_n704), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n700), .A2(new_n704), .A3(new_n829), .A4(KEYINPUT111), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n738), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT112), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n721), .A2(new_n685), .A3(new_n732), .A4(new_n733), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n654), .B2(new_n734), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n647), .A2(new_n648), .ZN(new_n838));
  INV_X1    g652(.A(new_n427), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n383), .A2(new_n839), .A3(new_n653), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n649), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT106), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n649), .A2(new_n840), .A3(KEYINPUT106), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n733), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n837), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n608), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n811), .B1(new_n839), .B2(new_n384), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n308), .A2(new_n597), .A3(new_n436), .A4(new_n849), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n644), .A2(new_n598), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n847), .A2(KEYINPUT110), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT110), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n745), .B(new_n836), .C1(new_n838), .C2(new_n845), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n598), .B(new_n644), .C1(new_n848), .C2(new_n850), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n639), .A2(new_n536), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n653), .B(KEYINPUT107), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n531), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT108), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n640), .A2(KEYINPUT108), .A3(new_n860), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n865), .A2(new_n678), .ZN(new_n866));
  INV_X1    g680(.A(new_n711), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT109), .A4(new_n732), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT109), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n731), .A2(new_n489), .A3(new_n497), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n865), .A2(new_n870), .A3(new_n499), .A4(new_n678), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n871), .B2(new_n711), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n656), .A2(new_n686), .A3(new_n722), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT52), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n656), .A2(new_n686), .A3(new_n722), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n868), .A2(new_n872), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n656), .A2(new_n722), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n881), .B2(KEYINPUT52), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n875), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n832), .A2(new_n884), .A3(new_n738), .A4(new_n833), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n835), .A2(new_n858), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n830), .A2(new_n856), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n740), .A3(new_n741), .A4(new_n847), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n875), .A2(new_n879), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n880), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n891), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT53), .B1(new_n881), .B2(KEYINPUT52), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n889), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n892), .B1(new_n896), .B2(new_n887), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n828), .A2(new_n897), .B1(G952), .B2(G953), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n798), .A2(new_n799), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(KEYINPUT49), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n694), .A2(new_n187), .A3(new_n499), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n747), .A2(new_n614), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n678), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(KEYINPUT49), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n900), .A2(new_n663), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT105), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n898), .A2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n268), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(G210), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n910), .B(new_n298), .C1(new_n886), .C2(new_n891), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n282), .A2(new_n246), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n270), .ZN(new_n913));
  XOR2_X1   g727(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n915), .A2(KEYINPUT56), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n909), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n886), .A2(new_n891), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(G210), .A3(G902), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT119), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n298), .B1(new_n886), .B2(new_n891), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n923), .A3(G210), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n917), .B1(new_n925), .B2(new_n915), .ZN(G51));
  XNOR2_X1  g740(.A(new_n496), .B(KEYINPUT57), .ZN(new_n927));
  INV_X1    g741(.A(new_n892), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n887), .B1(new_n886), .B2(new_n891), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n689), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n922), .A2(new_n758), .A3(new_n760), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n908), .B1(new_n932), .B2(new_n933), .ZN(G54));
  AND2_X1   g748(.A1(KEYINPUT58), .A2(G475), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n922), .A2(new_n625), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n625), .B1(new_n922), .B2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n908), .ZN(G60));
  AND2_X1   g752(.A1(new_n610), .A2(new_n611), .ZN(new_n939));
  XOR2_X1   g753(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n940));
  NOR2_X1   g754(.A1(new_n422), .A2(new_n298), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n939), .B(new_n942), .C1(new_n928), .C2(new_n929), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n909), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n939), .B1(new_n897), .B2(new_n942), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(G63));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n886), .B2(new_n891), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n639), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n909), .B1(new_n950), .B2(new_n533), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n947), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n950), .A2(new_n533), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(KEYINPUT61), .A3(new_n909), .A4(new_n951), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(G66));
  INV_X1    g771(.A(G224), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n434), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n888), .B(KEYINPUT121), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(G953), .ZN(new_n961));
  INV_X1    g775(.A(new_n912), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(G898), .B2(new_n268), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT122), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n961), .B(new_n964), .ZN(G69));
  OR2_X1    g779(.A1(new_n354), .A2(new_n355), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n572), .B(new_n966), .Z(new_n967));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n682), .A2(new_n968), .A3(new_n876), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n593), .A2(new_n733), .A3(new_n849), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n970), .A2(new_n659), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n969), .A2(new_n767), .A3(new_n776), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n682), .A2(new_n876), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT123), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n973), .A2(new_n976), .A3(KEYINPUT62), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n972), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n967), .B1(new_n978), .B2(G953), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n740), .A2(new_n741), .A3(new_n745), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n980), .A2(KEYINPUT124), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n867), .A2(new_n593), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n874), .B1(new_n765), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n776), .A2(new_n767), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n980), .A2(KEYINPUT124), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n967), .A2(G953), .ZN(new_n987));
  AOI22_X1  g801(.A1(new_n986), .A2(new_n987), .B1(new_n650), .B2(G953), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n979), .A2(new_n988), .ZN(new_n989));
  OAI221_X1 g803(.A(G953), .B1(new_n441), .B2(new_n650), .C1(new_n967), .C2(KEYINPUT125), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT126), .Z(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n989), .B(new_n992), .ZN(G72));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n978), .B2(new_n960), .ZN(new_n997));
  INV_X1    g811(.A(new_n576), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n545), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n995), .B1(new_n672), .B2(new_n585), .ZN(new_n1000));
  OAI22_X1  g814(.A1(new_n997), .A2(new_n999), .B1(new_n896), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n998), .A2(new_n545), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n960), .A2(new_n981), .A3(new_n984), .A4(new_n985), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n995), .ZN(new_n1005));
  OR3_X1    g819(.A1(new_n1005), .A2(KEYINPUT127), .A3(new_n908), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT127), .B1(new_n1005), .B2(new_n908), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(G57));
endmodule


