

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(n694), .A2(n689), .ZN(n691) );
  BUF_X1 U552 ( .A(n537), .Z(n518) );
  XNOR2_X1 U553 ( .A(n522), .B(KEYINPUT17), .ZN(n523) );
  XNOR2_X1 U554 ( .A(n524), .B(n523), .ZN(n537) );
  XNOR2_X1 U555 ( .A(KEYINPUT65), .B(G2104), .ZN(n527) );
  NOR2_X1 U556 ( .A1(n527), .A2(G2105), .ZN(n528) );
  NOR2_X1 U557 ( .A1(n534), .A2(n533), .ZN(G160) );
  OR2_X1 U558 ( .A1(n762), .A2(KEYINPUT33), .ZN(n519) );
  AND2_X1 U559 ( .A1(n981), .A2(n829), .ZN(n520) );
  OR2_X1 U560 ( .A1(n783), .A2(n782), .ZN(n521) );
  INV_X1 U561 ( .A(KEYINPUT26), .ZN(n690) );
  INV_X1 U562 ( .A(KEYINPUT98), .ZN(n699) );
  NOR2_X1 U563 ( .A1(n706), .A2(n705), .ZN(n713) );
  XNOR2_X1 U564 ( .A(KEYINPUT29), .B(KEYINPUT100), .ZN(n718) );
  INV_X1 U565 ( .A(n983), .ZN(n768) );
  NOR2_X1 U566 ( .A1(n769), .A2(n768), .ZN(n770) );
  INV_X1 U567 ( .A(KEYINPUT68), .ZN(n522) );
  NOR2_X1 U568 ( .A1(n817), .A2(n520), .ZN(n818) );
  NOR2_X1 U569 ( .A1(G651), .A2(G543), .ZN(n647) );
  XNOR2_X1 U570 ( .A(n544), .B(KEYINPUT88), .ZN(G164) );
  AND2_X1 U571 ( .A1(n527), .A2(G2105), .ZN(n883) );
  NAND2_X1 U572 ( .A1(G125), .A2(n883), .ZN(n526) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  NAND2_X1 U574 ( .A1(G137), .A2(n518), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n534) );
  XNOR2_X1 U576 ( .A(n528), .B(KEYINPUT66), .ZN(n614) );
  NAND2_X1 U577 ( .A1(n614), .A2(G101), .ZN(n529) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n529), .Z(n532) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n882) );
  NAND2_X1 U580 ( .A1(G113), .A2(n882), .ZN(n530) );
  XOR2_X1 U581 ( .A(KEYINPUT67), .B(n530), .Z(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U583 ( .A1(G114), .A2(n882), .ZN(n536) );
  NAND2_X1 U584 ( .A1(G126), .A2(n883), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n543) );
  NAND2_X1 U586 ( .A1(G138), .A2(n537), .ZN(n539) );
  NAND2_X1 U587 ( .A1(G102), .A2(n614), .ZN(n538) );
  NAND2_X1 U588 ( .A1(n539), .A2(n538), .ZN(n541) );
  INV_X1 U589 ( .A(KEYINPUT87), .ZN(n540) );
  XNOR2_X1 U590 ( .A(n541), .B(n540), .ZN(n542) );
  NOR2_X1 U591 ( .A1(n543), .A2(n542), .ZN(n544) );
  INV_X1 U592 ( .A(G651), .ZN(n548) );
  NOR2_X1 U593 ( .A1(G543), .A2(n548), .ZN(n545) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n545), .Z(n646) );
  NAND2_X1 U595 ( .A1(G65), .A2(n646), .ZN(n547) );
  NAND2_X1 U596 ( .A1(G91), .A2(n647), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n547), .A2(n546), .ZN(n553) );
  XOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .Z(n631) );
  NOR2_X1 U599 ( .A1(n631), .A2(n548), .ZN(n650) );
  NAND2_X1 U600 ( .A1(G78), .A2(n650), .ZN(n551) );
  NOR2_X1 U601 ( .A1(G651), .A2(n631), .ZN(n549) );
  XNOR2_X1 U602 ( .A(KEYINPUT64), .B(n549), .ZN(n654) );
  NAND2_X1 U603 ( .A1(G53), .A2(n654), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n552) );
  OR2_X1 U605 ( .A1(n553), .A2(n552), .ZN(G299) );
  AND2_X1 U606 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U607 ( .A(G132), .ZN(G219) );
  INV_X1 U608 ( .A(G120), .ZN(G236) );
  INV_X1 U609 ( .A(G69), .ZN(G235) );
  INV_X1 U610 ( .A(G108), .ZN(G238) );
  NAND2_X1 U611 ( .A1(n650), .A2(G77), .ZN(n554) );
  XNOR2_X1 U612 ( .A(n554), .B(KEYINPUT70), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G90), .A2(n647), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U615 ( .A(n557), .B(KEYINPUT9), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G64), .A2(n646), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G52), .A2(n654), .ZN(n560) );
  XNOR2_X1 U619 ( .A(KEYINPUT69), .B(n560), .ZN(n561) );
  NOR2_X1 U620 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U621 ( .A1(n647), .A2(G89), .ZN(n563) );
  XNOR2_X1 U622 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U623 ( .A1(G76), .A2(n650), .ZN(n564) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U625 ( .A(n566), .B(KEYINPUT5), .ZN(n573) );
  XNOR2_X1 U626 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n571) );
  NAND2_X1 U627 ( .A1(n646), .A2(G63), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT76), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G51), .A2(n654), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U633 ( .A(KEYINPUT7), .B(n574), .ZN(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U636 ( .A(n575), .B(KEYINPUT72), .ZN(n576) );
  XNOR2_X1 U637 ( .A(KEYINPUT10), .B(n576), .ZN(G223) );
  XNOR2_X1 U638 ( .A(KEYINPUT73), .B(G223), .ZN(n834) );
  NAND2_X1 U639 ( .A1(n834), .A2(G567), .ZN(n577) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  NAND2_X1 U641 ( .A1(G56), .A2(n646), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(n578), .Z(n584) );
  NAND2_X1 U643 ( .A1(n647), .A2(G81), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G68), .A2(n650), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(n582), .Z(n583) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G43), .A2(n654), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n975) );
  INV_X1 U651 ( .A(G860), .ZN(n601) );
  OR2_X1 U652 ( .A1(n975), .A2(n601), .ZN(G153) );
  INV_X1 U653 ( .A(G171), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G301), .A2(G868), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT74), .ZN(n597) );
  NAND2_X1 U656 ( .A1(n654), .A2(G54), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G92), .A2(n647), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G79), .A2(n650), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G66), .A2(n646), .ZN(n590) );
  XNOR2_X1 U661 ( .A(KEYINPUT75), .B(n590), .ZN(n591) );
  NOR2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U664 ( .A(n595), .B(KEYINPUT15), .ZN(n686) );
  BUF_X1 U665 ( .A(n686), .Z(n982) );
  OR2_X1 U666 ( .A1(G868), .A2(n982), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(G284) );
  INV_X1 U668 ( .A(G868), .ZN(n665) );
  XNOR2_X1 U669 ( .A(KEYINPUT78), .B(n665), .ZN(n598) );
  NOR2_X1 U670 ( .A1(G286), .A2(n598), .ZN(n600) );
  NOR2_X1 U671 ( .A1(G868), .A2(G299), .ZN(n599) );
  NOR2_X1 U672 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U673 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n602), .A2(n982), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT16), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT79), .B(n604), .Z(G148) );
  NAND2_X1 U677 ( .A1(n982), .A2(G868), .ZN(n605) );
  NOR2_X1 U678 ( .A1(G559), .A2(n605), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT80), .ZN(n608) );
  NOR2_X1 U680 ( .A1(n975), .A2(G868), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G111), .A2(n882), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G135), .A2(n518), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n883), .A2(G123), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT18), .B(n611), .Z(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n616) );
  BUF_X1 U688 ( .A(n614), .Z(n887) );
  NAND2_X1 U689 ( .A1(G99), .A2(n887), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n956) );
  XOR2_X1 U691 ( .A(n956), .B(G2096), .Z(n618) );
  XNOR2_X1 U692 ( .A(G2100), .B(KEYINPUT81), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(KEYINPUT82), .B(n619), .ZN(G156) );
  NAND2_X1 U695 ( .A1(n982), .A2(G559), .ZN(n663) );
  XNOR2_X1 U696 ( .A(n975), .B(n663), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n620), .A2(G860), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G67), .A2(n646), .ZN(n622) );
  NAND2_X1 U699 ( .A1(G93), .A2(n647), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U701 ( .A1(G80), .A2(n650), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G55), .A2(n654), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n625) );
  OR2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n666) );
  XOR2_X1 U705 ( .A(n627), .B(n666), .Z(G145) );
  NAND2_X1 U706 ( .A1(G651), .A2(G74), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G49), .A2(n654), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U709 ( .A1(n646), .A2(n630), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n631), .A2(G87), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U712 ( .A1(G88), .A2(n647), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G75), .A2(n650), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G62), .A2(n646), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G50), .A2(n654), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U718 ( .A1(n639), .A2(n638), .ZN(G166) );
  AND2_X1 U719 ( .A1(n646), .A2(G60), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G85), .A2(n647), .ZN(n641) );
  NAND2_X1 U721 ( .A1(G72), .A2(n650), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G47), .A2(n654), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U726 ( .A1(G61), .A2(n646), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G86), .A2(n647), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U729 ( .A1(n650), .A2(G73), .ZN(n651) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n651), .Z(n652) );
  NOR2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U732 ( .A1(G48), .A2(n654), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n656), .A2(n655), .ZN(G305) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(G288), .ZN(n662) );
  XOR2_X1 U735 ( .A(n666), .B(G290), .Z(n658) );
  XNOR2_X1 U736 ( .A(G305), .B(n975), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U738 ( .A(G166), .B(n659), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n660), .B(G299), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n662), .B(n661), .ZN(n903) );
  XOR2_X1 U741 ( .A(n903), .B(n663), .Z(n664) );
  NAND2_X1 U742 ( .A1(G868), .A2(n664), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U744 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2084), .A2(G2078), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n669), .B(KEYINPUT83), .ZN(n670) );
  XNOR2_X1 U747 ( .A(KEYINPUT20), .B(n670), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U752 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U753 ( .A1(G235), .A2(G236), .ZN(n674) );
  XNOR2_X1 U754 ( .A(n674), .B(KEYINPUT85), .ZN(n675) );
  NOR2_X1 U755 ( .A1(G238), .A2(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G57), .A2(n676), .ZN(n840) );
  NAND2_X1 U757 ( .A1(n840), .A2(G567), .ZN(n682) );
  NOR2_X1 U758 ( .A1(G219), .A2(G220), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U760 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U761 ( .A1(G96), .A2(n679), .ZN(n839) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n839), .ZN(n680) );
  XNOR2_X1 U763 ( .A(KEYINPUT84), .B(n680), .ZN(n681) );
  NAND2_X1 U764 ( .A1(n682), .A2(n681), .ZN(n841) );
  NAND2_X1 U765 ( .A1(G661), .A2(G483), .ZN(n683) );
  XNOR2_X1 U766 ( .A(KEYINPUT86), .B(n683), .ZN(n684) );
  NOR2_X1 U767 ( .A1(n841), .A2(n684), .ZN(n838) );
  NAND2_X1 U768 ( .A1(n838), .A2(G36), .ZN(G176) );
  INV_X1 U769 ( .A(G166), .ZN(G303) );
  INV_X1 U770 ( .A(n975), .ZN(n685) );
  NAND2_X1 U771 ( .A1(n686), .A2(n685), .ZN(n688) );
  NOR2_X1 U772 ( .A1(G1384), .A2(G164), .ZN(n784) );
  NAND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n785) );
  INV_X1 U774 ( .A(n785), .ZN(n687) );
  NAND2_X2 U775 ( .A1(n784), .A2(n687), .ZN(n694) );
  AND2_X1 U776 ( .A1(n694), .A2(G1341), .ZN(n701) );
  NOR2_X1 U777 ( .A1(n688), .A2(n701), .ZN(n692) );
  INV_X1 U778 ( .A(G1996), .ZN(n689) );
  XNOR2_X1 U779 ( .A(n691), .B(n690), .ZN(n703) );
  NAND2_X1 U780 ( .A1(n692), .A2(n703), .ZN(n693) );
  XOR2_X1 U781 ( .A(n693), .B(KEYINPUT97), .Z(n698) );
  INV_X1 U782 ( .A(n694), .ZN(n721) );
  NOR2_X1 U783 ( .A1(n721), .A2(G1348), .ZN(n696) );
  NOR2_X1 U784 ( .A1(G2067), .A2(n694), .ZN(n695) );
  NOR2_X1 U785 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U786 ( .A1(n698), .A2(n697), .ZN(n700) );
  XNOR2_X1 U787 ( .A(n700), .B(n699), .ZN(n706) );
  NOR2_X1 U788 ( .A1(n701), .A2(n975), .ZN(n702) );
  AND2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U790 ( .A1(n982), .A2(n704), .ZN(n705) );
  NAND2_X1 U791 ( .A1(G1956), .A2(n694), .ZN(n707) );
  XNOR2_X1 U792 ( .A(KEYINPUT96), .B(n707), .ZN(n710) );
  NAND2_X1 U793 ( .A1(n721), .A2(G2072), .ZN(n708) );
  XOR2_X1 U794 ( .A(KEYINPUT27), .B(n708), .Z(n709) );
  NAND2_X1 U795 ( .A1(n710), .A2(n709), .ZN(n714) );
  NOR2_X1 U796 ( .A1(G299), .A2(n714), .ZN(n711) );
  XOR2_X1 U797 ( .A(KEYINPUT99), .B(n711), .Z(n712) );
  NOR2_X1 U798 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U799 ( .A1(G299), .A2(n714), .ZN(n715) );
  XOR2_X1 U800 ( .A(KEYINPUT28), .B(n715), .Z(n716) );
  NOR2_X1 U801 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U802 ( .A(n719), .B(n718), .ZN(n725) );
  XNOR2_X1 U803 ( .A(G2078), .B(KEYINPUT25), .ZN(n720) );
  XNOR2_X1 U804 ( .A(n720), .B(KEYINPUT95), .ZN(n1004) );
  NOR2_X1 U805 ( .A1(n1004), .A2(n694), .ZN(n723) );
  NOR2_X1 U806 ( .A1(n721), .A2(G1961), .ZN(n722) );
  NOR2_X1 U807 ( .A1(n723), .A2(n722), .ZN(n731) );
  OR2_X1 U808 ( .A1(G301), .A2(n731), .ZN(n724) );
  NAND2_X1 U809 ( .A1(n725), .A2(n724), .ZN(n748) );
  NAND2_X1 U810 ( .A1(G8), .A2(n694), .ZN(n781) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n781), .ZN(n753) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n694), .ZN(n749) );
  NOR2_X1 U813 ( .A1(n753), .A2(n749), .ZN(n726) );
  NAND2_X1 U814 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U815 ( .A(KEYINPUT101), .B(n727), .ZN(n728) );
  XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n728), .ZN(n730) );
  INV_X1 U817 ( .A(G168), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U819 ( .A1(n731), .A2(G301), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U821 ( .A(n734), .B(KEYINPUT31), .ZN(n747) );
  INV_X1 U822 ( .A(G8), .ZN(n739) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n781), .ZN(n736) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n694), .ZN(n735) );
  NOR2_X1 U825 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n737), .A2(G303), .ZN(n738) );
  OR2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n741) );
  AND2_X1 U828 ( .A1(n747), .A2(n741), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n748), .A2(n740), .ZN(n744) );
  INV_X1 U830 ( .A(n741), .ZN(n742) );
  OR2_X1 U831 ( .A1(n742), .A2(G286), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n746) );
  XOR2_X1 U833 ( .A(KEYINPUT32), .B(KEYINPUT102), .Z(n745) );
  XNOR2_X1 U834 ( .A(n746), .B(n745), .ZN(n755) );
  NAND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n751) );
  NAND2_X1 U836 ( .A1(G8), .A2(n749), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U838 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U839 ( .A1(n755), .A2(n754), .ZN(n771) );
  OR2_X1 U840 ( .A1(G303), .A2(G1971), .ZN(n757) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n764) );
  INV_X1 U842 ( .A(n764), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n972) );
  NOR2_X1 U844 ( .A1(n771), .A2(n972), .ZN(n761) );
  INV_X1 U845 ( .A(KEYINPUT103), .ZN(n758) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NAND2_X1 U847 ( .A1(n758), .A2(n974), .ZN(n759) );
  OR2_X1 U848 ( .A1(n781), .A2(n759), .ZN(n760) );
  NOR2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n764), .A2(KEYINPUT33), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n758), .A2(n763), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n764), .A2(KEYINPUT103), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n781), .A2(n767), .ZN(n769) );
  XOR2_X1 U855 ( .A(G1981), .B(G305), .Z(n983) );
  NAND2_X1 U856 ( .A1(n519), .A2(n770), .ZN(n777) );
  INV_X1 U857 ( .A(n771), .ZN(n774) );
  NOR2_X1 U858 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n775), .A2(n781), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT104), .ZN(n783) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XOR2_X1 U865 ( .A(n779), .B(KEYINPUT24), .Z(n780) );
  NOR2_X1 U866 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U867 ( .A1(n784), .A2(n785), .ZN(n829) );
  NAND2_X1 U868 ( .A1(G95), .A2(n887), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G131), .A2(n518), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U871 ( .A(KEYINPUT92), .B(n788), .Z(n792) );
  NAND2_X1 U872 ( .A1(G107), .A2(n882), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G119), .A2(n883), .ZN(n789) );
  AND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U875 ( .A1(n792), .A2(n791), .ZN(n893) );
  NAND2_X1 U876 ( .A1(G1991), .A2(n893), .ZN(n802) );
  NAND2_X1 U877 ( .A1(G117), .A2(n882), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G129), .A2(n883), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U880 ( .A1(G105), .A2(n887), .ZN(n795) );
  XNOR2_X1 U881 ( .A(KEYINPUT38), .B(n795), .ZN(n796) );
  XNOR2_X1 U882 ( .A(KEYINPUT93), .B(n796), .ZN(n797) );
  NOR2_X1 U883 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G141), .A2(n518), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n899) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n899), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n822) );
  INV_X1 U888 ( .A(n822), .ZN(n815) );
  XOR2_X1 U889 ( .A(G2067), .B(KEYINPUT37), .Z(n803) );
  XNOR2_X1 U890 ( .A(KEYINPUT89), .B(n803), .ZN(n827) );
  NAND2_X1 U891 ( .A1(n887), .A2(G104), .ZN(n805) );
  NAND2_X1 U892 ( .A1(G140), .A2(n518), .ZN(n804) );
  NAND2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n806), .B(KEYINPUT90), .ZN(n807) );
  XNOR2_X1 U895 ( .A(KEYINPUT34), .B(n807), .ZN(n812) );
  NAND2_X1 U896 ( .A1(G116), .A2(n882), .ZN(n809) );
  NAND2_X1 U897 ( .A1(G128), .A2(n883), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U899 ( .A(KEYINPUT35), .B(n810), .Z(n811) );
  NOR2_X1 U900 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U901 ( .A(KEYINPUT36), .B(n813), .ZN(n878) );
  NOR2_X1 U902 ( .A1(n827), .A2(n878), .ZN(n814) );
  XNOR2_X1 U903 ( .A(KEYINPUT91), .B(n814), .ZN(n825) );
  NAND2_X1 U904 ( .A1(n815), .A2(n825), .ZN(n966) );
  NAND2_X1 U905 ( .A1(n829), .A2(n966), .ZN(n816) );
  XOR2_X1 U906 ( .A(KEYINPUT94), .B(n816), .Z(n817) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n981) );
  NAND2_X1 U908 ( .A1(n521), .A2(n818), .ZN(n832) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n899), .ZN(n947) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n893), .ZN(n958) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U912 ( .A1(n958), .A2(n819), .ZN(n820) );
  XOR2_X1 U913 ( .A(KEYINPUT105), .B(n820), .Z(n821) );
  NOR2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U915 ( .A1(n947), .A2(n823), .ZN(n824) );
  XNOR2_X1 U916 ( .A(n824), .B(KEYINPUT39), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n827), .A2(n878), .ZN(n959) );
  NAND2_X1 U919 ( .A1(n828), .A2(n959), .ZN(n830) );
  NAND2_X1 U920 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U921 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U922 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(n834), .A2(G2106), .ZN(n835) );
  XNOR2_X1 U924 ( .A(n835), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U926 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U928 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n841), .ZN(G319) );
  XOR2_X1 U934 ( .A(KEYINPUT107), .B(G2072), .Z(n843) );
  XNOR2_X1 U935 ( .A(G2090), .B(G2078), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U937 ( .A(n844), .B(G2100), .Z(n846) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2084), .ZN(n845) );
  XNOR2_X1 U939 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U940 ( .A(G2096), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U941 ( .A(KEYINPUT42), .B(G2678), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U943 ( .A(n850), .B(n849), .Z(G227) );
  XOR2_X1 U944 ( .A(G1976), .B(G1961), .Z(n852) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1971), .ZN(n851) );
  XNOR2_X1 U946 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U947 ( .A(n853), .B(G2474), .Z(n855) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U950 ( .A(KEYINPUT41), .B(G1966), .Z(n857) );
  XNOR2_X1 U951 ( .A(G1981), .B(G1956), .ZN(n856) );
  XNOR2_X1 U952 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U953 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U954 ( .A1(n883), .A2(G124), .ZN(n860) );
  XNOR2_X1 U955 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U956 ( .A1(G136), .A2(n518), .ZN(n861) );
  NAND2_X1 U957 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U958 ( .A(KEYINPUT108), .B(n863), .ZN(n867) );
  NAND2_X1 U959 ( .A1(G112), .A2(n882), .ZN(n865) );
  NAND2_X1 U960 ( .A1(G100), .A2(n887), .ZN(n864) );
  NAND2_X1 U961 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U962 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT110), .Z(n869) );
  XNOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n869), .B(n868), .ZN(n881) );
  NAND2_X1 U966 ( .A1(G115), .A2(n882), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G127), .A2(n883), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U969 ( .A(n872), .B(KEYINPUT47), .ZN(n874) );
  NAND2_X1 U970 ( .A1(G103), .A2(n887), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n877) );
  NAND2_X1 U972 ( .A1(G139), .A2(n518), .ZN(n875) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n875), .ZN(n876) );
  NOR2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n949) );
  XNOR2_X1 U975 ( .A(n949), .B(n878), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n879), .B(n956), .ZN(n880) );
  XNOR2_X1 U977 ( .A(n881), .B(n880), .ZN(n897) );
  NAND2_X1 U978 ( .A1(G118), .A2(n882), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G130), .A2(n883), .ZN(n884) );
  NAND2_X1 U980 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U981 ( .A(KEYINPUT109), .B(n886), .Z(n892) );
  NAND2_X1 U982 ( .A1(G142), .A2(n518), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G106), .A2(n887), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U985 ( .A(n890), .B(KEYINPUT45), .Z(n891) );
  NOR2_X1 U986 ( .A1(n892), .A2(n891), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U988 ( .A(G164), .B(n895), .ZN(n896) );
  XNOR2_X1 U989 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U990 ( .A(G162), .B(n898), .ZN(n901) );
  XNOR2_X1 U991 ( .A(n899), .B(G160), .ZN(n900) );
  XNOR2_X1 U992 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U993 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U994 ( .A(G171), .B(n982), .ZN(n904) );
  XNOR2_X1 U995 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U996 ( .A(n905), .B(G286), .ZN(n906) );
  NOR2_X1 U997 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U998 ( .A(G2451), .B(G2430), .Z(n908) );
  XNOR2_X1 U999 ( .A(G2438), .B(G2443), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n908), .B(n907), .ZN(n914) );
  XOR2_X1 U1001 ( .A(G2435), .B(G2454), .Z(n910) );
  XNOR2_X1 U1002 ( .A(G1341), .B(G1348), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n912) );
  XOR2_X1 U1004 ( .A(G2446), .B(G2427), .Z(n911) );
  XNOR2_X1 U1005 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1006 ( .A(n914), .B(n913), .Z(n915) );
  NAND2_X1 U1007 ( .A1(G14), .A2(n915), .ZN(n921) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n921), .ZN(n918) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1013 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G57), .ZN(G237) );
  INV_X1 U1016 ( .A(n921), .ZN(G401) );
  XOR2_X1 U1017 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n932) );
  XNOR2_X1 U1018 ( .A(G1981), .B(G6), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(G1956), .B(G20), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n930) );
  XOR2_X1 U1021 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT59), .B(G4), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n925), .B(n924), .ZN(n926) );
  XOR2_X1 U1024 ( .A(G1348), .B(n926), .Z(n928) );
  XNOR2_X1 U1025 ( .A(G19), .B(G1341), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n932), .B(n931), .ZN(n941) );
  XOR2_X1 U1029 ( .A(G1986), .B(G24), .Z(n934) );
  XOR2_X1 U1030 ( .A(G1971), .B(G22), .Z(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G23), .B(G1976), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1034 ( .A(KEYINPUT58), .B(n937), .Z(n939) );
  XNOR2_X1 U1035 ( .A(G1966), .B(G21), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(G5), .B(G1961), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1040 ( .A(KEYINPUT61), .B(n944), .Z(n945) );
  NOR2_X1 U1041 ( .A1(G16), .A2(n945), .ZN(n1027) );
  XOR2_X1 U1042 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1044 ( .A(KEYINPUT51), .B(n948), .Z(n964) );
  XNOR2_X1 U1045 ( .A(G2072), .B(n949), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G2078), .B(KEYINPUT114), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(n950), .B(G164), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n953), .B(KEYINPUT50), .ZN(n962) );
  XOR2_X1 U1050 ( .A(G160), .B(G2084), .Z(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT113), .B(n954), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1058 ( .A(KEYINPUT52), .B(n967), .Z(n968) );
  NOR2_X1 U1059 ( .A1(KEYINPUT55), .A2(n968), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(KEYINPUT115), .B(n969), .ZN(n970) );
  NAND2_X1 U1061 ( .A1(n970), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1062 ( .A(G1956), .B(G299), .ZN(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n979) );
  NAND2_X1 U1064 ( .A1(G1971), .A2(G303), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(G1341), .B(n975), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n990) );
  XOR2_X1 U1070 ( .A(n982), .B(G1348), .Z(n988) );
  XNOR2_X1 U1071 ( .A(G168), .B(G1966), .ZN(n984) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(n985), .B(KEYINPUT57), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(KEYINPUT121), .B(n986), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1076 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1077 ( .A(G1961), .B(G171), .Z(n991) );
  XNOR2_X1 U1078 ( .A(KEYINPUT122), .B(n991), .ZN(n992) );
  NOR2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n995) );
  XOR2_X1 U1080 ( .A(G16), .B(KEYINPUT56), .Z(n994) );
  NOR2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1082 ( .A(KEYINPUT123), .B(n996), .Z(n1023) );
  XNOR2_X1 U1083 ( .A(KEYINPUT118), .B(KEYINPUT55), .ZN(n1017) );
  XOR2_X1 U1084 ( .A(G2084), .B(G34), .Z(n997) );
  XNOR2_X1 U1085 ( .A(KEYINPUT54), .B(n997), .ZN(n1014) );
  XNOR2_X1 U1086 ( .A(G2090), .B(G35), .ZN(n1012) );
  XOR2_X1 U1087 ( .A(G2072), .B(G33), .Z(n998) );
  NAND2_X1 U1088 ( .A1(G28), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G25), .B(G1991), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(G2067), .B(KEYINPUT116), .Z(n1001) );
  XNOR2_X1 U1092 ( .A(G26), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G1996), .B(G32), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1004), .B(G27), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT117), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(KEYINPUT53), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(n1015), .B(KEYINPUT119), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(n1017), .B(n1016), .ZN(n1019) );
  INV_X1 U1104 ( .A(G29), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(G11), .A2(n1020), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(KEYINPUT120), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

