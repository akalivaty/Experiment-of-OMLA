//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NOR3_X1   g005(.A1(new_n191), .A2(KEYINPUT3), .A3(G107), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(KEYINPUT75), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT75), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT76), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n195), .A2(G104), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n191), .A2(KEYINPUT75), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n198), .B1(new_n202), .B2(KEYINPUT3), .ZN(new_n203));
  AOI21_X1  g017(.A(G107), .B1(new_n194), .B2(new_n196), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n204), .A2(KEYINPUT76), .A3(new_n205), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n193), .B(new_n197), .C1(new_n203), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT4), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G101), .ZN(new_n209));
  XNOR2_X1  g023(.A(G116), .B(G119), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT2), .B(G113), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n212), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n197), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n193), .B(new_n219), .C1(new_n203), .C2(new_n206), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT4), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT76), .B1(new_n204), .B2(new_n205), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT75), .B(G104), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n198), .B(KEYINPUT3), .C1(new_n223), .C2(G107), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n192), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n217), .B1(new_n225), .B2(new_n197), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n216), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT5), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n211), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G113), .ZN(new_n231));
  INV_X1    g045(.A(G116), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G119), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n233), .B2(new_n229), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n213), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  AOI211_X1 g050(.A(new_n192), .B(new_n218), .C1(new_n222), .C2(new_n224), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n191), .A2(G107), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n217), .B1(new_n202), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT79), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT79), .ZN(new_n241));
  INV_X1    g055(.A(new_n239), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n220), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n236), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n190), .B1(new_n228), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n243), .ZN(new_n246));
  INV_X1    g060(.A(new_n236), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n215), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n226), .B2(new_n208), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n207), .A2(G101), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n248), .A2(new_n189), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n245), .A2(KEYINPUT6), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT0), .A4(G128), .ZN(new_n260));
  XNOR2_X1  g074(.A(G143), .B(G146), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT0), .B(G128), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G125), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n266), .A2(new_n257), .A3(new_n259), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n257), .A2(new_n259), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n256), .A2(G143), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n269), .A2(new_n265), .B1(KEYINPUT1), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n264), .B1(new_n272), .B2(G125), .ZN(new_n273));
  INV_X1    g087(.A(G224), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G953), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n273), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n277), .B(new_n190), .C1(new_n228), .C2(new_n244), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n255), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT7), .B1(new_n274), .B2(G953), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n273), .B(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n246), .A2(new_n247), .B1(new_n250), .B2(new_n252), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(new_n189), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n239), .B1(new_n225), .B2(new_n219), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n284), .B(new_n236), .C1(KEYINPUT79), .C2(KEYINPUT81), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n189), .B(KEYINPUT8), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT81), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n240), .B2(new_n243), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n285), .B(new_n286), .C1(new_n288), .C2(new_n236), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n279), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G210), .B1(G237), .B2(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n279), .A2(new_n292), .A3(new_n290), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n188), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(G953), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n258), .A2(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n265), .A2(G143), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G134), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n232), .A2(G122), .ZN(new_n308));
  INV_X1    g122(.A(G122), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(G116), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n199), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT14), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT87), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n232), .A2(G122), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT14), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n309), .A2(G116), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n316), .B2(KEYINPUT14), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT88), .A3(G107), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT88), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n315), .B2(new_n318), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(new_n199), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n313), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n311), .B(new_n199), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT13), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n301), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n302), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n301), .A2(new_n330), .ZN(new_n333));
  OAI21_X1  g147(.A(G134), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n334), .A3(new_n306), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n300), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n313), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT88), .B1(new_n323), .B2(G107), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n326), .A2(new_n325), .A3(new_n199), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n335), .A3(new_n299), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G902), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT89), .ZN(new_n346));
  AOI21_X1  g160(.A(G902), .B1(new_n337), .B2(new_n342), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT89), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G478), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(KEYINPUT15), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n353), .B1(new_n347), .B2(new_n348), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G140), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G125), .ZN(new_n359));
  INV_X1    g173(.A(G125), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G140), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT16), .ZN(new_n362));
  OR3_X1    g176(.A1(new_n360), .A2(KEYINPUT16), .A3(G140), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G146), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(G146), .B1(new_n362), .B2(new_n363), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G237), .ZN(new_n368));
  INV_X1    g182(.A(G953), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G214), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n258), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n368), .A2(new_n369), .A3(G143), .A4(G214), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT17), .A3(G131), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(G131), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT17), .ZN(new_n377));
  INV_X1    g191(.A(G131), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n378), .A3(new_n372), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G113), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT85), .B(G104), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XOR2_X1   g198(.A(new_n384), .B(KEYINPUT86), .Z(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT18), .A2(G131), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT83), .B1(new_n373), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n371), .A2(new_n389), .A3(new_n372), .A4(new_n386), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n392));
  XNOR2_X1  g206(.A(G125), .B(G140), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n393), .A2(new_n256), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n256), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n394), .A2(new_n395), .B1(new_n373), .B2(new_n387), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n391), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n392), .B1(new_n391), .B2(new_n396), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n381), .B(new_n385), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n375), .A2(new_n380), .ZN(new_n400));
  INV_X1    g214(.A(new_n398), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n391), .A2(new_n392), .A3(new_n396), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n384), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n399), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n344), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G475), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n408));
  XNOR2_X1  g222(.A(new_n393), .B(KEYINPUT19), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n256), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n376), .A2(new_n379), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n364), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n397), .B2(new_n398), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n384), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n399), .ZN(new_n415));
  NOR2_X1   g229(.A1(G475), .A2(G902), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n408), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n403), .A2(new_n385), .B1(new_n413), .B2(new_n384), .ZN(new_n418));
  INV_X1    g232(.A(new_n416), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n418), .A2(KEYINPUT20), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n407), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT90), .B(G952), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(G953), .ZN(new_n423));
  NAND2_X1  g237(.A1(G234), .A2(G237), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(G898), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT91), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n424), .A2(G902), .A3(G953), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n357), .A2(new_n421), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n296), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT22), .B(G137), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n369), .A2(G221), .A3(G234), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n434), .B(new_n435), .Z(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n265), .B(G119), .C1(KEYINPUT69), .C2(KEYINPUT23), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT23), .ZN(new_n439));
  INV_X1    g253(.A(G119), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(G128), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT69), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n440), .B2(G128), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n438), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G110), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT24), .B(G110), .Z(new_n446));
  XNOR2_X1  g260(.A(G119), .B(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n445), .B(new_n448), .C1(new_n365), .C2(new_n366), .ZN(new_n449));
  OAI22_X1  g263(.A1(new_n444), .A2(G110), .B1(new_n447), .B2(new_n446), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n364), .A3(new_n395), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT70), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT70), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n437), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n449), .A2(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n436), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n298), .B1(G234), .B2(new_n344), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G902), .ZN(new_n459));
  XOR2_X1   g273(.A(KEYINPUT72), .B(KEYINPUT73), .Z(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g276(.A(new_n462), .B(KEYINPUT74), .Z(new_n463));
  AOI21_X1  g277(.A(KEYINPUT25), .B1(new_n457), .B2(new_n344), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT25), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n465), .B(G902), .C1(new_n454), .C2(new_n456), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n458), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT71), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT71), .B(new_n458), .C1(new_n464), .C2(new_n466), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT32), .ZN(new_n472));
  XOR2_X1   g286(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n473));
  NAND3_X1  g287(.A1(new_n368), .A2(new_n369), .A3(G210), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT26), .B(G101), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n263), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT11), .B1(new_n305), .B2(G137), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT11), .ZN(new_n481));
  INV_X1    g295(.A(G137), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(G134), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT64), .B1(new_n482), .B2(G134), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT64), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n305), .A3(G137), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n484), .A2(new_n378), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n485), .A2(new_n487), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n378), .B1(new_n490), .B2(new_n484), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n479), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n305), .A2(G137), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n482), .A2(G134), .ZN(new_n494));
  OAI21_X1  g308(.A(G131), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n272), .A2(new_n488), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(new_n249), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT28), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G131), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n263), .B1(new_n500), .B2(new_n488), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n261), .B2(G128), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(new_n267), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n488), .A2(new_n495), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n488), .A2(KEYINPUT65), .A3(new_n495), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n509), .A2(new_n249), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n478), .B1(new_n498), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n492), .B2(new_n496), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(new_n509), .B2(new_n512), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n478), .B(new_n497), .C1(new_n514), .C2(new_n249), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT31), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n497), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n505), .A2(new_n506), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n272), .A3(new_n508), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n512), .A3(new_n492), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n505), .A2(new_n504), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT30), .B1(new_n501), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n518), .B1(new_n524), .B2(new_n215), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT31), .A3(new_n478), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n511), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(G472), .A2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n472), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n511), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT31), .B1(new_n525), .B2(new_n478), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n249), .B1(new_n521), .B2(new_n523), .ZN(new_n533));
  NOR4_X1   g347(.A1(new_n533), .A2(new_n516), .A3(new_n477), .A4(new_n518), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT32), .A3(new_n528), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(new_n536), .A3(KEYINPUT68), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT68), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n535), .A2(new_n538), .A3(KEYINPUT32), .A4(new_n528), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n498), .A2(new_n510), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n477), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT29), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n497), .B1(new_n514), .B2(new_n249), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n477), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n498), .A2(KEYINPUT67), .A3(new_n478), .A4(new_n510), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n543), .A2(new_n544), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n215), .B1(new_n501), .B2(new_n522), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n498), .A2(new_n549), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n550), .A2(new_n544), .A3(new_n477), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n471), .B1(new_n540), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G221), .ZN(new_n556));
  INV_X1    g370(.A(new_n297), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n344), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT10), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n504), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n263), .B1(new_n226), .B2(new_n208), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n246), .A2(new_n561), .B1(new_n562), .B2(new_n252), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n271), .A2(KEYINPUT77), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT77), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n503), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n566), .A3(new_n268), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n220), .A2(new_n242), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT78), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT78), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n284), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n560), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n489), .A2(new_n491), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n563), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n240), .A2(new_n504), .A3(new_n243), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n574), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT12), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT12), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n580), .B(new_n574), .C1(new_n572), .C2(new_n576), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n575), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G110), .B(G140), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n369), .A2(G227), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  AOI211_X1 g400(.A(KEYINPUT79), .B(new_n239), .C1(new_n225), .C2(new_n219), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n241), .B1(new_n220), .B2(new_n242), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n561), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n209), .B(new_n479), .C1(new_n221), .C2(new_n226), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT10), .B1(new_n569), .B2(new_n571), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n578), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n585), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n575), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n586), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G469), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT80), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT80), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n591), .A2(new_n592), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n585), .B1(new_n600), .B2(new_n574), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n582), .A2(new_n585), .B1(new_n601), .B2(new_n593), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n599), .B(G469), .C1(new_n602), .C2(G902), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n574), .B1(new_n563), .B2(new_n573), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n591), .A2(new_n592), .A3(new_n578), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n585), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n575), .B(new_n594), .C1(new_n579), .C2(new_n581), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n597), .A3(new_n344), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n598), .A2(new_n603), .A3(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n433), .A2(new_n555), .A3(new_n559), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT92), .B(G101), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G3));
  AND2_X1   g427(.A1(new_n610), .A2(new_n559), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n343), .A2(KEYINPUT33), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n337), .A2(new_n342), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(G478), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n347), .A2(new_n351), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n351), .A2(new_n344), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n421), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(KEYINPUT93), .Z(new_n625));
  INV_X1    g439(.A(new_n430), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n279), .A2(new_n292), .A3(new_n290), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n292), .B1(new_n279), .B2(new_n290), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n187), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G472), .B1(new_n527), .B2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n535), .A2(new_n528), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n471), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n614), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT94), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT34), .B(G104), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n187), .B1(new_n627), .B2(new_n628), .ZN(new_n641));
  INV_X1    g455(.A(new_n408), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n418), .B2(new_n419), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n415), .A2(new_n408), .A3(new_n416), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT95), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n415), .A2(KEYINPUT95), .A3(new_n408), .A4(new_n416), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n649), .A2(new_n357), .A3(new_n626), .A4(new_n407), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n640), .B1(new_n641), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n352), .B1(new_n346), .B2(new_n349), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n407), .B1(new_n652), .B2(new_n355), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n653), .A2(new_n648), .A3(new_n430), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n296), .A2(KEYINPUT96), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n614), .A2(new_n635), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n452), .A2(new_n453), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n437), .A2(KEYINPUT36), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n461), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n469), .A2(new_n470), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n660), .B1(new_n633), .B2(new_n665), .ZN(new_n666));
  AND4_X1   g480(.A1(new_n660), .A2(new_n665), .A3(new_n632), .A4(new_n631), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(new_n559), .A3(new_n610), .A4(new_n433), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT98), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  INV_X1    g486(.A(new_n665), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n540), .B2(new_n554), .ZN(new_n674));
  INV_X1    g488(.A(G900), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n426), .B1(new_n675), .B2(new_n429), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n653), .A2(new_n648), .A3(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n296), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n674), .A2(new_n678), .A3(new_n610), .A4(new_n559), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XOR2_X1   g494(.A(new_n676), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n614), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n294), .A2(new_n295), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n525), .A2(new_n477), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n549), .A2(new_n477), .A3(new_n497), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n344), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n540), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n357), .A2(new_n421), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n665), .A3(new_n188), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n687), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n683), .A2(new_n684), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT100), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n683), .A2(new_n698), .A3(new_n684), .A4(new_n695), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT101), .B(G143), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G45));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n674), .A2(new_n559), .A3(new_n610), .ZN(new_n704));
  INV_X1    g518(.A(G475), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n405), .B2(new_n344), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT20), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n415), .A2(new_n707), .A3(new_n416), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n706), .B1(new_n643), .B2(new_n708), .ZN(new_n709));
  OR3_X1    g523(.A1(new_n709), .A2(new_n622), .A3(new_n676), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT102), .B1(new_n641), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n624), .A2(new_n676), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n296), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n703), .B1(new_n704), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n711), .A2(new_n714), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n614), .A2(KEYINPUT103), .A3(new_n674), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  AOI21_X1  g535(.A(G902), .B1(new_n606), .B2(new_n607), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(new_n597), .ZN(new_n723));
  OAI21_X1  g537(.A(G469), .B1(new_n722), .B2(KEYINPUT104), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n725), .B(G902), .C1(new_n606), .C2(new_n607), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n723), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n594), .B1(new_n593), .B2(new_n575), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n579), .A2(new_n581), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n728), .B1(new_n729), .B2(new_n601), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n725), .B1(new_n730), .B2(G902), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n721), .A3(G469), .A4(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n558), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n630), .A2(new_n734), .A3(new_n555), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT41), .B(G113), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT106), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n735), .B(new_n737), .ZN(G15));
  NAND3_X1  g552(.A1(new_n734), .A2(new_n656), .A3(new_n555), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  INV_X1    g554(.A(G472), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n548), .B2(new_n552), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n742), .B1(new_n537), .B2(new_n539), .ZN(new_n743));
  INV_X1    g557(.A(new_n431), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n673), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n734), .A2(new_n296), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  INV_X1    g561(.A(new_n471), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n478), .B1(new_n550), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n498), .A2(KEYINPUT107), .A3(new_n549), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n532), .A2(new_n534), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n749), .B(new_n528), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n751), .A2(new_n752), .B1(new_n517), .B2(new_n526), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT108), .B1(new_n756), .B2(new_n529), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n748), .A2(new_n631), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n758), .A2(new_n629), .A3(new_n693), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n734), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  NAND2_X1  g575(.A1(new_n727), .A2(new_n733), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n757), .A3(new_n665), .A4(new_n631), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n710), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n559), .A3(new_n296), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  NOR3_X1   g580(.A1(new_n627), .A2(new_n628), .A3(new_n188), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n597), .A2(new_n344), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n722), .B2(new_n597), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n601), .B2(new_n593), .ZN(new_n771));
  AND4_X1   g585(.A1(new_n770), .A2(new_n593), .A3(new_n575), .A4(new_n594), .ZN(new_n772));
  OAI211_X1 g586(.A(G469), .B(new_n586), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n558), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n555), .A2(new_n713), .A3(new_n767), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n778));
  INV_X1    g592(.A(new_n768), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n609), .A3(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n624), .A2(new_n776), .A3(new_n676), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n767), .A3(new_n559), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n536), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n535), .A2(KEYINPUT110), .A3(KEYINPUT32), .A4(new_n528), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n554), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n530), .B(KEYINPUT111), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n471), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n778), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n530), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n554), .A2(new_n785), .A3(new_n786), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n748), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n782), .A3(KEYINPUT112), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n777), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n777), .B(KEYINPUT113), .C1(new_n790), .C2(new_n795), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G131), .ZN(G33));
  NAND4_X1  g615(.A1(new_n555), .A2(new_n677), .A3(new_n767), .A4(new_n774), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  NAND2_X1  g617(.A1(new_n586), .A2(new_n595), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n597), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(KEYINPUT45), .B(new_n586), .C1(new_n771), .C2(new_n772), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n768), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(KEYINPUT46), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n609), .B1(new_n808), .B2(KEYINPUT46), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n559), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n681), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n294), .A2(new_n187), .A3(new_n295), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n421), .A2(new_n622), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT43), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n634), .A3(new_n665), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT44), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n813), .B(new_n819), .C1(new_n818), .C2(new_n817), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G137), .ZN(G39));
  NAND4_X1  g635(.A1(new_n743), .A2(new_n471), .A3(new_n713), .A4(new_n767), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n809), .A2(new_n810), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(KEYINPUT47), .A3(new_n559), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n811), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g641(.A(KEYINPUT114), .B(G140), .Z(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(G42));
  NAND2_X1  g643(.A1(new_n765), .A2(new_n679), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n693), .A2(new_n665), .A3(new_n676), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n692), .A2(new_n774), .A3(new_n296), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n719), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n716), .B2(new_n718), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n765), .B2(new_n679), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n735), .A2(new_n739), .A3(new_n746), .A4(new_n760), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n357), .A2(new_n846), .A3(new_n709), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n355), .B1(new_n350), .B2(new_n353), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT116), .B1(new_n421), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n847), .A2(new_n849), .A3(new_n624), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n629), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n610), .A3(new_n559), .A4(new_n635), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n669), .A2(new_n611), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n706), .A2(new_n676), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n649), .A2(new_n848), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n814), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n674), .A2(new_n610), .A3(new_n856), .A4(new_n559), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n764), .A2(new_n767), .A3(new_n774), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n802), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n798), .A2(new_n799), .A3(new_n845), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n843), .A2(new_n844), .A3(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n834), .A2(new_n835), .B1(new_n831), .B2(new_n838), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n798), .A2(new_n845), .A3(new_n860), .A4(new_n799), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT53), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n865), .A3(KEYINPUT54), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n844), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n860), .A2(new_n845), .A3(KEYINPUT53), .A4(new_n796), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n843), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n734), .A2(new_n767), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n816), .A2(new_n426), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n816), .A2(new_n877), .A3(new_n426), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n763), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n874), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n692), .A2(new_n471), .A3(new_n425), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n421), .A2(new_n623), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n874), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n758), .B1(new_n876), .B2(new_n878), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n687), .A2(new_n187), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n734), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT50), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n886), .A2(KEYINPUT50), .A3(new_n734), .A4(new_n887), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n885), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n762), .A2(new_n558), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n824), .A2(new_n826), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n886), .A2(new_n767), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n892), .A2(new_n896), .A3(KEYINPUT51), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n892), .A2(new_n896), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT51), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n892), .A2(new_n896), .A3(KEYINPUT119), .A4(KEYINPUT51), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n886), .A2(new_n296), .A3(new_n734), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n874), .A2(new_n882), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n904), .B(new_n423), .C1(new_n905), .C2(new_n625), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n874), .A2(new_n879), .A3(new_n789), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n907), .A2(KEYINPUT48), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(KEYINPUT48), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n899), .A2(new_n902), .A3(new_n903), .A4(new_n910), .ZN(new_n911));
  OAI22_X1  g725(.A1(new_n873), .A2(new_n911), .B1(G952), .B2(G953), .ZN(new_n912));
  INV_X1    g726(.A(new_n762), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n913), .A2(KEYINPUT49), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(KEYINPUT49), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n815), .A2(new_n559), .A3(new_n187), .ZN(new_n916));
  NOR4_X1   g730(.A1(new_n687), .A2(new_n471), .A3(new_n692), .A4(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT115), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n912), .A2(KEYINPUT120), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(G75));
  INV_X1    g738(.A(new_n837), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n719), .A2(new_n831), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n765), .A2(new_n679), .A3(new_n833), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n716), .B2(new_n718), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n928), .B2(KEYINPUT52), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT53), .B1(new_n861), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n868), .B1(new_n836), .B2(new_n842), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n344), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT56), .B1(new_n933), .B2(G210), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n255), .A2(new_n278), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n276), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT55), .Z(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n369), .A2(G952), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n934), .B2(new_n938), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n939), .A2(new_n942), .ZN(G51));
  NAND2_X1  g757(.A1(new_n867), .A2(new_n870), .ZN(new_n944));
  AND4_X1   g758(.A1(G902), .A2(new_n944), .A3(new_n807), .A4(new_n806), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT54), .B1(new_n930), .B2(new_n931), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n872), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n768), .B(KEYINPUT57), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n730), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n948), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n946), .B2(new_n872), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT121), .B1(new_n953), .B2(new_n730), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n940), .B1(new_n951), .B2(new_n954), .ZN(G54));
  NAND2_X1  g769(.A1(new_n944), .A2(G902), .ZN(new_n956));
  NAND2_X1  g770(.A1(KEYINPUT58), .A2(G475), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n418), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n957), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n944), .A2(G902), .A3(new_n415), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n941), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT122), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n958), .A2(KEYINPUT122), .A3(new_n941), .A4(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G60));
  XNOR2_X1  g779(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n621), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n873), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n615), .A2(new_n617), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT123), .Z(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n971), .A2(new_n967), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT54), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n871), .B1(new_n867), .B2(new_n870), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n972), .A2(new_n973), .A3(new_n941), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n941), .ZN(new_n979));
  INV_X1    g793(.A(new_n971), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n873), .B2(new_n968), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT125), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n978), .A2(new_n982), .ZN(G63));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT126), .Z(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT60), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n932), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n663), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n941), .B1(new_n988), .B2(new_n457), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n984), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n988), .A2(new_n457), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n993), .A2(KEYINPUT61), .A3(new_n941), .A4(new_n989), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(G66));
  OAI21_X1  g809(.A(G953), .B1(new_n428), .B2(new_n274), .ZN(new_n996));
  INV_X1    g810(.A(new_n853), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n845), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n996), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n935), .B1(G898), .B2(new_n369), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(G69));
  AOI21_X1  g816(.A(new_n369), .B1(G227), .B2(G900), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n514), .B(new_n409), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n839), .A2(new_n841), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n800), .A2(new_n719), .A3(new_n1005), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n794), .A2(new_n641), .A3(new_n693), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n813), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n820), .A2(new_n802), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1009), .A2(new_n827), .ZN(new_n1010));
  AOI21_X1  g824(.A(G953), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n369), .A2(G900), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT127), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n827), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1014), .A2(new_n802), .A3(new_n820), .A4(new_n1008), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n800), .A2(new_n719), .A3(new_n1005), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n369), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1012), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1004), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1004), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1005), .A2(new_n719), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT62), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1023), .A2(new_n1024), .A3(new_n699), .A4(new_n697), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1005), .A2(new_n719), .ZN(new_n1026));
  OAI21_X1  g840(.A(KEYINPUT62), .B1(new_n700), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n850), .A2(new_n814), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n555), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n820), .B1(new_n682), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1030), .A2(new_n827), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1025), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1022), .B1(new_n1032), .B2(new_n369), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1003), .B1(new_n1021), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1020), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1018), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1022), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1003), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1033), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1034), .A2(new_n1040), .ZN(G72));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  NAND2_X1  g857(.A1(new_n546), .A2(new_n515), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n862), .A2(new_n865), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1045), .A2(new_n941), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1006), .A2(new_n1010), .A3(new_n999), .ZN(new_n1047));
  AOI211_X1 g861(.A(new_n478), .B(new_n545), .C1(new_n1047), .C2(new_n1043), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1043), .B1(new_n1032), .B2(new_n998), .ZN(new_n1049));
  AOI211_X1 g863(.A(new_n1046), .B(new_n1048), .C1(new_n688), .C2(new_n1049), .ZN(G57));
endmodule


