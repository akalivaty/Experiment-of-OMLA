//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g0008(.A(new_n208), .B1(G68), .B2(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n203), .A2(G13), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT0), .Z(new_n233));
  NOR3_X1   g0033(.A1(new_n223), .A2(new_n230), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n211), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G222), .ZN(new_n257));
  INV_X1    g0057(.A(G223), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n255), .B(new_n257), .C1(new_n258), .C2(new_n256), .ZN(new_n259));
  AND2_X1   g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n229), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n259), .B(new_n261), .C1(G77), .C2(new_n255), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT65), .B1(new_n260), .B2(new_n229), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT65), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n263), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(new_n264), .B2(new_n268), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n262), .B(new_n273), .C1(new_n275), .C2(new_n215), .ZN(new_n276));
  XOR2_X1   g0076(.A(KEYINPUT67), .B(G179), .Z(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n229), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT66), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT66), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(G20), .B1(new_n225), .B2(G50), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n250), .A2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n287), .B1(new_n288), .B2(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G1), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n286), .A2(new_n294), .B1(new_n214), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n283), .A2(new_n285), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n296), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n214), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n276), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n279), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n276), .A2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n307), .B1(new_n308), .B2(new_n276), .C1(new_n309), .C2(new_n302), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n302), .A2(new_n309), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n310), .A2(KEYINPUT10), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT10), .B1(new_n310), .B2(new_n311), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n306), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n298), .A2(new_n293), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n301), .B2(new_n293), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT7), .A2(G20), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT72), .B1(new_n252), .B2(G33), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT72), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(new_n250), .A3(KEYINPUT3), .ZN(new_n321));
  AOI211_X1 g0121(.A(KEYINPUT73), .B(new_n318), .C1(new_n319), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT73), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n321), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n253), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n317), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n318), .B1(new_n319), .B2(new_n321), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT7), .B1(new_n327), .B2(G20), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(G68), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(G58), .B(G68), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(G20), .B1(G159), .B2(new_n289), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT7), .B1(new_n254), .B2(new_n228), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  AOI211_X1 g0134(.A(new_n334), .B(G20), .C1(new_n251), .C2(new_n253), .ZN(new_n335));
  OAI21_X1  g0135(.A(G68), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n331), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n282), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n316), .B1(new_n332), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT76), .ZN(new_n341));
  INV_X1    g0141(.A(new_n261), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n258), .A2(G1698), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n320), .B1(KEYINPUT3), .B2(new_n250), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n252), .A2(KEYINPUT72), .A3(G33), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n253), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n250), .A2(new_n204), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n256), .A2(KEYINPUT75), .A3(G223), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G226), .A2(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(new_n327), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n342), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n264), .A2(new_n268), .ZN(new_n355));
  INV_X1    g0155(.A(new_n272), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(G232), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n273), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n341), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n324), .A2(new_n253), .A3(new_n352), .ZN(new_n360));
  INV_X1    g0160(.A(new_n349), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT75), .B1(new_n327), .B2(new_n343), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n261), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(G232), .A2(new_n274), .B1(new_n269), .B2(new_n272), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(KEYINPUT76), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(G200), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n354), .A2(new_n358), .A3(G190), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n340), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT17), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n340), .B(KEYINPUT17), .C1(new_n367), .C2(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n354), .A2(new_n358), .A3(new_n278), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n359), .A2(new_n366), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n303), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT74), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n332), .A2(new_n339), .ZN(new_n378));
  INV_X1    g0178(.A(new_n316), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI211_X1 g0180(.A(KEYINPUT74), .B(new_n316), .C1(new_n332), .C2(new_n339), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(KEYINPUT18), .B(new_n376), .C1(new_n380), .C2(new_n381), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n373), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n228), .A2(G1), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n281), .A2(new_n387), .A3(new_n216), .ZN(new_n388));
  INV_X1    g0188(.A(new_n293), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n292), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(new_n281), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n298), .A2(new_n216), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G238), .A2(G1698), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n255), .B(new_n397), .C1(new_n220), .C2(G1698), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n261), .C1(G107), .C2(new_n255), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(new_n273), .C1(new_n217), .C2(new_n275), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G200), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n396), .B(new_n401), .C1(new_n308), .C2(new_n400), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n291), .A2(G77), .B1(G20), .B2(new_n224), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n214), .B2(new_n290), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(new_n285), .A3(new_n283), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT11), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT11), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n286), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT71), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n387), .A2(G13), .A3(new_n224), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT12), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n296), .A2(new_n280), .A3(G68), .A4(new_n229), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT68), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n414), .A3(KEYINPUT69), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT69), .B1(new_n412), .B2(new_n414), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n409), .B(new_n410), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n412), .A2(new_n414), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT69), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n415), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n410), .B1(new_n423), .B2(new_n409), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n274), .A2(G238), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n215), .A2(new_n256), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n220), .A2(G1698), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n427), .B1(new_n254), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n261), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n273), .A2(new_n426), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT13), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n273), .A2(new_n426), .A3(new_n432), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT70), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT14), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n437), .A2(G169), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n437), .B2(G169), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G179), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n425), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n437), .A2(new_n308), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n423), .A2(new_n409), .ZN(new_n448));
  INV_X1    g0248(.A(G200), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n434), .B2(new_n436), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n400), .A2(new_n278), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n400), .A2(new_n303), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n395), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n446), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  AND4_X1   g0256(.A1(new_n314), .A2(new_n386), .A3(new_n402), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n204), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n327), .A2(new_n228), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT79), .B(G116), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n291), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n228), .A2(G107), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n464), .B(KEYINPUT23), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n228), .A2(G87), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n458), .B1(new_n254), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n460), .A2(new_n463), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n468), .A2(KEYINPUT24), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(KEYINPUT24), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n282), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n298), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n295), .A2(G33), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n300), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n210), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n298), .A2(new_n210), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT25), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT83), .B1(new_n471), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n470), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n468), .A2(KEYINPUT24), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n281), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT83), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n475), .A2(new_n477), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  NOR2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n295), .B(G45), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n355), .A2(G264), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT84), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n355), .A2(new_n491), .A3(G264), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n205), .A2(new_n256), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n207), .A2(G1698), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n327), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G294), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n261), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n486), .A2(new_n487), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n269), .A2(G45), .A3(new_n272), .A4(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n493), .A2(G179), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n489), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n342), .B1(new_n496), .B2(new_n497), .ZN(new_n504));
  OAI21_X1  g0304(.A(G169), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT85), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n502), .A2(KEYINPUT85), .A3(new_n505), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n479), .A2(new_n485), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n217), .A2(G1698), .ZN(new_n511));
  OR2_X1    g0311(.A1(G238), .A2(G1698), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n327), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n462), .A2(G33), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n261), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT80), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n205), .B1(new_n271), .B2(G1), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n295), .A2(new_n263), .A3(G45), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n355), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n342), .B1(new_n513), .B2(new_n514), .ZN(new_n522));
  INV_X1    g0322(.A(new_n520), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT80), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n277), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n327), .A2(new_n228), .A3(G68), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n228), .B1(new_n427), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n204), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n528), .B1(new_n427), .B2(G20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n527), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n281), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n298), .A2(new_n391), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n474), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n391), .B(KEYINPUT81), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n521), .A2(new_n303), .A3(new_n524), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n526), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n525), .A2(G190), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n521), .A2(G200), .A3(new_n524), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n535), .B(new_n536), .C1(new_n204), .C2(new_n474), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n510), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n324), .A2(G244), .A3(new_n253), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(new_n553), .B1(G33), .B2(G283), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT4), .B1(new_n254), .B2(new_n205), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n254), .A2(new_n217), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n553), .A2(G1698), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n555), .A2(G1698), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n261), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n355), .A2(G257), .A3(new_n488), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n501), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT77), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n342), .B1(new_n554), .B2(new_n558), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT77), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n565), .A2(new_n566), .A3(new_n562), .ZN(new_n567));
  OAI21_X1  g0367(.A(G190), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n210), .A2(KEYINPUT6), .A3(G97), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n206), .A2(new_n210), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(new_n530), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n571), .B2(KEYINPUT6), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(G20), .B1(G77), .B2(new_n289), .ZN(new_n573));
  OAI21_X1  g0373(.A(G107), .B1(new_n333), .B2(new_n335), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n282), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n474), .A2(new_n206), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n472), .A2(G97), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n560), .A2(new_n563), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G200), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n568), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n560), .A2(KEYINPUT77), .A3(new_n563), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n566), .B1(new_n565), .B2(new_n562), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n303), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT78), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n579), .B2(new_n278), .ZN(new_n586));
  INV_X1    g0386(.A(new_n578), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n560), .A2(KEYINPUT78), .A3(new_n277), .A4(new_n563), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n584), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n504), .B1(new_n490), .B2(new_n492), .ZN(new_n590));
  AOI21_X1  g0390(.A(G200), .B1(new_n590), .B2(new_n501), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n503), .A2(G190), .A3(new_n504), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n482), .B(new_n484), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n581), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n298), .A2(new_n461), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n472), .A2(G116), .A3(new_n282), .A4(new_n473), .ZN(new_n596));
  AOI21_X1  g0396(.A(G20), .B1(G33), .B2(G283), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(G33), .B2(new_n206), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n281), .B(new_n598), .C1(new_n462), .C2(new_n228), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT20), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n595), .B(new_n596), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n207), .A2(new_n256), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n211), .A2(G1698), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n324), .A2(new_n253), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n254), .A2(G303), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n261), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n355), .A2(G270), .A3(new_n488), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n501), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n603), .A2(G169), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n611), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(new_n603), .A3(G179), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n603), .A2(KEYINPUT21), .A3(new_n611), .A4(G169), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n603), .B1(new_n615), .B2(G190), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(G200), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT82), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT82), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n619), .A2(new_n623), .A3(new_n620), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n618), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n457), .A2(new_n551), .A3(new_n594), .A4(new_n625), .ZN(G372));
  NAND2_X1  g0426(.A1(new_n378), .A2(new_n379), .ZN(new_n627));
  XNOR2_X1  g0427(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n627), .A2(new_n376), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n627), .B2(new_n376), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n451), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n446), .B1(new_n632), .B2(new_n455), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n633), .B2(new_n373), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n312), .A2(new_n313), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n457), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n547), .B1(new_n525), .B2(G190), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n516), .A2(new_n520), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G200), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n482), .A2(new_n484), .B1(new_n505), .B2(new_n502), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n581), .B(new_n593), .C1(new_n644), .C2(new_n618), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n645), .B2(new_n589), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT26), .B1(new_n550), .B2(new_n589), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n525), .A2(new_n277), .B1(new_n538), .B2(new_n541), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n639), .A2(new_n303), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n305), .B(new_n636), .C1(new_n637), .C2(new_n652), .ZN(G369));
  NAND2_X1  g0453(.A1(new_n508), .A2(new_n509), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n471), .A2(new_n478), .A3(KEYINPUT83), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n297), .A2(G20), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OR3_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .A3(G1), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT27), .B1(new_n659), .B2(G1), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT87), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT87), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n655), .B2(new_n656), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n657), .A2(new_n668), .A3(new_n593), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT88), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT88), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n510), .A2(new_n667), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n603), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n625), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n618), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n675), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n667), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n644), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n677), .A2(new_n667), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n670), .A2(new_n671), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT89), .ZN(G399));
  NOR2_X1   g0487(.A1(new_n531), .A2(G116), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT90), .ZN(new_n689));
  INV_X1    g0489(.A(new_n231), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n689), .A2(new_n295), .A3(new_n691), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT91), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT91), .ZN(new_n694));
  INV_X1    g0494(.A(new_n691), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n693), .B(new_n694), .C1(new_n226), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n609), .A2(G179), .A3(new_n501), .A4(new_n610), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n524), .B2(new_n521), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n699), .B(new_n590), .C1(new_n564), .C2(new_n567), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT30), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n700), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n615), .A2(new_n278), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n590), .A2(new_n501), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n579), .A4(new_n639), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n667), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n594), .A2(new_n551), .A3(new_n625), .A4(new_n682), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT31), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n713), .A3(new_n667), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n682), .B1(new_n646), .B2(new_n651), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n718), .B1(new_n720), .B2(KEYINPUT93), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n648), .A2(new_n649), .B1(new_n638), .B2(new_n640), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n589), .A3(new_n581), .A4(new_n593), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n510), .A2(new_n618), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n657), .A2(new_n677), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n594), .A2(new_n727), .A3(KEYINPUT94), .A4(new_n723), .ZN(new_n728));
  INV_X1    g0528(.A(new_n650), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n642), .B1(new_n550), .B2(new_n589), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n584), .A2(new_n587), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n586), .A2(new_n588), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT26), .A4(new_n641), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n726), .A2(new_n728), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n682), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT29), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n717), .A2(new_n721), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n697), .B1(new_n740), .B2(G1), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT95), .ZN(G364));
  NOR2_X1   g0542(.A1(new_n228), .A2(G179), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n744));
  INV_X1    g0544(.A(G303), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n277), .A2(new_n228), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G190), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G311), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n747), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n308), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT97), .B(G326), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n254), .B(new_n751), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n308), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n756), .B1(G322), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n747), .A2(new_n308), .A3(G200), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT98), .B(G317), .Z(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT33), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n760), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n743), .A2(new_n748), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n746), .B(new_n764), .C1(G329), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G283), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n743), .A2(new_n308), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(G294), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n757), .A2(new_n443), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n767), .B1(new_n768), .B2(new_n769), .C1(new_n770), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n206), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n765), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(KEYINPUT32), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n749), .A2(KEYINPUT96), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n749), .A2(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n775), .B(new_n779), .C1(new_n783), .C2(G77), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n214), .B2(new_n754), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(KEYINPUT32), .B2(new_n778), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n769), .A2(new_n210), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n758), .A2(new_n219), .B1(new_n204), .B2(new_n744), .ZN(new_n789));
  INV_X1    g0589(.A(new_n761), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G68), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n786), .A2(new_n255), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n774), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n229), .B1(G20), .B2(new_n303), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n255), .A2(G355), .A3(new_n231), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n322), .A2(new_n325), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n690), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G45), .B2(new_n227), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n245), .A2(new_n271), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n796), .B1(G116), .B2(new_n231), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G13), .A2(G33), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n794), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n804), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n678), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n295), .B1(new_n658), .B2(G45), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n691), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n795), .A2(new_n806), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n680), .A2(new_n811), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(G330), .B2(new_n678), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(G396));
  OR3_X1    g0615(.A1(new_n454), .A2(KEYINPUT102), .A3(new_n682), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT102), .B1(new_n454), .B2(new_n682), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n454), .B(KEYINPUT101), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n667), .A2(new_n395), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n402), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n719), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n717), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT103), .ZN(new_n826));
  INV_X1    g0626(.A(new_n811), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(KEYINPUT103), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT104), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n717), .A2(new_n824), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n826), .A2(KEYINPUT104), .A3(new_n827), .A4(new_n828), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n769), .A2(new_n224), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n783), .A2(G159), .B1(G143), .B2(new_n759), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n837), .B2(new_n754), .C1(new_n288), .C2(new_n761), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT34), .ZN(new_n839));
  INV_X1    g0639(.A(new_n797), .ZN(new_n840));
  INV_X1    g0640(.A(new_n744), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(G50), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n839), .B(new_n842), .C1(new_n843), .C2(new_n765), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n835), .B(new_n844), .C1(G58), .C2(new_n772), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n753), .A2(G303), .B1(new_n759), .B2(G294), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n204), .B2(new_n769), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n761), .A2(KEYINPUT100), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n761), .A2(KEYINPUT100), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n847), .B1(new_n850), .B2(G283), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n255), .B(new_n775), .C1(G311), .C2(new_n766), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(new_n461), .C2(new_n782), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G107), .B2(new_n841), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n794), .B1(new_n845), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n794), .A2(new_n802), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n811), .B1(G77), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT99), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n855), .B(new_n859), .C1(new_n803), .C2(new_n822), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n834), .A2(new_n860), .ZN(G384));
  INV_X1    g0661(.A(KEYINPUT108), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n368), .B1(new_n375), .B2(new_n449), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT107), .B1(new_n627), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n627), .A2(new_n376), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT107), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n340), .B(new_n866), .C1(new_n367), .C2(new_n368), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT106), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n665), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n627), .A2(KEYINPUT74), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n340), .A2(new_n377), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT37), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n665), .B(KEYINPUT106), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n380), .B2(new_n381), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n382), .A2(new_n876), .A3(new_n877), .A4(new_n369), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n372), .B(new_n371), .C1(new_n629), .C2(new_n630), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n874), .A2(new_n878), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n862), .B1(new_n880), .B2(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n382), .A2(new_n369), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n876), .A2(new_n865), .A3(new_n864), .A4(new_n867), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n883), .A2(new_n884), .B1(new_n885), .B2(KEYINPUT37), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n879), .A2(new_n873), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT108), .B(new_n882), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n329), .A2(new_n331), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n338), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n890), .A2(new_n286), .A3(new_n332), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n376), .B1(new_n891), .B2(new_n316), .ZN(new_n892));
  INV_X1    g0692(.A(new_n665), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n891), .B2(new_n316), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n892), .A2(new_n894), .A3(new_n369), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n878), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n897), .B(KEYINPUT38), .C1(new_n386), .C2(new_n894), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n881), .A2(new_n888), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n446), .B2(new_n451), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n632), .B(KEYINPUT105), .C1(new_n902), .C2(new_n425), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n425), .A2(new_n682), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n900), .B1(new_n425), .B2(new_n682), .C1(new_n446), .C2(new_n451), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n822), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n715), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT40), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT109), .B1(new_n715), .B2(new_n907), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n905), .A2(new_n822), .A3(new_n906), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT109), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n912), .A2(new_n712), .A3(new_n714), .A4(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n386), .A2(new_n894), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n883), .A2(new_n884), .B1(new_n895), .B2(KEYINPUT37), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n882), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n898), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n915), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n910), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n716), .A2(new_n457), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(G330), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n631), .A2(new_n875), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n819), .A2(new_n682), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n719), .B2(new_n823), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n905), .A2(new_n906), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n925), .B1(new_n930), .B2(new_n919), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n899), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n446), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(new_n667), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n918), .A2(new_n898), .A3(KEYINPUT39), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n636), .A2(new_n305), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n738), .A2(new_n721), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(new_n457), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n938), .B(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n924), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n295), .B2(new_n658), .ZN(new_n944));
  INV_X1    g0744(.A(G116), .ZN(new_n945));
  OAI211_X1 g0745(.A(G20), .B(new_n265), .C1(new_n572), .C2(KEYINPUT35), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n945), .B(new_n946), .C1(KEYINPUT35), .C2(new_n572), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT36), .Z(new_n948));
  OAI21_X1  g0748(.A(G77), .B1(new_n219), .B2(new_n224), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n226), .A2(new_n949), .B1(G50), .B2(new_n224), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(G1), .A3(new_n297), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n944), .A2(new_n948), .A3(new_n951), .ZN(G367));
  OAI211_X1 g0752(.A(new_n581), .B(new_n589), .C1(new_n578), .C2(new_n682), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n731), .A2(new_n732), .A3(new_n667), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT42), .B1(new_n685), .B2(new_n956), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n685), .A2(KEYINPUT42), .A3(new_n956), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n510), .A2(new_n581), .B1(new_n731), .B2(new_n732), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n957), .B(new_n958), .C1(new_n667), .C2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n723), .B1(new_n548), .B2(new_n682), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n729), .A2(new_n547), .A3(new_n667), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n960), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n960), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n681), .B1(new_n953), .B2(new_n954), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n691), .B(KEYINPUT41), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n685), .A2(new_n683), .A3(new_n955), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n973), .A2(KEYINPUT110), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(KEYINPUT110), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n955), .B1(new_n685), .B2(new_n683), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT44), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n974), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n681), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n685), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT111), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT111), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n685), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n988), .C1(new_n674), .C2(new_n684), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(new_n680), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n680), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n739), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n978), .A2(new_n980), .A3(new_n681), .A4(new_n981), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n984), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n972), .B1(new_n994), .B2(new_n740), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n970), .B1(new_n995), .B2(new_n810), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n850), .A2(G294), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n841), .A2(KEYINPUT46), .A3(G116), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n744), .B2(new_n461), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n769), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(G97), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n758), .A2(new_n745), .B1(new_n210), .B2(new_n773), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n753), .A2(G311), .ZN(new_n1005));
  NOR4_X1   g0805(.A1(new_n1003), .A2(new_n797), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(G317), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(new_n768), .B2(new_n782), .C1(new_n1007), .C2(new_n765), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n782), .A2(new_n214), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n850), .A2(G159), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G58), .A2(new_n841), .B1(new_n772), .B2(G68), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1001), .A2(G77), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n255), .B1(new_n837), .B2(new_n765), .C1(new_n758), .C2(new_n288), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G143), .B2(new_n753), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1008), .B1(new_n1009), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n794), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n961), .A2(new_n804), .A3(new_n962), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n798), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n805), .B1(new_n231), .B2(new_n391), .C1(new_n1020), .C2(new_n241), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n811), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n996), .A2(new_n1022), .ZN(G387));
  AOI21_X1  g0823(.A(new_n809), .B1(new_n990), .B2(new_n991), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n674), .A2(new_n807), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n540), .A2(new_n772), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n841), .A2(G77), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n288), .B2(new_n765), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT112), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1002), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1027), .B(new_n1031), .C1(new_n1030), .C2(new_n1029), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n797), .B1(new_n749), .B2(new_n224), .C1(new_n293), .C2(new_n761), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G50), .B2(new_n759), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(new_n776), .C2(new_n754), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT113), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n850), .A2(G311), .B1(G322), .B2(new_n753), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n745), .B2(new_n782), .C1(new_n1007), .C2(new_n758), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT48), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n768), .B2(new_n773), .C1(new_n770), .C2(new_n744), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT49), .Z(new_n1041));
  OAI221_X1 g0841(.A(new_n840), .B1(new_n461), .B2(new_n769), .C1(new_n765), .C2(new_n755), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n827), .B(new_n1025), .C1(new_n1043), .C2(new_n794), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n798), .B1(new_n238), .B2(new_n271), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n689), .A2(new_n231), .A3(new_n255), .ZN(new_n1046));
  AOI211_X1 g0846(.A(G45), .B(new_n689), .C1(G68), .C2(G77), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n293), .A2(G50), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1045), .A2(new_n1046), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n231), .A2(G107), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n805), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1024), .B1(new_n1044), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n992), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n990), .A2(new_n739), .A3(new_n991), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n691), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1053), .A2(new_n1056), .ZN(G393));
  NAND3_X1  g0857(.A1(new_n984), .A2(KEYINPUT114), .A3(new_n993), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT114), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n982), .A2(new_n1059), .A3(new_n983), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n691), .B(new_n994), .C1(new_n1061), .C2(new_n992), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n753), .A2(G150), .B1(new_n759), .B2(G159), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT51), .Z(new_n1064));
  NAND2_X1  g0864(.A1(new_n772), .A2(G77), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n850), .A2(G50), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n224), .A2(new_n744), .B1(new_n769), .B2(new_n204), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1067), .B(new_n840), .C1(G143), .C2(new_n766), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n389), .B2(new_n783), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n753), .A2(G317), .B1(new_n759), .B2(G311), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT52), .Z(new_n1072));
  NAND2_X1  g0872(.A1(new_n750), .A2(G294), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n772), .A2(new_n462), .B1(new_n766), .B2(G322), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n841), .A2(G283), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n255), .B(new_n1076), .C1(G303), .C2(new_n850), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1070), .B1(new_n1077), .B2(new_n788), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT116), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n794), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n805), .B1(new_n206), .B2(new_n231), .C1(new_n1020), .C2(new_n248), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n955), .A2(new_n807), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT115), .ZN(new_n1083));
  AND4_X1   g0883(.A1(new_n811), .A2(new_n1080), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1061), .B2(new_n810), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1062), .A2(new_n1085), .ZN(G390));
  NAND4_X1  g0886(.A1(new_n712), .A2(G330), .A3(new_n714), .A4(new_n822), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(new_n929), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n735), .A2(new_n682), .A3(new_n822), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n926), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n929), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n935), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1092), .A2(new_n899), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n935), .B1(new_n927), .B2(new_n1091), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n933), .B2(new_n936), .ZN(new_n1096));
  OAI211_X1 g0896(.A(KEYINPUT117), .B(new_n1088), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n933), .A2(new_n936), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1095), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1088), .A2(KEYINPUT117), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1088), .A2(KEYINPUT117), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1092), .A2(new_n899), .A3(new_n1093), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1097), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n810), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1098), .A2(new_n802), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n856), .A2(new_n293), .ZN(new_n1108));
  INV_X1    g0908(.A(G128), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n754), .A2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT54), .B(G143), .Z(new_n1111));
  AOI22_X1  g0911(.A1(new_n850), .A2(G137), .B1(new_n783), .B2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT120), .ZN(new_n1113));
  OR3_X1    g0913(.A1(new_n744), .A2(KEYINPUT53), .A3(new_n288), .ZN(new_n1114));
  OAI21_X1  g0914(.A(KEYINPUT53), .B1(new_n744), .B2(new_n288), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1114), .B(new_n1115), .C1(new_n214), .C2(new_n769), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n254), .B(new_n1116), .C1(G132), .C2(new_n759), .ZN(new_n1117));
  INV_X1    g0917(.A(G125), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1113), .B(new_n1117), .C1(new_n1118), .C2(new_n765), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1110), .B(new_n1119), .C1(G159), .C2(new_n772), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n254), .B1(new_n765), .B2(new_n770), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n782), .A2(new_n206), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n754), .A2(new_n768), .B1(new_n758), .B2(new_n945), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1122), .A2(new_n1123), .A3(new_n835), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n850), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1065), .C1(new_n210), .C2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1121), .B(new_n1126), .C1(G87), .C2(new_n841), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n794), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1107), .A2(new_n811), .A3(new_n1108), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1106), .A2(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1087), .A2(new_n929), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1087), .A2(new_n929), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n927), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1090), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1087), .A2(new_n929), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1088), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT119), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n716), .A2(new_n457), .A3(G330), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT118), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1088), .A2(new_n1134), .A3(KEYINPUT119), .A4(new_n1135), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(new_n941), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n1097), .A3(new_n1104), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1142), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n695), .B1(new_n1105), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1130), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G378));
  NAND2_X1  g0947(.A1(new_n840), .A2(new_n270), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1028), .B1(new_n768), .B2(new_n765), .C1(new_n758), .C2(new_n210), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n540), .B2(new_n750), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1001), .A2(G58), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n206), .B2(new_n761), .C1(new_n945), .C2(new_n754), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1148), .B(new_n1153), .C1(G68), .C2(new_n772), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT58), .Z(new_n1155));
  NOR2_X1   g0955(.A1(G33), .A2(G41), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT121), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1148), .A2(new_n214), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(G124), .B2(new_n766), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n776), .B2(new_n769), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n761), .A2(new_n843), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1109), .A2(new_n758), .B1(new_n749), .B2(new_n837), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1161), .B(new_n1162), .C1(new_n841), .C2(new_n1111), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n1118), .B2(new_n754), .C1(new_n288), .C2(new_n773), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT59), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1155), .B(new_n1158), .C1(new_n1160), .C2(new_n1165), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1166), .A2(new_n794), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n857), .A2(G50), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n314), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n314), .A2(new_n1170), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n893), .A2(new_n302), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n803), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR4_X1   g0977(.A1(new_n1167), .A2(new_n827), .A3(new_n1168), .A4(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1176), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT122), .B1(new_n1180), .B2(new_n1174), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n911), .A2(new_n915), .A3(new_n919), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n913), .B1(new_n899), .B2(new_n908), .ZN(new_n1183));
  OAI211_X1 g0983(.A(G330), .B(new_n1181), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(G330), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n910), .B2(new_n920), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1181), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1180), .A2(KEYINPUT122), .A3(new_n1174), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1184), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT123), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n938), .A2(KEYINPUT124), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT124), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n931), .A2(new_n937), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1190), .A2(new_n1193), .A3(new_n1191), .A4(new_n1195), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1179), .B1(new_n1199), .B2(new_n809), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1140), .A2(new_n941), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1142), .B1(new_n1097), .B2(new_n1104), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1197), .B(new_n1198), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n695), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1105), .A2(new_n1144), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1201), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n938), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1190), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n938), .B(new_n1184), .C1(new_n1186), .C2(new_n1189), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(KEYINPUT57), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1200), .B1(new_n1205), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(G375));
  AOI22_X1  g1014(.A1(new_n759), .A2(G137), .B1(G159), .B2(new_n841), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1215), .B(new_n797), .C1(new_n843), .C2(new_n754), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n850), .B2(new_n1111), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1151), .B1(new_n1109), .B2(new_n765), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1217), .B(new_n1219), .C1(new_n288), .C2(new_n749), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G50), .B2(new_n772), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n850), .A2(new_n462), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n783), .A2(G107), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1012), .A2(new_n254), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT125), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n841), .A2(G97), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n758), .A2(new_n768), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n765), .A2(new_n745), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1026), .B1(new_n754), .B2(new_n770), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n794), .B1(new_n1221), .B2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n811), .B(new_n1232), .C1(new_n1091), .C2(new_n803), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n224), .B2(new_n856), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1235), .B2(new_n810), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n971), .B1(new_n1235), .B2(new_n1207), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(new_n1144), .ZN(G381));
  NAND4_X1  g1038(.A1(new_n996), .A2(new_n1062), .A3(new_n1022), .A4(new_n1085), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(G375), .A2(G378), .A3(G381), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G384), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(G393), .A2(G396), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(G407));
  NAND2_X1  g1043(.A1(new_n666), .A2(G213), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT126), .Z(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1213), .A2(new_n1146), .A3(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(G407), .A2(G213), .A3(new_n1247), .ZN(G409));
  AND2_X1   g1048(.A1(G393), .A2(G396), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(new_n1242), .ZN(new_n1250));
  AND4_X1   g1050(.A1(new_n996), .A2(new_n1062), .A3(new_n1022), .A4(new_n1085), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n996), .A2(new_n1022), .B1(new_n1062), .B2(new_n1085), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(G390), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1250), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1255), .A3(new_n1239), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT60), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1235), .B2(new_n1207), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n691), .A3(new_n1142), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1235), .A2(new_n1207), .A3(new_n1258), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1236), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1241), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G384), .B(new_n1236), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1146), .B(new_n1200), .C1(new_n1205), .C2(new_n1212), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1210), .A2(new_n1211), .A3(new_n810), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1179), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1208), .A2(new_n971), .A3(new_n1198), .A4(new_n1197), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT127), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1268), .A2(new_n1272), .A3(new_n1179), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1274), .A2(new_n1146), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1244), .B(new_n1266), .C1(new_n1267), .C2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n691), .A3(new_n1212), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1200), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(G378), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1274), .A2(new_n1146), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1246), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1265), .A2(new_n1277), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1276), .A2(new_n1277), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n666), .A2(G213), .A3(G2897), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1266), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1245), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(G2897), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1286), .B1(new_n1291), .B2(new_n1283), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1257), .B1(new_n1285), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT63), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1265), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1257), .B1(new_n1283), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1244), .B1(new_n1267), .B2(new_n1275), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1266), .A2(new_n1287), .B1(new_n1289), .B2(G2897), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1294), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1276), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1286), .B(new_n1296), .C1(new_n1299), .C2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1293), .A2(new_n1301), .ZN(G405));
  NOR2_X1   g1102(.A1(new_n1213), .A2(G378), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1303), .A2(new_n1267), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1257), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1304), .A2(new_n1257), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1265), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1304), .A2(new_n1257), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(new_n1266), .A3(new_n1305), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(G402));
endmodule


