//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT91), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT15), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT92), .ZN(new_n208));
  NOR3_X1   g007(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(new_n208), .B2(new_n209), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n205), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  OAI22_X1  g013(.A1(new_n207), .A2(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT15), .A3(new_n202), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(KEYINPUT93), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(KEYINPUT93), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n219), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  AOI21_X1  g023(.A(G1gat), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G8gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(KEYINPUT94), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT95), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n229), .B(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n217), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n230), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n232), .B(new_n233), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n235), .B(KEYINPUT96), .Z(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT13), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n234), .A4(new_n235), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT11), .B(G169gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(G197gat), .ZN(new_n246));
  XOR2_X1   g045(.A(G113gat), .B(G141gat), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n238), .A2(new_n242), .A3(new_n249), .A4(new_n243), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n254));
  INV_X1    g053(.A(G183gat), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT68), .B1(new_n255), .B2(KEYINPUT27), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT27), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(G183gat), .ZN(new_n259));
  INV_X1    g058(.A(G190gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(new_n258), .B2(G183gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n255), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n254), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT69), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n268), .B(new_n254), .C1(new_n261), .C2(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n258), .A2(G183gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT27), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT28), .A4(new_n260), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT26), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(G169gat), .B2(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(KEYINPUT26), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n273), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT23), .ZN(new_n283));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n283), .A2(KEYINPUT65), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT65), .B1(new_n283), .B2(new_n284), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  NOR2_X1   g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n274), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(KEYINPUT24), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n255), .A2(new_n260), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(KEYINPUT24), .A3(new_n292), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(KEYINPUT66), .C1(KEYINPUT24), .C2(new_n292), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n277), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n287), .A2(new_n294), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G176gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n276), .A2(KEYINPUT64), .ZN(new_n304));
  OAI211_X1 g103(.A(KEYINPUT23), .B(new_n275), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  AND4_X1   g104(.A1(new_n301), .A2(new_n305), .A3(new_n284), .A4(new_n299), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n291), .A2(new_n293), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n300), .A2(KEYINPUT25), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n282), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G113gat), .B(G120gat), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT70), .B1(new_n310), .B2(KEYINPUT1), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313));
  INV_X1    g112(.A(G113gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(G120gat), .ZN(new_n315));
  INV_X1    g114(.A(G120gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(G113gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n312), .B(new_n313), .C1(new_n315), .C2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n311), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n320), .B1(new_n311), .B2(new_n318), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n309), .B(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT34), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT33), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G15gat), .B(G43gat), .Z(new_n332));
  XNOR2_X1  g131(.A(G71gat), .B(G99gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT32), .A3(new_n329), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(KEYINPUT32), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(new_n331), .A3(new_n334), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n328), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n328), .B1(new_n336), .B2(new_n338), .ZN(new_n341));
  OR3_X1    g140(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT36), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n336), .A2(new_n338), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT34), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n327), .B(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n343), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n328), .A2(new_n336), .A3(KEYINPUT72), .A4(new_n338), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT36), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n282), .A2(new_n308), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n282), .B2(new_n308), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n273), .A2(new_n281), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n294), .A2(new_n297), .ZN(new_n360));
  INV_X1    g159(.A(new_n286), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n283), .A2(KEYINPUT65), .A3(new_n284), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n299), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT25), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n306), .A2(new_n307), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n358), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT75), .A3(new_n352), .ZN(new_n368));
  XNOR2_X1  g167(.A(G197gat), .B(G204gat), .ZN(new_n369));
  INV_X1    g168(.A(G211gat), .ZN(new_n370));
  INV_X1    g169(.A(G218gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(KEYINPUT22), .B2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G211gat), .B(G218gat), .Z(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT29), .B1(new_n282), .B2(new_n308), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n353), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n357), .A2(new_n368), .A3(new_n375), .A4(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n358), .B(new_n352), .C1(new_n355), .C2(new_n356), .ZN(new_n382));
  INV_X1    g181(.A(new_n375), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n282), .A2(new_n308), .A3(new_n353), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT74), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n382), .A2(KEYINPUT74), .A3(new_n383), .A4(new_n384), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(G8gat), .B(G36gat), .Z(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G64gat), .ZN(new_n391));
  INV_X1    g190(.A(G92gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n381), .A2(KEYINPUT30), .A3(new_n389), .A4(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n387), .A2(new_n388), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT75), .B1(new_n367), .B2(new_n352), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n377), .A2(new_n376), .A3(new_n353), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n399), .A2(new_n380), .A3(new_n375), .A4(new_n357), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n379), .A2(KEYINPUT76), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n393), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n401), .A3(new_n400), .A4(new_n394), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(G148gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(G141gat), .ZN(new_n412));
  INV_X1    g211(.A(G141gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G148gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G155gat), .B(G162gat), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n417));
  INV_X1    g216(.A(G155gat), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT2), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n415), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT78), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT2), .B1(new_n412), .B2(new_n414), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n416), .ZN(new_n423));
  INV_X1    g222(.A(G162gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(G155gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n418), .A2(G162gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G141gat), .B(G148gat), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n427), .B(KEYINPUT78), .C1(new_n428), .C2(KEYINPUT2), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n420), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n430), .B(new_n431), .C1(new_n322), .C2(new_n323), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT82), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n322), .B2(new_n323), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n311), .A2(new_n318), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n319), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n321), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n431), .A4(new_n430), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  AOI211_X1 g241(.A(KEYINPUT3), .B(new_n420), .C1(new_n423), .C2(new_n429), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT3), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n429), .ZN(new_n445));
  INV_X1    g244(.A(new_n420), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT80), .B1(new_n448), .B2(new_n324), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT3), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n430), .A2(new_n444), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(KEYINPUT80), .A3(new_n324), .A4(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n410), .B(new_n442), .C1(new_n449), .C2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n450), .A2(new_n438), .A3(new_n321), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n434), .ZN(new_n458));
  INV_X1    g257(.A(new_n410), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI211_X1 g259(.A(KEYINPUT83), .B(new_n410), .C1(new_n457), .C2(new_n434), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n455), .A2(new_n462), .A3(KEYINPUT5), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT0), .B(G57gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(G85gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n324), .A3(new_n452), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT80), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n453), .ZN(new_n471));
  INV_X1    g270(.A(new_n435), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n434), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT4), .B1(new_n439), .B2(new_n430), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT5), .ZN(new_n475));
  AND4_X1   g274(.A1(KEYINPUT84), .A2(new_n471), .A3(new_n410), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n459), .B1(new_n470), .B2(new_n453), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT84), .B1(new_n477), .B2(new_n475), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n463), .B(new_n467), .C1(new_n476), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT85), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n471), .A2(new_n410), .A3(new_n475), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(KEYINPUT84), .A3(new_n475), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n485), .A2(new_n486), .A3(new_n467), .A4(new_n463), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n463), .B1(new_n476), .B2(new_n478), .ZN(new_n488));
  INV_X1    g287(.A(new_n467), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n480), .A2(new_n487), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n467), .B1(new_n485), .B2(new_n463), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n405), .A2(KEYINPUT77), .A3(new_n406), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n404), .A2(new_n409), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G228gat), .A2(G233gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n375), .A2(new_n358), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n430), .B1(new_n499), .B2(new_n444), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n375), .B1(new_n452), .B2(new_n358), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n502), .B(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n506));
  OR3_X1    g305(.A1(new_n505), .A2(new_n506), .A3(G22gat), .ZN(new_n507));
  XOR2_X1   g306(.A(G78gat), .B(G106gat), .Z(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT31), .B(G50gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n505), .B2(new_n506), .ZN(new_n512));
  OAI21_X1  g311(.A(G22gat), .B1(new_n505), .B2(new_n506), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n507), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n507), .B2(new_n513), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n351), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n519));
  NOR2_X1   g318(.A1(KEYINPUT88), .A2(KEYINPUT40), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n473), .A2(new_n474), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n471), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n459), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n457), .A2(new_n410), .A3(new_n434), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(KEYINPUT39), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT39), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n527), .A3(new_n459), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n528), .A3(new_n467), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n529), .A2(KEYINPUT88), .A3(KEYINPUT40), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(KEYINPUT88), .B2(KEYINPUT40), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n490), .B(new_n521), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n496), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT77), .B1(new_n405), .B2(new_n406), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n532), .B1(new_n535), .B2(new_n404), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n514), .A2(new_n515), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT38), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n389), .A2(new_n401), .A3(new_n400), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(KEYINPUT37), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n389), .A2(new_n541), .A3(new_n401), .A4(new_n400), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n357), .A2(new_n368), .A3(new_n383), .A4(new_n378), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n382), .A2(new_n375), .A3(new_n384), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT37), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n545), .A2(new_n393), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n540), .A2(new_n542), .B1(new_n547), .B2(new_n538), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT38), .B1(new_n381), .B2(new_n389), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n492), .B(new_n494), .C1(new_n549), .C2(new_n393), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n537), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n519), .B1(new_n536), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n393), .B1(new_n539), .B2(new_n538), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n495), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n538), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT37), .B1(new_n396), .B2(new_n402), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(KEYINPUT38), .A3(new_n542), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n516), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n404), .A2(new_n409), .A3(new_n496), .ZN(new_n560));
  NAND2_X1  g359(.A1(KEYINPUT88), .A2(KEYINPUT40), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n529), .B(new_n561), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n562), .A2(new_n493), .A3(new_n520), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n564), .A3(KEYINPUT89), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n518), .B1(new_n552), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT35), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n537), .B(new_n567), .C1(new_n340), .C2(new_n341), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT90), .ZN(new_n569));
  OR3_X1    g368(.A1(new_n497), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n497), .B2(new_n568), .ZN(new_n571));
  INV_X1    g370(.A(new_n560), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n516), .B1(new_n347), .B2(new_n348), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n495), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n570), .A2(new_n571), .B1(new_n574), .B2(KEYINPUT35), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n253), .B1(new_n566), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT97), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT10), .ZN(new_n581));
  XOR2_X1   g380(.A(G57gat), .B(G64gat), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT98), .B1(G71gat), .B2(G78gat), .ZN(new_n585));
  OR3_X1    g384(.A1(KEYINPUT98), .A2(G71gat), .A3(G78gat), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT9), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n589), .A2(KEYINPUT99), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(KEYINPUT99), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n590), .A2(new_n591), .A3(new_n582), .A4(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n598), .B2(new_n392), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G99gat), .ZN(new_n601));
  INV_X1    g400(.A(G106gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n597), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n597), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n596), .A2(new_n606), .A3(new_n599), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n607), .A2(new_n605), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n594), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n587), .A2(new_n593), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n607), .B2(new_n604), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n581), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n609), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT102), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n618), .A3(new_n615), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n580), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n610), .A2(new_n612), .A3(new_n579), .ZN(new_n621));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n276), .ZN(new_n623));
  INV_X1    g422(.A(G204gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n620), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n579), .B(KEYINPUT103), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n616), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n625), .B1(new_n630), .B2(new_n621), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(KEYINPUT97), .B(new_n253), .C1(new_n566), .C2(new_n575), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n578), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n594), .A2(KEYINPUT21), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n594), .A2(KEYINPUT21), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n232), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n255), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G127gat), .B(G155gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(G211gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n643), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n638), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n637), .A3(new_n646), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n222), .A2(new_n609), .A3(new_n608), .ZN(new_n654));
  AND2_X1   g453(.A1(G232gat), .A2(G233gat), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n217), .A2(new_n614), .B1(KEYINPUT41), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G134gat), .B(G162gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT101), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n657), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n655), .A2(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g460(.A(G190gat), .B(G218gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n660), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n653), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n634), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n495), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g469(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n224), .A2(new_n226), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n667), .A2(new_n560), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G8gat), .B1(new_n666), .B2(new_n572), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(G1325gat));
  INV_X1    g477(.A(new_n351), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n667), .A2(G15gat), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n340), .A2(new_n341), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(G15gat), .B1(new_n667), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n680), .A2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n666), .A2(new_n537), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT43), .B(G22gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  AND2_X1   g486(.A1(new_n351), .A2(new_n517), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n559), .A2(new_n564), .A3(KEYINPUT89), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT89), .B1(new_n559), .B2(new_n564), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n692));
  INV_X1    g491(.A(new_n575), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n688), .B(new_n694), .C1(new_n689), .C2(new_n690), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n664), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g498(.A(KEYINPUT44), .B(new_n664), .C1(new_n566), .C2(new_n575), .ZN(new_n700));
  INV_X1    g499(.A(new_n632), .ZN(new_n701));
  INV_X1    g500(.A(new_n253), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n652), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n699), .A2(new_n668), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n700), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n697), .B2(new_n698), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n708), .A2(KEYINPUT105), .A3(new_n668), .A4(new_n703), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n706), .A2(G29gat), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n578), .A2(new_n664), .A3(new_n633), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n652), .A2(new_n701), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n711), .A2(new_n212), .A3(new_n668), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT45), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n578), .A2(new_n664), .A3(new_n633), .A4(new_n712), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n495), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(new_n717), .A3(new_n212), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n710), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n710), .A2(KEYINPUT106), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n560), .A3(new_n703), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n711), .A2(new_n213), .A3(new_n560), .A4(new_n712), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n725), .A2(G36gat), .B1(new_n726), .B2(KEYINPUT46), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n726), .B2(KEYINPUT46), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n715), .A2(G36gat), .A3(new_n572), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(KEYINPUT107), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n727), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n727), .A2(KEYINPUT108), .A3(new_n729), .A4(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(G1329gat));
  NOR3_X1   g536(.A1(new_n715), .A2(G43gat), .A3(new_n681), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n708), .A2(new_n679), .A3(new_n703), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT47), .B1(new_n741), .B2(KEYINPUT109), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n742), .A2(new_n745), .ZN(G1330gat));
  XNOR2_X1  g545(.A(new_n715), .B(KEYINPUT110), .ZN(new_n747));
  INV_X1    g546(.A(G50gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n748), .A3(new_n516), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n708), .A2(new_n516), .A3(new_n703), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G50gat), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n750), .B1(new_n749), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(G1331gat));
  NOR3_X1   g554(.A1(new_n653), .A2(new_n664), .A3(new_n253), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n696), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(new_n701), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n668), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n701), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n572), .B(new_n761), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1333gat));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n758), .A2(new_n765), .A3(new_n682), .ZN(new_n766));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT111), .B1(new_n761), .B2(new_n681), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n758), .A2(G71gat), .A3(new_n679), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT50), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n773), .A3(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n516), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g576(.A(KEYINPUT44), .B1(new_n696), .B2(new_n664), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n652), .A2(new_n253), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n778), .A2(new_n707), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n701), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n782), .A2(new_n598), .A3(new_n495), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n696), .A2(new_n664), .A3(new_n779), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT51), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n696), .A2(new_n786), .A3(new_n664), .A4(new_n779), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(new_n668), .A3(new_n701), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n783), .B1(new_n598), .B2(new_n789), .ZN(G1336gat));
  OAI21_X1  g589(.A(G92gat), .B1(new_n782), .B2(new_n572), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n788), .A2(new_n392), .A3(new_n701), .A4(new_n560), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT52), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n782), .B2(new_n351), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n788), .A2(new_n601), .A3(new_n701), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n681), .B2(new_n799), .ZN(G1338gat));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n701), .A3(new_n516), .A4(new_n787), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n602), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n781), .A2(G106gat), .A3(new_n701), .A4(new_n516), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT112), .ZN(new_n805));
  XNOR2_X1  g604(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(KEYINPUT112), .A3(new_n806), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1339gat));
  NOR2_X1   g609(.A1(new_n239), .A2(new_n241), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n235), .B1(new_n230), .B2(new_n234), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n248), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n252), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n616), .A2(new_n628), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n620), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n625), .B1(new_n629), .B2(KEYINPUT54), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n626), .B1(new_n819), .B2(KEYINPUT55), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n817), .B2(new_n818), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n664), .A2(new_n814), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n253), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n814), .A2(new_n701), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n664), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n653), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n664), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n652), .A2(new_n830), .A3(new_n632), .A4(new_n702), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(new_n573), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n560), .A2(new_n495), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT114), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n314), .A3(new_n253), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n681), .A2(new_n516), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n839), .A2(new_n834), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n702), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n837), .A2(new_n842), .ZN(G1340gat));
  NAND3_X1  g642(.A1(new_n836), .A2(new_n316), .A3(new_n701), .ZN(new_n844));
  OAI21_X1  g643(.A(G120gat), .B1(new_n841), .B2(new_n632), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1341gat));
  NAND3_X1  g645(.A1(new_n840), .A2(G127gat), .A3(new_n652), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT115), .ZN(new_n848));
  AOI21_X1  g647(.A(G127gat), .B1(new_n835), .B2(new_n652), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n851), .A3(new_n664), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(KEYINPUT56), .Z(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n841), .B2(new_n830), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n822), .A2(KEYINPUT116), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n857), .B(new_n821), .C1(new_n817), .C2(new_n818), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n820), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n820), .A2(new_n856), .A3(KEYINPUT117), .A4(new_n858), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n253), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n664), .B1(new_n863), .B2(new_n827), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n653), .B1(new_n864), .B2(new_n825), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n831), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n516), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT57), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n537), .B1(new_n829), .B2(new_n831), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n351), .A2(new_n834), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G141gat), .B1(new_n874), .B2(new_n702), .ZN(new_n875));
  INV_X1    g674(.A(new_n869), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n872), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n413), .A3(new_n253), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n411), .A3(new_n701), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  INV_X1    g681(.A(new_n828), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n652), .B1(new_n883), .B2(new_n824), .ZN(new_n884));
  AND4_X1   g683(.A1(new_n652), .A2(new_n830), .A3(new_n632), .A4(new_n702), .ZN(new_n885));
  OAI211_X1 g684(.A(KEYINPUT57), .B(new_n516), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT118), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n869), .A2(new_n888), .A3(KEYINPUT57), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT119), .B1(new_n867), .B2(new_n870), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n537), .B1(new_n865), .B2(new_n831), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT57), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n701), .A3(new_n873), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n411), .B1(new_n896), .B2(KEYINPUT120), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n895), .A2(new_n898), .A3(new_n701), .A4(new_n873), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n882), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n874), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT59), .B(new_n411), .C1(new_n901), .C2(new_n701), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n881), .B1(new_n900), .B2(new_n902), .ZN(G1345gat));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n652), .ZN(new_n904));
  XNOR2_X1  g703(.A(KEYINPUT79), .B(G155gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n653), .A2(new_n905), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n904), .A2(new_n905), .B1(new_n877), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT121), .ZN(G1346gat));
  AOI21_X1  g707(.A(G162gat), .B1(new_n877), .B2(new_n664), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n874), .A2(new_n424), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n664), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n572), .A2(new_n668), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n833), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n275), .A3(new_n253), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n832), .A2(new_n838), .A3(new_n912), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT122), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(KEYINPUT122), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n253), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n914), .B1(new_n919), .B2(new_n275), .ZN(G1348gat));
  AOI21_X1  g719(.A(G176gat), .B1(new_n913), .B2(new_n701), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n632), .A2(new_n303), .A3(new_n304), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n918), .B2(new_n922), .ZN(G1349gat));
  NAND3_X1  g722(.A1(new_n916), .A2(new_n652), .A3(new_n917), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT123), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n916), .A2(new_n926), .A3(new_n652), .A4(new_n917), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(G183gat), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n652), .A3(new_n270), .A4(new_n271), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g730(.A(new_n260), .B1(new_n918), .B2(new_n664), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n932), .A2(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(KEYINPUT61), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n913), .A2(new_n260), .A3(new_n664), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT124), .Z(new_n936));
  NAND3_X1  g735(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(G1351gat));
  NAND2_X1  g736(.A1(new_n912), .A2(new_n351), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n876), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT125), .Z(new_n940));
  INV_X1    g739(.A(G197gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n941), .A3(new_n253), .ZN(new_n942));
  INV_X1    g741(.A(new_n895), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(new_n702), .A3(new_n938), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n942), .B1(new_n944), .B2(new_n941), .ZN(G1352gat));
  NAND2_X1  g744(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n939), .A2(new_n624), .A3(new_n701), .A4(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n943), .A2(new_n632), .A3(new_n938), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n624), .ZN(G1353gat));
  NAND4_X1  g750(.A1(new_n895), .A2(new_n652), .A3(new_n351), .A4(new_n912), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G211gat), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT63), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n370), .A3(new_n652), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(KEYINPUT63), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n954), .A2(KEYINPUT63), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n952), .A2(G211gat), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n956), .A3(new_n959), .ZN(G1354gat));
  NAND3_X1  g759(.A1(new_n940), .A2(new_n371), .A3(new_n664), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n943), .A2(new_n830), .A3(new_n938), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n371), .ZN(G1355gat));
endmodule


