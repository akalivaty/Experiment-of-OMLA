

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590;

  XNOR2_X1 U323 ( .A(n417), .B(n416), .ZN(n543) );
  XNOR2_X1 U324 ( .A(n415), .B(KEYINPUT48), .ZN(n416) );
  XOR2_X1 U325 ( .A(KEYINPUT97), .B(n462), .Z(n291) );
  INV_X1 U326 ( .A(G92GAT), .ZN(n315) );
  XNOR2_X1 U327 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n418) );
  XNOR2_X1 U328 ( .A(n340), .B(n451), .ZN(n341) );
  XNOR2_X1 U329 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U330 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U331 ( .A(n342), .B(n341), .ZN(n344) );
  XNOR2_X1 U332 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U333 ( .A(n325), .B(n432), .Z(n519) );
  XNOR2_X1 U334 ( .A(n456), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U335 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U336 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n482), .B(n481), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(G127GAT), .B(G134GAT), .Z(n293) );
  XNOR2_X1 U339 ( .A(G120GAT), .B(KEYINPUT0), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n308) );
  XOR2_X1 U341 ( .A(G155GAT), .B(KEYINPUT2), .Z(n295) );
  XNOR2_X1 U342 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n429) );
  XOR2_X1 U344 ( .A(G85GAT), .B(n429), .Z(n297) );
  XOR2_X1 U345 ( .A(G113GAT), .B(G1GAT), .Z(n346) );
  XNOR2_X1 U346 ( .A(G29GAT), .B(n346), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U348 ( .A(G57GAT), .B(KEYINPUT1), .Z(n299) );
  NAND2_X1 U349 ( .A1(G225GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U351 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U352 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n303) );
  XNOR2_X1 U353 ( .A(G141GAT), .B(G148GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n304), .B(KEYINPUT4), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n545) );
  INV_X1 U358 ( .A(n545), .ZN(n517) );
  XOR2_X1 U359 ( .A(KEYINPUT80), .B(KEYINPUT95), .Z(n310) );
  XNOR2_X1 U360 ( .A(G190GAT), .B(G204GAT), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n320) );
  XOR2_X1 U362 ( .A(G176GAT), .B(G64GAT), .Z(n333) );
  XOR2_X1 U363 ( .A(G183GAT), .B(KEYINPUT17), .Z(n312) );
  XNOR2_X1 U364 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n440) );
  XOR2_X1 U366 ( .A(n333), .B(n440), .Z(n314) );
  NAND2_X1 U367 ( .A1(G226GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U369 ( .A(G169GAT), .B(G8GAT), .Z(n345) );
  XNOR2_X1 U370 ( .A(G36GAT), .B(n345), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n325) );
  XOR2_X1 U372 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n322) );
  XNOR2_X1 U373 ( .A(G197GAT), .B(G211GAT), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U375 ( .A(G218GAT), .B(KEYINPUT21), .Z(n323) );
  XOR2_X1 U376 ( .A(n324), .B(n323), .Z(n432) );
  XOR2_X1 U377 ( .A(G92GAT), .B(KEYINPUT75), .Z(n327) );
  XNOR2_X1 U378 ( .A(G99GAT), .B(G85GAT), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n389) );
  XNOR2_X1 U380 ( .A(n389), .B(KEYINPUT32), .ZN(n330) );
  INV_X1 U381 ( .A(n330), .ZN(n329) );
  INV_X1 U382 ( .A(KEYINPUT76), .ZN(n328) );
  NAND2_X1 U383 ( .A1(n329), .A2(n328), .ZN(n332) );
  NAND2_X1 U384 ( .A1(n330), .A2(KEYINPUT76), .ZN(n331) );
  NAND2_X1 U385 ( .A1(n332), .A2(n331), .ZN(n336) );
  XNOR2_X1 U386 ( .A(n333), .B(KEYINPUT33), .ZN(n334) );
  XOR2_X1 U387 ( .A(n334), .B(KEYINPUT31), .Z(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n342) );
  XOR2_X1 U389 ( .A(G78GAT), .B(G148GAT), .Z(n338) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(G204GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n431) );
  XNOR2_X1 U392 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n339), .B(KEYINPUT13), .ZN(n372) );
  XNOR2_X1 U394 ( .A(n431), .B(n372), .ZN(n340) );
  XOR2_X1 U395 ( .A(G120GAT), .B(G71GAT), .Z(n451) );
  AND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n410) );
  XNOR2_X1 U398 ( .A(n410), .B(KEYINPUT41), .ZN(n550) );
  XOR2_X1 U399 ( .A(G197GAT), .B(G15GAT), .Z(n348) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U402 ( .A(G141GAT), .B(G22GAT), .Z(n426) );
  XOR2_X1 U403 ( .A(n349), .B(n426), .Z(n354) );
  XOR2_X1 U404 ( .A(KEYINPUT67), .B(KEYINPUT72), .Z(n351) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U407 ( .A(KEYINPUT29), .B(n352), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n364) );
  XOR2_X1 U409 ( .A(G43GAT), .B(G29GAT), .Z(n356) );
  XNOR2_X1 U410 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U412 ( .A(n357), .B(KEYINPUT70), .Z(n359) );
  XNOR2_X1 U413 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n402) );
  XOR2_X1 U415 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n361) );
  XNOR2_X1 U416 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U418 ( .A(n402), .B(n362), .Z(n363) );
  XOR2_X1 U419 ( .A(n364), .B(n363), .Z(n576) );
  INV_X1 U420 ( .A(n576), .ZN(n546) );
  AND2_X1 U421 ( .A1(n550), .A2(n546), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n365), .B(KEYINPUT46), .ZN(n387) );
  XOR2_X1 U423 ( .A(G15GAT), .B(G127GAT), .Z(n438) );
  XOR2_X1 U424 ( .A(G155GAT), .B(G78GAT), .Z(n367) );
  XNOR2_X1 U425 ( .A(G71GAT), .B(G183GAT), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U427 ( .A(n438), .B(n368), .Z(n370) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n371), .B(KEYINPUT84), .ZN(n374) );
  XOR2_X1 U431 ( .A(n372), .B(KEYINPUT85), .Z(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U433 ( .A(G64GAT), .B(G211GAT), .Z(n376) );
  XNOR2_X1 U434 ( .A(G22GAT), .B(G1GAT), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n386) );
  XOR2_X1 U437 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n380) );
  XNOR2_X1 U438 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U440 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n382) );
  XNOR2_X1 U441 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U443 ( .A(n384), .B(n383), .Z(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n570) );
  NOR2_X1 U445 ( .A1(n387), .A2(n570), .ZN(n403) );
  INV_X1 U446 ( .A(G162GAT), .ZN(n388) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U448 ( .A(G190GAT), .B(G134GAT), .Z(n439) );
  XNOR2_X1 U449 ( .A(n439), .B(G218GAT), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U451 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n393) );
  NAND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n392) );
  XOR2_X1 U453 ( .A(n393), .B(n392), .Z(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n400) );
  XOR2_X1 U455 ( .A(KEYINPUT79), .B(KEYINPUT9), .Z(n397) );
  XNOR2_X1 U456 ( .A(KEYINPUT10), .B(KEYINPUT77), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U458 ( .A(G106GAT), .B(n398), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U460 ( .A(n402), .B(n401), .Z(n556) );
  INV_X1 U461 ( .A(n556), .ZN(n405) );
  NAND2_X1 U462 ( .A1(n403), .A2(n405), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n404), .B(KEYINPUT47), .ZN(n414) );
  INV_X1 U464 ( .A(KEYINPUT65), .ZN(n409) );
  XOR2_X1 U465 ( .A(n405), .B(KEYINPUT36), .Z(n586) );
  NAND2_X1 U466 ( .A1(n570), .A2(n586), .ZN(n407) );
  XOR2_X1 U467 ( .A(KEYINPUT111), .B(KEYINPUT45), .Z(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n412) );
  XOR2_X1 U470 ( .A(KEYINPUT73), .B(n576), .Z(n561) );
  NAND2_X1 U471 ( .A1(n410), .A2(n561), .ZN(n411) );
  NOR2_X1 U472 ( .A1(n412), .A2(n411), .ZN(n413) );
  NOR2_X1 U473 ( .A1(n414), .A2(n413), .ZN(n417) );
  XOR2_X1 U474 ( .A(KEYINPUT64), .B(KEYINPUT112), .Z(n415) );
  NAND2_X1 U475 ( .A1(n519), .A2(n543), .ZN(n419) );
  NOR2_X1 U476 ( .A1(n517), .A2(n420), .ZN(n575) );
  XOR2_X1 U477 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n422) );
  XNOR2_X1 U478 ( .A(KEYINPUT91), .B(KEYINPUT89), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n436) );
  XOR2_X1 U480 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n424) );
  XNOR2_X1 U481 ( .A(G50GAT), .B(KEYINPUT24), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U483 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U486 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n468) );
  NAND2_X1 U490 ( .A1(n575), .A2(n468), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n437), .B(KEYINPUT55), .ZN(n455) );
  XNOR2_X1 U492 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U494 ( .A(G113GAT), .B(KEYINPUT0), .Z(n443) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U497 ( .A(n445), .B(n444), .Z(n450) );
  XOR2_X1 U498 ( .A(G176GAT), .B(KEYINPUT88), .Z(n447) );
  XNOR2_X1 U499 ( .A(KEYINPUT87), .B(KEYINPUT20), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(n448), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U503 ( .A(n452), .B(n451), .Z(n454) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G99GAT), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(n526) );
  NAND2_X1 U506 ( .A1(n455), .A2(n526), .ZN(n571) );
  NOR2_X1 U507 ( .A1(n571), .A2(n405), .ZN(n458) );
  INV_X1 U508 ( .A(G190GAT), .ZN(n456) );
  XOR2_X1 U509 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n459) );
  XNOR2_X1 U510 ( .A(n468), .B(n459), .ZN(n522) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n519), .Z(n470) );
  NOR2_X1 U512 ( .A1(n522), .A2(n470), .ZN(n460) );
  NAND2_X1 U513 ( .A1(n517), .A2(n460), .ZN(n528) );
  XNOR2_X1 U514 ( .A(KEYINPUT96), .B(n528), .ZN(n461) );
  NOR2_X1 U515 ( .A1(n526), .A2(n461), .ZN(n462) );
  XOR2_X1 U516 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n466) );
  NAND2_X1 U517 ( .A1(n526), .A2(n519), .ZN(n463) );
  XOR2_X1 U518 ( .A(KEYINPUT99), .B(n463), .Z(n464) );
  NAND2_X1 U519 ( .A1(n464), .A2(n468), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U521 ( .A(KEYINPUT25), .B(n467), .ZN(n472) );
  NOR2_X1 U522 ( .A1(n526), .A2(n468), .ZN(n469) );
  XOR2_X1 U523 ( .A(KEYINPUT26), .B(n469), .Z(n573) );
  NOR2_X1 U524 ( .A1(n573), .A2(n470), .ZN(n542) );
  XNOR2_X1 U525 ( .A(n542), .B(KEYINPUT98), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U527 ( .A1(n517), .A2(n473), .ZN(n474) );
  NOR2_X1 U528 ( .A1(n291), .A2(n474), .ZN(n485) );
  NOR2_X1 U529 ( .A1(n570), .A2(n485), .ZN(n475) );
  NAND2_X1 U530 ( .A1(n586), .A2(n475), .ZN(n476) );
  XOR2_X1 U531 ( .A(KEYINPUT37), .B(n476), .Z(n515) );
  INV_X1 U532 ( .A(n561), .ZN(n529) );
  NAND2_X1 U533 ( .A1(n410), .A2(n529), .ZN(n488) );
  NOR2_X1 U534 ( .A1(n515), .A2(n488), .ZN(n478) );
  XNOR2_X1 U535 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(n501) );
  NAND2_X1 U537 ( .A1(n501), .A2(n526), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n480) );
  XNOR2_X1 U539 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n490) );
  XOR2_X1 U541 ( .A(KEYINPUT16), .B(KEYINPUT86), .Z(n484) );
  NAND2_X1 U542 ( .A1(n570), .A2(n405), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n487) );
  INV_X1 U544 ( .A(n485), .ZN(n486) );
  NAND2_X1 U545 ( .A1(n487), .A2(n486), .ZN(n505) );
  NOR2_X1 U546 ( .A1(n488), .A2(n505), .ZN(n496) );
  NAND2_X1 U547 ( .A1(n517), .A2(n496), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1324GAT) );
  NAND2_X1 U549 ( .A1(n519), .A2(n496), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n493) );
  NAND2_X1 U552 ( .A1(n496), .A2(n526), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n495) );
  XOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT102), .Z(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n496), .A2(n522), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  NAND2_X1 U559 ( .A1(n501), .A2(n517), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n519), .A2(n501), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT107), .Z(n503) );
  NAND2_X1 U564 ( .A1(n501), .A2(n522), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  INV_X1 U567 ( .A(n550), .ZN(n564) );
  NOR2_X1 U568 ( .A1(n564), .A2(n546), .ZN(n504) );
  XOR2_X1 U569 ( .A(KEYINPUT108), .B(n504), .Z(n516) );
  NOR2_X1 U570 ( .A1(n516), .A2(n505), .ZN(n511) );
  NAND2_X1 U571 ( .A1(n517), .A2(n511), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n519), .A2(n511), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT109), .Z(n510) );
  NAND2_X1 U576 ( .A1(n511), .A2(n526), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n510), .B(n509), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U579 ( .A1(n511), .A2(n522), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n517), .A2(n523), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n523), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n526), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT113), .Z(n531) );
  NAND2_X1 U593 ( .A1(n526), .A2(n543), .ZN(n527) );
  NOR2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n539), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U598 ( .A1(n539), .A2(n550), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n539), .A2(n570), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(KEYINPUT114), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U607 ( .A1(n539), .A2(n556), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n557), .A2(n546), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n549) );
  XNOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n554) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n557), .A2(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n557), .A2(n570), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n571), .A2(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT123), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NOR2_X1 U629 ( .A1(n571), .A2(n564), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n566) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  INV_X1 U635 ( .A(n570), .ZN(n583) );
  NOR2_X1 U636 ( .A1(n583), .A2(n571), .ZN(n572) );
  XOR2_X1 U637 ( .A(G183GAT), .B(n572), .Z(G1350GAT) );
  INV_X1 U638 ( .A(n573), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n585) );
  NOR2_X1 U640 ( .A1(n576), .A2(n585), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n410), .A2(n585), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n589) );
  INV_X1 U651 ( .A(n585), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

