

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775;

  INV_X1 U371 ( .A(n636), .ZN(n349) );
  XOR2_X1 U372 ( .A(G143), .B(G122), .Z(n568) );
  NAND2_X2 U373 ( .A1(n596), .A2(n694), .ZN(n348) );
  XNOR2_X2 U374 ( .A(n348), .B(KEYINPUT92), .ZN(n433) );
  NOR2_X2 U375 ( .A1(n653), .A2(n455), .ZN(n454) );
  XNOR2_X2 U376 ( .A(n640), .B(n639), .ZN(n429) );
  NAND2_X2 U377 ( .A1(n774), .A2(n675), .ZN(n474) );
  XNOR2_X2 U378 ( .A(n462), .B(KEYINPUT32), .ZN(n774) );
  XNOR2_X2 U379 ( .A(n632), .B(KEYINPUT66), .ZN(n633) );
  AND2_X2 U380 ( .A1(n350), .A2(n349), .ZN(n640) );
  XNOR2_X1 U381 ( .A(n634), .B(n351), .ZN(n350) );
  INV_X1 U382 ( .A(n635), .ZN(n351) );
  NOR2_X1 U383 ( .A1(n682), .A2(n684), .ZN(n697) );
  XNOR2_X1 U384 ( .A(G113), .B(G104), .ZN(n567) );
  XNOR2_X1 U385 ( .A(n557), .B(n445), .ZN(n759) );
  XOR2_X1 U386 ( .A(G122), .B(KEYINPUT7), .Z(n560) );
  NOR2_X1 U387 ( .A1(n622), .A2(n601), .ZN(n684) );
  BUF_X1 U388 ( .A(G110), .Z(n398) );
  XNOR2_X1 U389 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n352) );
  XOR2_X1 U390 ( .A(KEYINPUT48), .B(KEYINPUT89), .Z(n353) );
  XNOR2_X2 U391 ( .A(n528), .B(G469), .ZN(n602) );
  XNOR2_X2 U392 ( .A(n461), .B(n633), .ZN(n644) );
  NOR2_X1 U393 ( .A1(n691), .A2(n508), .ZN(n692) );
  AND2_X1 U394 ( .A1(n364), .A2(n418), .ZN(n373) );
  NOR2_X1 U395 ( .A1(n609), .A2(n706), .ZN(n610) );
  INV_X1 U396 ( .A(n646), .ZN(n707) );
  XNOR2_X1 U397 ( .A(n503), .B(G472), .ZN(n660) );
  INV_X1 U398 ( .A(n373), .ZN(n368) );
  INV_X1 U399 ( .A(n600), .ZN(n682) );
  NAND2_X1 U400 ( .A1(n622), .A2(n601), .ZN(n600) );
  AND2_X2 U401 ( .A1(n359), .A2(n358), .ZN(n438) );
  AND2_X1 U402 ( .A1(n368), .A2(G478), .ZN(n356) );
  NAND2_X1 U403 ( .A1(n360), .A2(n368), .ZN(n359) );
  NOR2_X1 U404 ( .A1(n429), .A2(KEYINPUT44), .ZN(n652) );
  NOR2_X1 U405 ( .A1(n611), .A2(n602), .ZN(n375) );
  NOR2_X1 U406 ( .A1(n539), .A2(n629), .ZN(n385) );
  XNOR2_X1 U407 ( .A(n759), .B(G146), .ZN(n532) );
  INV_X1 U408 ( .A(KEYINPUT21), .ZN(n383) );
  INV_X1 U409 ( .A(KEYINPUT38), .ZN(n366) );
  INV_X1 U410 ( .A(G472), .ZN(n369) );
  INV_X1 U411 ( .A(G137), .ZN(n446) );
  INV_X1 U412 ( .A(KEYINPUT46), .ZN(n380) );
  INV_X1 U413 ( .A(G116), .ZN(n485) );
  INV_X1 U414 ( .A(G210), .ZN(n363) );
  INV_X1 U415 ( .A(KEYINPUT69), .ZN(n382) );
  NAND2_X1 U416 ( .A1(n357), .A2(G469), .ZN(n735) );
  INV_X1 U417 ( .A(n359), .ZN(n357) );
  NAND2_X1 U418 ( .A1(n692), .A2(n388), .ZN(n387) );
  NAND2_X1 U419 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U420 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U421 ( .A1(n413), .A2(KEYINPUT87), .ZN(n390) );
  NAND2_X1 U422 ( .A1(n413), .A2(n395), .ZN(n394) );
  NOR2_X1 U423 ( .A1(n378), .A2(n448), .ZN(n377) );
  XNOR2_X1 U424 ( .A(n381), .B(n380), .ZN(n379) );
  NAND2_X1 U425 ( .A1(n775), .A2(n772), .ZN(n381) );
  XNOR2_X1 U426 ( .A(n615), .B(KEYINPUT86), .ZN(n378) );
  AND2_X1 U427 ( .A1(n457), .A2(n706), .ZN(n671) );
  XNOR2_X1 U428 ( .A(n361), .B(n352), .ZN(n775) );
  NOR2_X1 U429 ( .A1(n722), .A2(n362), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n502), .B(n501), .ZN(n772) );
  INV_X1 U431 ( .A(n375), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n488), .B(n415), .ZN(n693) );
  AND2_X1 U433 ( .A1(n499), .A2(n496), .ZN(n411) );
  AND2_X1 U434 ( .A1(n450), .A2(n365), .ZN(n623) );
  AND2_X1 U435 ( .A1(n708), .A2(n486), .ZN(n487) );
  XNOR2_X1 U436 ( .A(KEYINPUT103), .B(n643), .ZN(n645) );
  XNOR2_X1 U437 ( .A(n604), .B(n382), .ZN(n556) );
  AND2_X1 U438 ( .A1(n384), .A2(n702), .ZN(n604) );
  XNOR2_X1 U439 ( .A(n619), .B(n366), .ZN(n365) );
  XNOR2_X1 U440 ( .A(n602), .B(KEYINPUT1), .ZN(n646) );
  XNOR2_X1 U441 ( .A(n385), .B(KEYINPUT81), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n555), .B(n483), .ZN(n648) );
  OR2_X1 U443 ( .A1(n667), .A2(G902), .ZN(n503) );
  XNOR2_X1 U444 ( .A(n577), .B(n430), .ZN(n621) );
  XNOR2_X1 U445 ( .A(n532), .B(n504), .ZN(n667) );
  XNOR2_X1 U446 ( .A(n532), .B(n493), .ZN(n732) );
  NAND2_X1 U447 ( .A1(n404), .A2(G475), .ZN(n420) );
  XNOR2_X1 U448 ( .A(n541), .B(n383), .ZN(n702) );
  XNOR2_X1 U449 ( .A(n583), .B(n447), .ZN(n557) );
  XNOR2_X1 U450 ( .A(n386), .B(KEYINPUT20), .ZN(n552) );
  NAND2_X1 U451 ( .A1(n522), .A2(n521), .ZN(n583) );
  NAND2_X1 U452 ( .A1(n592), .A2(G214), .ZN(n694) );
  INV_X1 U453 ( .A(n664), .ZN(n540) );
  NAND2_X1 U454 ( .A1(n664), .A2(G234), .ZN(n386) );
  XNOR2_X1 U455 ( .A(n516), .B(KEYINPUT94), .ZN(n664) );
  XNOR2_X1 U456 ( .A(n587), .B(n446), .ZN(n445) );
  NAND2_X1 U457 ( .A1(n727), .A2(n395), .ZN(n389) );
  NAND2_X1 U458 ( .A1(n727), .A2(KEYINPUT87), .ZN(n393) );
  INV_X1 U459 ( .A(KEYINPUT16), .ZN(n471) );
  XNOR2_X1 U460 ( .A(G113), .B(G101), .ZN(n533) );
  INV_X1 U461 ( .A(KEYINPUT22), .ZN(n464) );
  INV_X1 U462 ( .A(G128), .ZN(n519) );
  INV_X1 U463 ( .A(G143), .ZN(n520) );
  XOR2_X1 U464 ( .A(G131), .B(G140), .Z(n575) );
  XOR2_X1 U465 ( .A(G125), .B(G146), .Z(n588) );
  XNOR2_X1 U466 ( .A(G119), .B(G137), .ZN(n542) );
  XNOR2_X1 U467 ( .A(G902), .B(KEYINPUT15), .ZN(n516) );
  XOR2_X1 U468 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n635) );
  XNOR2_X1 U469 ( .A(n354), .B(n468), .ZN(n456) );
  NAND2_X1 U470 ( .A1(n469), .A2(n399), .ZN(n354) );
  NAND2_X1 U471 ( .A1(n355), .A2(n360), .ZN(n742) );
  AND2_X1 U472 ( .A1(n368), .A2(G217), .ZN(n355) );
  NAND2_X1 U473 ( .A1(n356), .A2(n360), .ZN(n739) );
  INV_X1 U474 ( .A(n404), .ZN(n358) );
  NOR2_X1 U475 ( .A1(n737), .A2(n745), .ZN(G54) );
  NOR2_X1 U476 ( .A1(n744), .A2(n745), .ZN(G66) );
  NAND2_X1 U477 ( .A1(n367), .A2(n360), .ZN(n437) );
  INV_X2 U478 ( .A(n691), .ZN(n360) );
  INV_X1 U479 ( .A(n722), .ZN(n714) );
  NAND2_X1 U480 ( .A1(n492), .A2(n750), .ZN(n364) );
  NOR2_X1 U481 ( .A1(n373), .A2(n363), .ZN(n371) );
  NAND2_X1 U482 ( .A1(n411), .A2(n365), .ZN(n620) );
  NAND2_X1 U483 ( .A1(n365), .A2(n694), .ZN(n452) );
  NOR2_X1 U484 ( .A1(n365), .A2(n694), .ZN(n695) );
  NOR2_X1 U485 ( .A1(n373), .A2(n420), .ZN(n367) );
  XNOR2_X2 U486 ( .A(n374), .B(n513), .ZN(n691) );
  NOR2_X1 U487 ( .A1(n373), .A2(n369), .ZN(n370) );
  NAND2_X1 U488 ( .A1(n370), .A2(n372), .ZN(n494) );
  NAND2_X1 U489 ( .A1(n371), .A2(n372), .ZN(n491) );
  INV_X1 U490 ( .A(n691), .ZN(n372) );
  NAND2_X1 U491 ( .A1(n750), .A2(n410), .ZN(n374) );
  XNOR2_X2 U492 ( .A(n453), .B(KEYINPUT45), .ZN(n750) );
  NAND2_X1 U493 ( .A1(n375), .A2(n612), .ZN(n616) );
  XNOR2_X1 U494 ( .A(n376), .B(n353), .ZN(n624) );
  NAND2_X1 U495 ( .A1(n379), .A2(n377), .ZN(n376) );
  INV_X1 U496 ( .A(n702), .ZN(n642) );
  NAND2_X1 U497 ( .A1(n391), .A2(n387), .ZN(n444) );
  NAND2_X1 U498 ( .A1(n396), .A2(n392), .ZN(n391) );
  INV_X1 U499 ( .A(KEYINPUT87), .ZN(n395) );
  INV_X1 U500 ( .A(n692), .ZN(n396) );
  BUF_X1 U501 ( .A(n429), .Z(n397) );
  NAND2_X1 U502 ( .A1(n442), .A2(n439), .ZN(n440) );
  XNOR2_X1 U503 ( .A(n474), .B(KEYINPUT91), .ZN(n399) );
  XNOR2_X1 U504 ( .A(n474), .B(n649), .ZN(n400) );
  XNOR2_X1 U505 ( .A(n470), .B(n591), .ZN(n731) );
  XNOR2_X1 U506 ( .A(n754), .B(n583), .ZN(n470) );
  BUF_X1 U507 ( .A(n654), .Z(n401) );
  BUF_X1 U508 ( .A(n774), .Z(n402) );
  BUF_X1 U509 ( .A(n731), .Z(n403) );
  NAND2_X1 U510 ( .A1(n498), .A2(n604), .ZN(n497) );
  INV_X1 U511 ( .A(n648), .ZN(n498) );
  INV_X1 U512 ( .A(n687), .ZN(n449) );
  INV_X1 U513 ( .A(KEYINPUT67), .ZN(n441) );
  XNOR2_X1 U514 ( .A(G101), .B(KEYINPUT97), .ZN(n524) );
  BUF_X1 U515 ( .A(n693), .Z(n723) );
  NOR2_X1 U516 ( .A1(n696), .A2(n451), .ZN(n450) );
  XNOR2_X1 U517 ( .A(G116), .B(G107), .ZN(n562) );
  INV_X1 U518 ( .A(KEYINPUT9), .ZN(n473) );
  INV_X1 U519 ( .A(G134), .ZN(n447) );
  INV_X1 U520 ( .A(KEYINPUT76), .ZN(n513) );
  XNOR2_X1 U521 ( .A(n620), .B(KEYINPUT39), .ZN(n625) );
  XNOR2_X1 U522 ( .A(n553), .B(n484), .ZN(n483) );
  XNOR2_X1 U523 ( .A(n554), .B(KEYINPUT25), .ZN(n484) );
  NAND2_X1 U524 ( .A1(n431), .A2(KEYINPUT118), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n712), .B(KEYINPUT113), .ZN(n481) );
  INV_X1 U526 ( .A(n713), .ZN(n480) );
  INV_X1 U527 ( .A(KEYINPUT71), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n479), .B(n477), .ZN(n715) );
  XNOR2_X1 U529 ( .A(n478), .B(KEYINPUT114), .ZN(n477) );
  NAND2_X1 U530 ( .A1(n481), .A2(n480), .ZN(n479) );
  INV_X1 U531 ( .A(KEYINPUT51), .ZN(n478) );
  NOR2_X1 U532 ( .A1(G902), .A2(G237), .ZN(n518) );
  NOR2_X1 U533 ( .A1(G953), .A2(G237), .ZN(n569) );
  XNOR2_X1 U534 ( .A(G131), .B(KEYINPUT5), .ZN(n529) );
  XOR2_X1 U535 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n571) );
  XNOR2_X1 U536 ( .A(n398), .B(G128), .ZN(n543) );
  XNOR2_X1 U537 ( .A(n526), .B(n527), .ZN(n493) );
  NOR2_X1 U538 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U539 ( .A(n603), .B(n500), .ZN(n499) );
  NOR2_X1 U540 ( .A1(n602), .A2(n497), .ZN(n496) );
  INV_X1 U541 ( .A(KEYINPUT30), .ZN(n500) );
  XNOR2_X1 U542 ( .A(n648), .B(n482), .ZN(n703) );
  INV_X1 U543 ( .A(KEYINPUT104), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n494), .B(n419), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n561), .B(n472), .ZN(n563) );
  XNOR2_X1 U546 ( .A(n562), .B(n473), .ZN(n472) );
  NOR2_X1 U547 ( .A1(n404), .A2(G475), .ZN(n436) );
  XNOR2_X1 U548 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n501) );
  NAND2_X1 U549 ( .A1(n625), .A2(n682), .ZN(n502) );
  XNOR2_X1 U550 ( .A(n638), .B(KEYINPUT35), .ZN(n639) );
  XNOR2_X1 U551 ( .A(n458), .B(KEYINPUT99), .ZN(n457) );
  AND2_X1 U552 ( .A1(n708), .A2(n460), .ZN(n459) );
  XNOR2_X1 U553 ( .A(n491), .B(n417), .ZN(n490) );
  INV_X1 U554 ( .A(KEYINPUT53), .ZN(n506) );
  XOR2_X1 U555 ( .A(n738), .B(n416), .Z(n404) );
  AND2_X1 U556 ( .A1(n592), .A2(G210), .ZN(n405) );
  INV_X1 U557 ( .A(G953), .ZN(n753) );
  XNOR2_X1 U558 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n406) );
  AND2_X1 U559 ( .A1(n569), .A2(G210), .ZN(n407) );
  AND2_X1 U560 ( .A1(G224), .A2(n753), .ZN(n408) );
  XNOR2_X1 U561 ( .A(n660), .B(KEYINPUT6), .ZN(n626) );
  AND2_X1 U562 ( .A1(n647), .A2(n505), .ZN(n409) );
  AND2_X1 U563 ( .A1(n666), .A2(n515), .ZN(n410) );
  AND2_X1 U564 ( .A1(n706), .A2(n648), .ZN(n412) );
  NAND2_X1 U565 ( .A1(n514), .A2(n727), .ZN(n413) );
  AND2_X1 U566 ( .A1(n466), .A2(n753), .ZN(n414) );
  XOR2_X1 U567 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n415) );
  XNOR2_X1 U568 ( .A(KEYINPUT59), .B(KEYINPUT93), .ZN(n416) );
  XNOR2_X1 U569 ( .A(n403), .B(n730), .ZN(n417) );
  XOR2_X1 U570 ( .A(n517), .B(KEYINPUT65), .Z(n418) );
  XOR2_X1 U571 ( .A(n667), .B(KEYINPUT62), .Z(n419) );
  NOR2_X1 U572 ( .A1(G952), .A2(n753), .ZN(n745) );
  INV_X1 U573 ( .A(n745), .ZN(n439) );
  XOR2_X1 U574 ( .A(n668), .B(KEYINPUT63), .Z(n421) );
  XOR2_X1 U575 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n422) );
  INV_X1 U576 ( .A(KEYINPUT118), .ZN(n727) );
  XNOR2_X2 U577 ( .A(n465), .B(n423), .ZN(n754) );
  XNOR2_X2 U578 ( .A(n582), .B(n424), .ZN(n423) );
  XNOR2_X2 U579 ( .A(n425), .B(n471), .ZN(n424) );
  XNOR2_X2 U580 ( .A(KEYINPUT73), .B(G122), .ZN(n425) );
  XNOR2_X2 U581 ( .A(n426), .B(G107), .ZN(n582) );
  XNOR2_X2 U582 ( .A(G104), .B(G110), .ZN(n426) );
  XNOR2_X2 U583 ( .A(n427), .B(n533), .ZN(n465) );
  XNOR2_X2 U584 ( .A(n428), .B(n485), .ZN(n427) );
  XNOR2_X2 U585 ( .A(G119), .B(KEYINPUT3), .ZN(n428) );
  NAND2_X1 U586 ( .A1(n429), .A2(KEYINPUT44), .ZN(n641) );
  XNOR2_X1 U587 ( .A(n397), .B(G122), .ZN(n773) );
  XOR2_X1 U588 ( .A(KEYINPUT13), .B(G475), .Z(n430) );
  XNOR2_X1 U589 ( .A(KEYINPUT117), .B(n726), .ZN(n431) );
  BUF_X1 U590 ( .A(n750), .Z(n432) );
  XNOR2_X1 U591 ( .A(n443), .B(n464), .ZN(n463) );
  NAND2_X1 U592 ( .A1(n656), .A2(n645), .ZN(n443) );
  INV_X1 U593 ( .A(n644), .ZN(n656) );
  NAND2_X1 U594 ( .A1(n490), .A2(n439), .ZN(n489) );
  XNOR2_X1 U595 ( .A(n652), .B(n441), .ZN(n469) );
  NOR2_X1 U596 ( .A1(n644), .A2(n693), .ZN(n634) );
  XNOR2_X2 U597 ( .A(n433), .B(n406), .ZN(n631) );
  NOR2_X1 U598 ( .A1(n597), .A2(n433), .ZN(n598) );
  NOR2_X2 U599 ( .A1(n438), .A2(n434), .ZN(n467) );
  NAND2_X1 U600 ( .A1(n437), .A2(n435), .ZN(n434) );
  NOR2_X1 U601 ( .A1(n436), .A2(n745), .ZN(n435) );
  XNOR2_X1 U602 ( .A(n509), .B(KEYINPUT83), .ZN(n508) );
  XNOR2_X1 U603 ( .A(n440), .B(n421), .ZN(G57) );
  NAND2_X1 U604 ( .A1(n444), .A2(n414), .ZN(n507) );
  NAND2_X1 U605 ( .A1(n449), .A2(n618), .ZN(n448) );
  INV_X1 U606 ( .A(n694), .ZN(n451) );
  NOR2_X1 U607 ( .A1(n697), .A2(n452), .ZN(n698) );
  NAND2_X1 U608 ( .A1(n456), .A2(n454), .ZN(n453) );
  INV_X1 U609 ( .A(n663), .ZN(n455) );
  NAND2_X1 U610 ( .A1(n659), .A2(n459), .ZN(n458) );
  INV_X1 U611 ( .A(n602), .ZN(n460) );
  NOR2_X2 U612 ( .A1(n631), .A2(n630), .ZN(n461) );
  NAND2_X1 U613 ( .A1(n654), .A2(n412), .ZN(n675) );
  AND2_X1 U614 ( .A1(n463), .A2(n646), .ZN(n654) );
  NAND2_X1 U615 ( .A1(n463), .A2(n409), .ZN(n462) );
  XNOR2_X1 U616 ( .A(n465), .B(n531), .ZN(n504) );
  XNOR2_X1 U617 ( .A(n623), .B(KEYINPUT41), .ZN(n722) );
  XNOR2_X1 U618 ( .A(n467), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U619 ( .A1(n558), .A2(G217), .ZN(n559) );
  XNOR2_X1 U620 ( .A(n548), .B(n547), .ZN(n558) );
  NAND2_X1 U621 ( .A1(n707), .A2(n487), .ZN(n488) );
  NAND2_X1 U622 ( .A1(n511), .A2(n510), .ZN(n509) );
  XNOR2_X1 U623 ( .A(n586), .B(n476), .ZN(n590) );
  XNOR2_X1 U624 ( .A(n587), .B(n408), .ZN(n476) );
  INV_X1 U625 ( .A(n626), .ZN(n486) );
  NAND2_X1 U626 ( .A1(n707), .A2(n708), .ZN(n657) );
  XNOR2_X1 U627 ( .A(n489), .B(n422), .ZN(G51) );
  AND2_X1 U628 ( .A1(n495), .A2(n540), .ZN(n492) );
  XNOR2_X1 U629 ( .A(n762), .B(KEYINPUT75), .ZN(n495) );
  INV_X1 U630 ( .A(n703), .ZN(n505) );
  XNOR2_X1 U631 ( .A(n507), .B(n506), .ZN(G75) );
  INV_X1 U632 ( .A(KEYINPUT2), .ZN(n510) );
  NAND2_X1 U633 ( .A1(n750), .A2(n512), .ZN(n511) );
  INV_X1 U634 ( .A(n762), .ZN(n512) );
  BUF_X1 U635 ( .A(n656), .Z(n659) );
  XOR2_X1 U636 ( .A(KEYINPUT117), .B(n726), .Z(n514) );
  XOR2_X1 U637 ( .A(KEYINPUT82), .B(n665), .Z(n515) );
  INV_X1 U638 ( .A(KEYINPUT91), .ZN(n649) );
  INV_X1 U639 ( .A(KEYINPUT0), .ZN(n632) );
  XNOR2_X1 U640 ( .A(n575), .B(n523), .ZN(n525) );
  XNOR2_X1 U641 ( .A(n530), .B(n407), .ZN(n531) );
  XNOR2_X1 U642 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U643 ( .A1(n666), .A2(n690), .ZN(n762) );
  INV_X1 U644 ( .A(KEYINPUT110), .ZN(n668) );
  NAND2_X1 U645 ( .A1(KEYINPUT2), .A2(n540), .ZN(n517) );
  XOR2_X1 U646 ( .A(KEYINPUT74), .B(n518), .Z(n592) );
  BUF_X1 U647 ( .A(n582), .Z(n527) );
  XOR2_X2 U648 ( .A(KEYINPUT4), .B(KEYINPUT64), .Z(n587) );
  NAND2_X1 U649 ( .A1(G143), .A2(n519), .ZN(n522) );
  NAND2_X1 U650 ( .A1(n520), .A2(G128), .ZN(n521) );
  AND2_X1 U651 ( .A1(G227), .A2(n753), .ZN(n523) );
  NOR2_X1 U652 ( .A1(n732), .A2(G902), .ZN(n528) );
  XNOR2_X1 U653 ( .A(n529), .B(KEYINPUT100), .ZN(n530) );
  NAND2_X1 U654 ( .A1(G234), .A2(G237), .ZN(n534) );
  XNOR2_X1 U655 ( .A(n534), .B(KEYINPUT14), .ZN(n535) );
  NAND2_X1 U656 ( .A1(n535), .A2(G952), .ZN(n720) );
  NOR2_X1 U657 ( .A1(G953), .A2(n720), .ZN(n629) );
  NAND2_X1 U658 ( .A1(G902), .A2(n535), .ZN(n536) );
  XOR2_X1 U659 ( .A(KEYINPUT96), .B(n536), .Z(n537) );
  NAND2_X1 U660 ( .A1(G953), .A2(n537), .ZN(n627) );
  XOR2_X1 U661 ( .A(KEYINPUT105), .B(n627), .Z(n538) );
  NOR2_X1 U662 ( .A1(G900), .A2(n538), .ZN(n539) );
  NAND2_X1 U663 ( .A1(n552), .A2(G221), .ZN(n541) );
  XOR2_X1 U664 ( .A(KEYINPUT10), .B(n588), .Z(n574) );
  XNOR2_X1 U665 ( .A(n542), .B(KEYINPUT24), .ZN(n546) );
  XOR2_X1 U666 ( .A(KEYINPUT23), .B(G140), .Z(n544) );
  XNOR2_X1 U667 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U668 ( .A(n546), .B(n545), .Z(n550) );
  XOR2_X1 U669 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n548) );
  NAND2_X1 U670 ( .A1(G234), .A2(n753), .ZN(n547) );
  NAND2_X1 U671 ( .A1(G221), .A2(n558), .ZN(n549) );
  XNOR2_X1 U672 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U673 ( .A(n574), .B(n551), .ZN(n743) );
  NOR2_X1 U674 ( .A1(G902), .A2(n743), .ZN(n555) );
  XOR2_X1 U675 ( .A(KEYINPUT98), .B(KEYINPUT78), .Z(n554) );
  NAND2_X1 U676 ( .A1(n552), .A2(G217), .ZN(n553) );
  NAND2_X1 U677 ( .A1(n556), .A2(n648), .ZN(n609) );
  INV_X1 U678 ( .A(n557), .ZN(n564) );
  XNOR2_X1 U679 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U680 ( .A(n564), .B(n563), .Z(n740) );
  NOR2_X1 U681 ( .A1(G902), .A2(n740), .ZN(n566) );
  XNOR2_X1 U682 ( .A(KEYINPUT102), .B(G478), .ZN(n565) );
  XNOR2_X1 U683 ( .A(n566), .B(n565), .ZN(n622) );
  XNOR2_X1 U684 ( .A(n568), .B(n567), .ZN(n573) );
  NAND2_X1 U685 ( .A1(n569), .A2(G214), .ZN(n570) );
  XNOR2_X1 U686 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U687 ( .A(n573), .B(n572), .ZN(n576) );
  XNOR2_X1 U688 ( .A(n575), .B(n574), .ZN(n760) );
  XNOR2_X1 U689 ( .A(n576), .B(n760), .ZN(n738) );
  NOR2_X1 U690 ( .A1(G902), .A2(n738), .ZN(n577) );
  XNOR2_X1 U691 ( .A(n621), .B(KEYINPUT101), .ZN(n601) );
  NOR2_X1 U692 ( .A1(n609), .A2(n600), .ZN(n578) );
  NAND2_X1 U693 ( .A1(n486), .A2(n578), .ZN(n597) );
  NOR2_X1 U694 ( .A1(n707), .A2(n597), .ZN(n579) );
  NAND2_X1 U695 ( .A1(n694), .A2(n579), .ZN(n580) );
  XNOR2_X1 U696 ( .A(n580), .B(KEYINPUT43), .ZN(n581) );
  XNOR2_X1 U697 ( .A(KEYINPUT106), .B(n581), .ZN(n594) );
  XOR2_X1 U698 ( .A(KEYINPUT18), .B(KEYINPUT95), .Z(n585) );
  XNOR2_X1 U699 ( .A(KEYINPUT79), .B(KEYINPUT17), .ZN(n584) );
  XNOR2_X1 U700 ( .A(n585), .B(n584), .ZN(n586) );
  INV_X1 U701 ( .A(n588), .ZN(n589) );
  XNOR2_X1 U702 ( .A(n590), .B(n589), .ZN(n591) );
  NAND2_X1 U703 ( .A1(n731), .A2(n664), .ZN(n593) );
  XNOR2_X2 U704 ( .A(n593), .B(n405), .ZN(n596) );
  BUF_X1 U705 ( .A(n596), .Z(n619) );
  INV_X1 U706 ( .A(n619), .ZN(n605) );
  NAND2_X1 U707 ( .A1(n594), .A2(n605), .ZN(n595) );
  XNOR2_X1 U708 ( .A(n595), .B(KEYINPUT107), .ZN(n771) );
  XOR2_X1 U709 ( .A(KEYINPUT36), .B(n598), .Z(n599) );
  NOR2_X1 U710 ( .A1(n646), .A2(n599), .ZN(n687) );
  NAND2_X1 U711 ( .A1(KEYINPUT47), .A2(n697), .ZN(n607) );
  NAND2_X1 U712 ( .A1(n660), .A2(n694), .ZN(n603) );
  OR2_X1 U713 ( .A1(n621), .A2(n622), .ZN(n636) );
  NOR2_X1 U714 ( .A1(n605), .A2(n636), .ZN(n606) );
  NAND2_X1 U715 ( .A1(n411), .A2(n606), .ZN(n678) );
  NAND2_X1 U716 ( .A1(n607), .A2(n678), .ZN(n608) );
  XOR2_X1 U717 ( .A(KEYINPUT84), .B(n608), .Z(n614) );
  INV_X1 U718 ( .A(n660), .ZN(n706) );
  XOR2_X1 U719 ( .A(KEYINPUT28), .B(n610), .Z(n611) );
  INV_X1 U720 ( .A(n631), .ZN(n612) );
  NAND2_X1 U721 ( .A1(KEYINPUT47), .A2(n616), .ZN(n613) );
  NAND2_X1 U722 ( .A1(n614), .A2(n613), .ZN(n615) );
  INV_X1 U723 ( .A(n616), .ZN(n679) );
  NOR2_X1 U724 ( .A1(KEYINPUT47), .A2(n697), .ZN(n617) );
  NAND2_X1 U725 ( .A1(n679), .A2(n617), .ZN(n618) );
  NAND2_X1 U726 ( .A1(n622), .A2(n621), .ZN(n696) );
  NOR2_X1 U727 ( .A1(n771), .A2(n624), .ZN(n666) );
  NAND2_X1 U728 ( .A1(n684), .A2(n625), .ZN(n690) );
  NOR2_X1 U729 ( .A1(n648), .A2(n642), .ZN(n708) );
  NOR2_X1 U730 ( .A1(n627), .A2(G898), .ZN(n628) );
  NOR2_X1 U731 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U732 ( .A(KEYINPUT88), .B(KEYINPUT80), .Z(n638) );
  XNOR2_X1 U733 ( .A(n641), .B(KEYINPUT90), .ZN(n651) );
  OR2_X1 U734 ( .A1(n696), .A2(n642), .ZN(n643) );
  NOR2_X1 U735 ( .A1(n646), .A2(n486), .ZN(n647) );
  NAND2_X1 U736 ( .A1(n400), .A2(KEYINPUT44), .ZN(n650) );
  NAND2_X1 U737 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U738 ( .A1(n401), .A2(n703), .ZN(n655) );
  NOR2_X1 U739 ( .A1(n486), .A2(n655), .ZN(n669) );
  NOR2_X1 U740 ( .A1(n706), .A2(n657), .ZN(n713) );
  NAND2_X1 U741 ( .A1(n659), .A2(n713), .ZN(n658) );
  XNOR2_X1 U742 ( .A(KEYINPUT31), .B(n658), .ZN(n685) );
  NOR2_X1 U743 ( .A1(n685), .A2(n671), .ZN(n661) );
  NOR2_X1 U744 ( .A1(n697), .A2(n661), .ZN(n662) );
  NOR2_X1 U745 ( .A1(n669), .A2(n662), .ZN(n663) );
  NAND2_X1 U746 ( .A1(KEYINPUT2), .A2(n690), .ZN(n665) );
  XOR2_X1 U747 ( .A(G101), .B(n669), .Z(G3) );
  NAND2_X1 U748 ( .A1(n671), .A2(n682), .ZN(n670) );
  XNOR2_X1 U749 ( .A(n670), .B(G104), .ZN(G6) );
  XOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n673) );
  NAND2_X1 U751 ( .A1(n671), .A2(n684), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U753 ( .A(G107), .B(n674), .ZN(G9) );
  XNOR2_X1 U754 ( .A(n675), .B(n398), .ZN(G12) );
  XOR2_X1 U755 ( .A(G128), .B(KEYINPUT29), .Z(n677) );
  NAND2_X1 U756 ( .A1(n684), .A2(n679), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n677), .B(n676), .ZN(G30) );
  XNOR2_X1 U758 ( .A(G143), .B(n678), .ZN(G45) );
  XOR2_X1 U759 ( .A(G146), .B(KEYINPUT111), .Z(n681) );
  NAND2_X1 U760 ( .A1(n679), .A2(n682), .ZN(n680) );
  XNOR2_X1 U761 ( .A(n681), .B(n680), .ZN(G48) );
  NAND2_X1 U762 ( .A1(n685), .A2(n682), .ZN(n683) );
  XNOR2_X1 U763 ( .A(n683), .B(G113), .ZN(G15) );
  NAND2_X1 U764 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U765 ( .A(n686), .B(G116), .ZN(G18) );
  XNOR2_X1 U766 ( .A(n687), .B(KEYINPUT112), .ZN(n688) );
  XNOR2_X1 U767 ( .A(n688), .B(KEYINPUT37), .ZN(n689) );
  XNOR2_X1 U768 ( .A(G125), .B(n689), .ZN(G27) );
  XNOR2_X1 U769 ( .A(G134), .B(n690), .ZN(G36) );
  NOR2_X1 U770 ( .A1(n696), .A2(n695), .ZN(n699) );
  NOR2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U772 ( .A1(n723), .A2(n700), .ZN(n701) );
  XNOR2_X1 U773 ( .A(n701), .B(KEYINPUT115), .ZN(n717) );
  NOR2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U775 ( .A(n704), .B(KEYINPUT49), .ZN(n705) );
  NAND2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n711) );
  NOR2_X1 U777 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U778 ( .A(n709), .B(KEYINPUT50), .ZN(n710) );
  NOR2_X1 U779 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U782 ( .A(KEYINPUT52), .B(n718), .Z(n719) );
  NOR2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U784 ( .A(KEYINPUT116), .B(n721), .ZN(n725) );
  NOR2_X1 U785 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U786 ( .A(KEYINPUT85), .B(KEYINPUT55), .Z(n729) );
  XNOR2_X1 U787 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n728) );
  XNOR2_X1 U788 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U789 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n734) );
  XNOR2_X1 U790 ( .A(n732), .B(KEYINPUT57), .ZN(n733) );
  XNOR2_X1 U791 ( .A(n734), .B(n733), .ZN(n736) );
  XNOR2_X1 U792 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U793 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U794 ( .A1(n745), .A2(n741), .ZN(G63) );
  XNOR2_X1 U795 ( .A(n743), .B(n742), .ZN(n744) );
  XOR2_X1 U796 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n747) );
  NAND2_X1 U797 ( .A1(G224), .A2(G953), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U799 ( .A(KEYINPUT122), .B(n748), .ZN(n749) );
  NAND2_X1 U800 ( .A1(n749), .A2(G898), .ZN(n752) );
  NAND2_X1 U801 ( .A1(n432), .A2(n753), .ZN(n751) );
  NAND2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n758) );
  OR2_X1 U803 ( .A1(n753), .A2(G898), .ZN(n756) );
  BUF_X1 U804 ( .A(n754), .Z(n755) );
  NAND2_X1 U805 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U806 ( .A(n758), .B(n757), .Z(G69) );
  XNOR2_X1 U807 ( .A(KEYINPUT124), .B(n759), .ZN(n761) );
  XNOR2_X1 U808 ( .A(n761), .B(n760), .ZN(n764) );
  XNOR2_X1 U809 ( .A(n764), .B(n762), .ZN(n763) );
  NOR2_X1 U810 ( .A1(G953), .A2(n763), .ZN(n769) );
  XNOR2_X1 U811 ( .A(n764), .B(KEYINPUT125), .ZN(n765) );
  XNOR2_X1 U812 ( .A(G227), .B(n765), .ZN(n767) );
  NAND2_X1 U813 ( .A1(G900), .A2(G953), .ZN(n766) );
  NOR2_X1 U814 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U815 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U816 ( .A(KEYINPUT126), .B(n770), .ZN(G72) );
  XOR2_X1 U817 ( .A(G140), .B(n771), .Z(G42) );
  XNOR2_X1 U818 ( .A(G131), .B(n772), .ZN(G33) );
  XNOR2_X1 U819 ( .A(n773), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U820 ( .A(n402), .B(G119), .ZN(G21) );
  XNOR2_X1 U821 ( .A(G137), .B(n775), .ZN(G39) );
endmodule

