//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G107), .C2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  AND2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n206), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT0), .Z(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n231), .A2(new_n204), .A3(new_n232), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n227), .A2(new_n230), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G264), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT16), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(KEYINPUT73), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT73), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n254), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n252), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT7), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(G20), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n207), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n223), .A2(new_n207), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G58), .A2(G68), .ZN(new_n264));
  OAI21_X1  g0064(.A(G20), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT72), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(new_n267), .A3(G159), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n266), .B2(G159), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n250), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n232), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n254), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n256), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n261), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G68), .ZN(new_n279));
  INV_X1    g0079(.A(new_n271), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(KEYINPUT16), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n272), .A2(new_n274), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT64), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OR3_X1    g0085(.A1(new_n284), .A2(new_n223), .A3(KEYINPUT8), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n204), .A2(G1), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G13), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n274), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(KEYINPUT65), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n288), .A2(KEYINPUT65), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n290), .B1(new_n295), .B2(new_n287), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n282), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G41), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(G1), .A3(G13), .ZN(new_n299));
  INV_X1    g0099(.A(G223), .ZN(new_n300));
  INV_X1    g0100(.A(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n219), .A2(G1698), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n256), .A2(new_n302), .A3(new_n275), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G87), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n307));
  INV_X1    g0107(.A(G274), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n299), .A2(G232), .A3(new_n307), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NOR4_X1   g0114(.A1(new_n306), .A2(new_n314), .A3(new_n310), .A4(new_n309), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n297), .B(KEYINPUT18), .C1(new_n313), .C2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT18), .ZN(new_n317));
  INV_X1    g0117(.A(G13), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n318), .A2(new_n204), .A3(G1), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n285), .B2(new_n286), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n274), .ZN(new_n321));
  INV_X1    g0121(.A(new_n294), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(new_n292), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n285), .A2(new_n286), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n271), .B1(new_n278), .B2(G68), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n291), .B1(new_n326), .B2(KEYINPUT16), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n325), .B1(new_n327), .B2(new_n272), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n313), .A2(new_n315), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n317), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n304), .A2(new_n305), .ZN(new_n333));
  INV_X1    g0133(.A(new_n299), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n309), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n310), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  NOR4_X1   g0138(.A1(new_n306), .A2(new_n338), .A3(new_n310), .A4(new_n309), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n337), .A2(new_n339), .A3(new_n325), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n340), .A2(new_n282), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n340), .B2(new_n282), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n340), .A2(new_n282), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n344), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n340), .A2(new_n282), .A3(new_n341), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT75), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n331), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT76), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n224), .A2(G1698), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G226), .B2(G1698), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n356), .A2(new_n276), .B1(new_n251), .B2(new_n212), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n309), .B1(new_n357), .B2(new_n334), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n299), .A2(new_n307), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G238), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT13), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n358), .A2(new_n364), .A3(new_n361), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(G179), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT70), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n366), .B(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G169), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n370), .A2(KEYINPUT14), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(KEYINPUT14), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n319), .A2(new_n207), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT12), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n207), .B2(new_n323), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n266), .A2(G50), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n204), .A2(G33), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n378), .B1(new_n204), .B2(G68), .C1(new_n220), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n274), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT11), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT11), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n383), .A3(new_n274), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n376), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT71), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n373), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n385), .B1(new_n369), .B2(new_n338), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n332), .B1(new_n363), .B2(new_n365), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G20), .A2(G77), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT15), .B(G87), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n204), .A2(new_n251), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n392), .B1(new_n393), .B2(new_n379), .C1(new_n394), .C2(new_n283), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n274), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n319), .A2(new_n220), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n397), .B(KEYINPUT66), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n396), .B(new_n398), .C1(new_n220), .C2(new_n323), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G238), .A2(G1698), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n260), .B(new_n400), .C1(new_n224), .C2(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n334), .C1(G107), .C2(new_n260), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n309), .B1(new_n360), .B2(G244), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n399), .B1(G190), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n332), .B2(new_n405), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n354), .A2(new_n388), .A3(new_n391), .A4(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n204), .B1(new_n264), .B2(new_n218), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(G150), .B2(new_n266), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n287), .B2(new_n379), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(new_n274), .B1(new_n218), .B2(new_n319), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n218), .B2(new_n323), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT9), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n301), .A2(G222), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n260), .B(new_n415), .C1(new_n300), .C2(new_n301), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n334), .C1(G77), .C2(new_n260), .ZN(new_n417));
  INV_X1    g0217(.A(new_n309), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n219), .C2(new_n359), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n338), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(G200), .B2(new_n419), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT68), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT10), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n422), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n419), .A2(new_n312), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n413), .B(new_n428), .C1(G179), .C2(new_n419), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT67), .B1(new_n405), .B2(G169), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(G179), .B2(new_n404), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n405), .A2(KEYINPUT67), .A3(new_n314), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n399), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n427), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n353), .A2(KEYINPUT76), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n408), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT21), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n301), .A2(G257), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G264), .A2(G1698), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n256), .A2(new_n275), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n334), .C1(G303), .C2(new_n260), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT5), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G41), .ZN(new_n444));
  INV_X1    g0244(.A(G41), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT5), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n444), .A2(new_n446), .A3(new_n203), .A4(G45), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(G270), .A3(new_n299), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n203), .A2(G45), .A3(G274), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n445), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT78), .B1(new_n445), .B2(KEYINPUT5), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n450), .B(new_n444), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n442), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G169), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n203), .A2(G33), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n291), .A2(new_n289), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(G20), .B1(G33), .B2(G283), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT77), .B(G97), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G33), .ZN(new_n462));
  AOI221_X4 g0262(.A(KEYINPUT81), .B1(new_n458), .B2(G20), .C1(new_n273), .C2(new_n232), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT81), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n458), .A2(G20), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n274), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n462), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT20), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n462), .B(KEYINPUT20), .C1(new_n463), .C2(new_n466), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n289), .A2(G116), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI211_X1 g0273(.A(new_n438), .B(new_n455), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n459), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n274), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT81), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n274), .A2(new_n464), .A3(new_n465), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT20), .B1(new_n479), .B2(new_n462), .ZN(new_n480));
  INV_X1    g0280(.A(new_n470), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n473), .B(new_n475), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n455), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT21), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT82), .ZN(new_n486));
  INV_X1    g0286(.A(new_n454), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n482), .A2(G179), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(G190), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n454), .A2(G200), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n471), .A3(new_n473), .A4(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n485), .A2(new_n486), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  AOI211_X1 g0292(.A(new_n472), .B(new_n459), .C1(new_n469), .C2(new_n470), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n438), .B1(new_n493), .B2(new_n455), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n482), .A2(KEYINPUT21), .A3(new_n483), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n494), .A2(new_n488), .A3(new_n495), .A4(new_n491), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT82), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n208), .A2(new_n301), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n221), .A2(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n256), .A2(new_n499), .A3(new_n275), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G116), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n299), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n449), .B(KEYINPUT80), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n203), .A2(G45), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n299), .A2(G250), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(new_n332), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(G190), .B2(new_n508), .ZN(new_n510));
  NAND3_X1  g0310(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n204), .ZN(new_n512));
  XOR2_X1   g0312(.A(KEYINPUT77), .B(G97), .Z(new_n513));
  INV_X1    g0313(.A(G107), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n210), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n260), .A2(new_n204), .A3(G68), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n461), .A2(new_n379), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n516), .B(new_n517), .C1(KEYINPUT19), .C2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n274), .B1(new_n319), .B2(new_n393), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n321), .A2(G87), .A3(new_n456), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n510), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n457), .A2(new_n393), .ZN(new_n524));
  OR3_X1    g0324(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n520), .A2(new_n524), .B1(new_n312), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n508), .A2(new_n314), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n256), .A2(new_n275), .A3(G244), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G283), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n531), .A2(G1698), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n534), .A2(new_n256), .A3(new_n275), .A4(G244), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n256), .A2(new_n275), .A3(G250), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n301), .B1(new_n537), .B2(KEYINPUT4), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n334), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n447), .A2(G257), .A3(new_n299), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n453), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n539), .A2(new_n338), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(G200), .B1(new_n539), .B2(new_n542), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n319), .A2(new_n212), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n457), .B2(new_n212), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n514), .B1(new_n258), .B2(new_n261), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n513), .A2(KEYINPUT6), .A3(new_n514), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n212), .A2(new_n514), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n204), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n394), .A2(new_n220), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n549), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n548), .B1(new_n557), .B2(new_n291), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n545), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n550), .A2(new_n554), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G20), .ZN(new_n561));
  INV_X1    g0361(.A(new_n556), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n258), .A2(new_n261), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n514), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n547), .B1(new_n564), .B2(new_n274), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n539), .A2(new_n314), .A3(new_n542), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n530), .A2(new_n531), .B1(G33), .B2(G283), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n531), .B1(new_n260), .B2(G250), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n567), .B(new_n535), .C1(new_n301), .C2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n541), .B1(new_n569), .B2(new_n334), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n566), .B1(new_n570), .B2(G169), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT79), .B1(new_n559), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n539), .A2(new_n542), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n312), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n558), .A2(new_n566), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT79), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n576), .B(new_n577), .C1(new_n558), .C2(new_n545), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n529), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT25), .B1(new_n289), .B2(G107), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT25), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n319), .A2(new_n581), .A3(new_n514), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n582), .C1(new_n457), .C2(new_n514), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT84), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n321), .A2(G107), .A3(new_n456), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT84), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n580), .A4(new_n582), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n203), .B(G45), .C1(new_n443), .C2(G41), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n445), .A2(KEYINPUT5), .ZN(new_n590));
  OAI211_X1 g0390(.A(G264), .B(new_n299), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT85), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT85), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n447), .A2(new_n593), .A3(G264), .A4(new_n299), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n211), .A2(new_n301), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n213), .A2(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n256), .A2(new_n596), .A3(new_n275), .A4(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(G294), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n251), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n334), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n595), .A2(new_n453), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G200), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT24), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n256), .A2(new_n275), .A3(new_n204), .A4(G87), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT22), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n260), .A2(KEYINPUT22), .A3(new_n204), .A4(G87), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT23), .ZN(new_n610));
  OAI211_X1 g0410(.A(G20), .B(new_n514), .C1(new_n610), .C2(KEYINPUT83), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT83), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(KEYINPUT23), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(KEYINPUT83), .B(new_n610), .C1(new_n204), .C2(G107), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n614), .A2(new_n616), .B1(new_n458), .B2(new_n379), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n604), .B1(new_n609), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n379), .A2(new_n458), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n610), .A2(KEYINPUT83), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n612), .A2(KEYINPUT23), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(G20), .A4(new_n514), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n619), .B1(new_n622), .B2(new_n615), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n623), .A2(KEYINPUT24), .A3(new_n607), .A4(new_n608), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n618), .A2(new_n274), .A3(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n592), .A2(new_n594), .B1(new_n600), .B2(new_n334), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(G190), .A3(new_n453), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n588), .A2(new_n603), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n625), .A2(new_n588), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n602), .A2(new_n312), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n314), .A3(new_n453), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n629), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n625), .A2(new_n588), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(KEYINPUT86), .A3(new_n632), .A4(new_n631), .ZN(new_n636));
  AOI211_X1 g0436(.A(KEYINPUT87), .B(new_n628), .C1(new_n634), .C2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT87), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n636), .ZN(new_n639));
  INV_X1    g0439(.A(new_n628), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n498), .B(new_n579), .C1(new_n637), .C2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n437), .A2(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n433), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n391), .A2(new_n644), .B1(new_n373), .B2(new_n387), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n347), .B1(new_n342), .B2(new_n346), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n333), .A2(new_n334), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(G190), .A3(new_n418), .A4(new_n336), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n296), .B(new_n648), .C1(new_n332), .C2(new_n311), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n272), .B2(new_n327), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n351), .B(KEYINPUT75), .C1(new_n650), .C2(new_n345), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n331), .B1(new_n645), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT89), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(KEYINPUT89), .B(new_n331), .C1(new_n645), .C2(new_n653), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n427), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n429), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n494), .A2(new_n488), .A3(new_n495), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n635), .A2(new_n632), .A3(new_n631), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT88), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT88), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n635), .A2(new_n664), .A3(new_n632), .A4(new_n631), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n522), .A2(new_n510), .B1(new_n526), .B2(new_n527), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n559), .A2(new_n572), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n666), .A2(new_n640), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n528), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n529), .B2(new_n576), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n667), .A2(KEYINPUT26), .A3(new_n572), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n436), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n660), .A2(new_n677), .ZN(G369));
  INV_X1    g0478(.A(KEYINPUT91), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n318), .A2(G20), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n203), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n630), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n639), .A2(new_n640), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT87), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n639), .A2(new_n638), .A3(new_n640), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n662), .A2(new_n687), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n679), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n641), .A2(new_n637), .B1(new_n630), .B2(new_n687), .ZN(new_n695));
  INV_X1    g0495(.A(new_n693), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(KEYINPUT91), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n661), .A2(new_n493), .A3(new_n687), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n498), .B1(new_n493), .B2(new_n687), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n663), .A2(new_n665), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n686), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n661), .A2(new_n686), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n698), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n228), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G1), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n461), .A2(new_n210), .A3(new_n514), .A4(new_n458), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(new_n231), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n686), .B1(new_n669), .B2(new_n675), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT29), .B1(new_n722), .B2(KEYINPUT94), .ZN(new_n723));
  INV_X1    g0523(.A(G330), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n487), .A2(G179), .A3(new_n508), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n626), .A2(new_n539), .A3(new_n542), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n442), .A2(G179), .A3(new_n448), .A4(new_n453), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n525), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n570), .A3(KEYINPUT30), .A4(new_n626), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n508), .A2(G179), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n574), .A3(new_n454), .A4(new_n602), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n686), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT93), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT92), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT93), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n735), .A2(new_n742), .A3(new_n736), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n738), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n739), .A2(new_n740), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n742), .B1(new_n735), .B2(new_n736), .ZN(new_n746));
  AOI211_X1 g0546(.A(KEYINPUT93), .B(KEYINPUT31), .C1(new_n734), .C2(new_n686), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n690), .A2(new_n691), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(new_n498), .A3(new_n579), .A4(new_n687), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n724), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT95), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n639), .A2(new_n661), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n639), .B2(new_n661), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n668), .A2(new_n640), .A3(new_n667), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n675), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT94), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n759), .A2(new_n687), .B1(new_n722), .B2(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n723), .B(new_n752), .C1(new_n761), .C2(KEYINPUT29), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n720), .B1(new_n762), .B2(G1), .ZN(G364));
  AOI21_X1  g0563(.A(new_n717), .B1(G45), .B2(new_n680), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n705), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n232), .B1(G20), .B2(new_n312), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n714), .A2(new_n260), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n231), .A2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(G45), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n773), .B(new_n774), .C1(new_n245), .C2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n228), .A2(G355), .A3(new_n260), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n776), .B(new_n777), .C1(G116), .C2(new_n228), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n765), .B(new_n770), .C1(new_n772), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n314), .A2(new_n332), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n204), .A2(new_n338), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n204), .A2(G190), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n332), .A2(G179), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n782), .A2(new_n218), .B1(new_n785), .B2(new_n514), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n204), .B1(new_n787), .B2(G190), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G97), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n314), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n781), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n276), .B1(new_n797), .B2(G58), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n781), .A2(new_n784), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n783), .A2(new_n795), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G87), .A2(new_n800), .B1(new_n802), .B2(G77), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n791), .A2(new_n794), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n780), .A2(new_n783), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n786), .B(new_n804), .C1(G68), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G283), .ZN(new_n810));
  INV_X1    g0610(.A(G329), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n785), .A2(new_n810), .B1(new_n788), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n782), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(G326), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n793), .A2(G294), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n260), .B1(new_n800), .B2(G303), .ZN(new_n816));
  INV_X1    g0616(.A(G317), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(KEYINPUT33), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n806), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n814), .A2(new_n815), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n809), .B(new_n821), .C1(G322), .C2(new_n797), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n771), .B1(new_n807), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n764), .B1(new_n705), .B2(G330), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n705), .A2(G330), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n779), .A2(new_n823), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n644), .A2(new_n687), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n399), .A2(new_n686), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n407), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n433), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n721), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(new_n752), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n765), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n785), .A2(new_n210), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n794), .B1(new_n808), .B2(new_n788), .ZN(new_n839));
  INV_X1    g0639(.A(G303), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n782), .A2(new_n840), .B1(new_n801), .B2(new_n458), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G283), .B2(new_n806), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n842), .A2(KEYINPUT96), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(KEYINPUT96), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n838), .B(new_n839), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n260), .B1(new_n800), .B2(G107), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(new_n599), .C2(new_n796), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT97), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G143), .A2(new_n797), .B1(new_n802), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n850), .B2(new_n782), .C1(new_n851), .C2(new_n805), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n276), .B1(new_n852), .B2(new_n853), .ZN(new_n855));
  INV_X1    g0655(.A(new_n788), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(G132), .ZN(new_n857));
  INV_X1    g0657(.A(new_n785), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G50), .A2(new_n800), .B1(new_n858), .B2(G68), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n855), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n854), .B(new_n860), .C1(G58), .C2(new_n793), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n771), .B1(new_n848), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n771), .A2(new_n766), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n220), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n833), .A2(new_n766), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n862), .A2(new_n764), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n837), .A2(new_n866), .ZN(G384));
  OAI211_X1 g0667(.A(new_n739), .B(new_n737), .C1(new_n642), .C2(new_n686), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n387), .A2(new_n686), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n388), .A2(new_n869), .A3(new_n391), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n389), .A2(new_n390), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n387), .B(new_n686), .C1(new_n373), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n833), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n327), .B1(KEYINPUT16), .B2(new_n326), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n296), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n329), .A2(new_n684), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n875), .B1(new_n879), .B2(new_n349), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n297), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n881), .A2(new_n875), .A3(new_n349), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n684), .B1(new_n652), .B2(new_n331), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n874), .B(new_n883), .C1(new_n884), .C2(new_n877), .ZN(new_n885));
  INV_X1    g0685(.A(new_n684), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n353), .A2(new_n886), .A3(new_n877), .ZN(new_n887));
  INV_X1    g0687(.A(new_n883), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n868), .B(new_n873), .C1(new_n885), .C2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n342), .A2(new_n346), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n328), .B(new_n684), .C1(new_n331), .C2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n875), .B1(new_n881), .B2(new_n349), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n882), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n874), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n868), .A4(new_n873), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n892), .A2(G330), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n868), .A2(G330), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n436), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n892), .A2(new_n868), .A3(new_n900), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n437), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT100), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n723), .B1(new_n761), .B2(KEYINPUT29), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(new_n437), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n659), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n908), .B(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n721), .A2(new_n832), .B1(new_n644), .B2(new_n687), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n877), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n684), .B(new_n915), .C1(new_n652), .C2(new_n331), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n874), .B1(new_n916), .B2(new_n883), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n893), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n870), .A2(new_n872), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n316), .A2(new_n330), .A3(new_n684), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n899), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(KEYINPUT99), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT99), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n918), .B2(KEYINPUT39), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n899), .A2(KEYINPUT39), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n373), .A2(new_n387), .A3(new_n687), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n922), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n912), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n203), .B2(new_n680), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n560), .B(KEYINPUT98), .Z(new_n935));
  INV_X1    g0735(.A(KEYINPUT35), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n204), .B(new_n232), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n937), .B(G116), .C1(new_n936), .C2(new_n935), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  OAI21_X1  g0739(.A(G77), .B1(new_n223), .B2(new_n207), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n940), .A2(new_n231), .B1(G50), .B2(new_n207), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n318), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(new_n939), .A3(new_n942), .ZN(G367));
  OAI21_X1  g0743(.A(new_n668), .B1(new_n565), .B2(new_n687), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n572), .A2(new_n686), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n707), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT103), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n711), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n694), .B2(new_n697), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n946), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT42), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n576), .B1(new_n944), .B2(new_n639), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n687), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n522), .A2(new_n687), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT101), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n671), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT102), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(new_n529), .C2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n961), .B2(new_n960), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n957), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n966), .B1(new_n957), .B2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n949), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n970), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n947), .A2(new_n948), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n968), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n715), .B(KEYINPUT41), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT44), .B1(new_n712), .B2(new_n946), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  INV_X1    g0778(.A(new_n946), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n951), .C2(new_n710), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT45), .B1(new_n712), .B2(new_n946), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n951), .A2(new_n982), .A3(new_n710), .A4(new_n979), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n977), .B(new_n980), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n707), .ZN(new_n985));
  INV_X1    g0785(.A(new_n697), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT91), .B1(new_n695), .B2(new_n696), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n711), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n710), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n988), .A2(new_n989), .A3(new_n946), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n982), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n712), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n993), .A2(new_n708), .A3(new_n977), .A4(new_n980), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n698), .A2(new_n711), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n951), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(KEYINPUT104), .A3(new_n706), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n706), .B(KEYINPUT104), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n985), .A2(new_n994), .A3(new_n762), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n976), .B1(new_n1000), .B2(new_n762), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n680), .A2(G45), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(G1), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT105), .Z(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n971), .B(new_n974), .C1(new_n1001), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n773), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n237), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n772), .B1(new_n228), .B2(new_n393), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n788), .A2(new_n850), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n813), .A2(G143), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n793), .A2(G68), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(new_n851), .C2(new_n796), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT107), .Z(new_n1014));
  NAND2_X1  g0814(.A1(new_n806), .A2(G159), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n858), .A2(G77), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(KEYINPUT108), .A3(new_n260), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT108), .B1(new_n1016), .B2(new_n260), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G50), .B2(new_n802), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1010), .B(new_n1020), .C1(G58), .C2(new_n800), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n858), .A2(new_n513), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n800), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT46), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n799), .B2(new_n458), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(new_n599), .C2(new_n805), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT106), .Z(new_n1027));
  NAND2_X1  g0827(.A1(new_n813), .A2(G311), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n796), .A2(new_n840), .B1(new_n801), .B2(new_n810), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G317), .B2(new_n856), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n276), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G107), .B2(new_n793), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1021), .B1(new_n1022), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n771), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n764), .B1(new_n1008), .B2(new_n1009), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT109), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n769), .B2(new_n964), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1006), .A2(new_n1038), .ZN(G387));
  OR2_X1    g0839(.A1(new_n999), .A2(new_n762), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n999), .A2(new_n762), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n715), .A3(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G322), .A2(new_n813), .B1(new_n806), .B2(G311), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n840), .B2(new_n801), .C1(new_n817), .C2(new_n796), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT48), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n810), .B2(new_n792), .C1(new_n599), .C2(new_n799), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT49), .Z(new_n1047));
  AOI21_X1  g0847(.A(new_n260), .B1(new_n856), .B2(G326), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n458), .B2(new_n785), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT111), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n799), .A2(new_n220), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G68), .B2(new_n802), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n212), .B2(new_n785), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n287), .A2(new_n805), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n260), .B1(new_n788), .B2(new_n851), .C1(new_n218), .C2(new_n796), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n782), .A2(new_n789), .B1(new_n792), .B2(new_n393), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n771), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n764), .C1(new_n698), .C2(new_n769), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n718), .A2(new_n228), .A3(new_n260), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n718), .B(KEYINPUT110), .Z(new_n1062));
  NOR2_X1   g0862(.A1(new_n207), .A2(new_n220), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT50), .B1(new_n283), .B2(G50), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n775), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n283), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1066));
  NOR4_X1   g0866(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n773), .B1(new_n241), .B2(new_n775), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1061), .B1(G107), .B2(new_n228), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1060), .B1(new_n772), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n999), .B2(new_n1005), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1042), .A2(new_n1071), .ZN(G393));
  INV_X1    g0872(.A(KEYINPUT112), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n985), .A2(new_n1073), .A3(new_n994), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n984), .A2(KEYINPUT112), .A3(new_n707), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n1041), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n715), .A3(new_n1000), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(KEYINPUT114), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT114), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1076), .A2(new_n1079), .A3(new_n715), .A4(new_n1000), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1005), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n782), .A2(new_n851), .B1(new_n796), .B2(new_n789), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT51), .Z(new_n1085));
  OAI22_X1  g0885(.A1(new_n799), .A2(new_n207), .B1(new_n801), .B2(new_n283), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1085), .A2(new_n838), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n806), .A2(G50), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n856), .A2(G143), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n276), .B1(new_n793), .B2(G77), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n782), .A2(new_n817), .B1(new_n796), .B2(new_n808), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT52), .Z(new_n1093));
  AOI22_X1  g0893(.A1(G107), .A2(new_n858), .B1(new_n856), .B2(G322), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1094), .B(new_n276), .C1(new_n810), .C2(new_n799), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT113), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1093), .B(new_n1096), .C1(G303), .C2(new_n806), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n599), .B2(new_n801), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n792), .A2(new_n458), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1091), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n771), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n979), .A2(new_n768), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n772), .B1(new_n228), .B2(new_n461), .C1(new_n1007), .C2(new_n248), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n764), .A4(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1081), .A2(new_n1083), .A3(new_n1104), .ZN(G390));
  NOR3_X1   g0905(.A1(new_n899), .A2(new_n926), .A3(KEYINPUT39), .ZN(new_n1106));
  OAI21_X1  g0906(.A(KEYINPUT39), .B1(new_n885), .B2(new_n889), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT99), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n923), .A2(new_n924), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n766), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n287), .A2(new_n863), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n260), .B1(new_n785), .B2(new_n218), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT116), .Z(new_n1114));
  AOI22_X1  g0914(.A1(G128), .A2(new_n813), .B1(new_n797), .B2(G132), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT54), .B(G143), .Z(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1114), .B(new_n1115), .C1(new_n801), .C2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n805), .A2(new_n850), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n800), .A2(G150), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT53), .ZN(new_n1121));
  INV_X1    g0921(.A(G125), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1122), .A2(new_n788), .B1(new_n792), .B2(new_n789), .ZN(new_n1123));
  NOR4_X1   g0923(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n801), .A2(new_n461), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G87), .A2(new_n800), .B1(new_n858), .B2(G68), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n813), .A2(G283), .B1(new_n856), .B2(G294), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n806), .A2(G107), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n260), .B1(new_n793), .B2(G77), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1125), .B(new_n1130), .C1(G116), .C2(new_n797), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n771), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1111), .A2(new_n764), .A3(new_n1112), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n919), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n930), .B1(new_n913), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n925), .B(new_n1135), .C1(new_n927), .C2(new_n928), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n687), .B(new_n832), .C1(new_n757), .C2(new_n676), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1134), .B1(new_n1137), .B2(new_n829), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n899), .A2(new_n930), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n752), .A2(new_n834), .A3(new_n919), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1136), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1110), .B2(new_n1135), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n903), .A2(new_n873), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1133), .B1(new_n1146), .B2(new_n1004), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1134), .B1(new_n902), .B2(new_n833), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1137), .A2(new_n829), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1148), .A2(new_n1149), .A3(new_n1142), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n642), .A2(new_n686), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n744), .A2(new_n748), .ZN(new_n1152));
  OAI211_X1 g0952(.A(G330), .B(new_n834), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1134), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT115), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT115), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1153), .A2(new_n1156), .A3(new_n1134), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1157), .A3(new_n1145), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1150), .B1(new_n1158), .B2(new_n914), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n660), .B(new_n904), .C1(new_n909), .C2(new_n437), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1136), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1145), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n716), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(new_n914), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1150), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1160), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1146), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1147), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(G378));
  NAND2_X1  g0973(.A1(new_n427), .A2(new_n429), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1175), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n427), .A2(new_n429), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n413), .A2(new_n886), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1176), .A2(new_n413), .A3(new_n886), .A4(new_n1178), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n766), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G41), .B1(new_n813), .B2(G116), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n223), .B2(new_n785), .C1(new_n514), .C2(new_n796), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1052), .B(new_n1186), .C1(G283), .C2(new_n856), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n805), .A2(new_n212), .B1(new_n801), .B2(new_n393), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT117), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n276), .A3(new_n1012), .A4(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT58), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n445), .B1(new_n254), .B2(new_n251), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1190), .A2(new_n1191), .B1(new_n218), .B2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT118), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G128), .A2(new_n797), .B1(new_n802), .B2(G137), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n800), .A2(new_n1116), .B1(new_n793), .B2(G150), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n813), .A2(G125), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G132), .B2(new_n806), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT59), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G33), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(G41), .B1(new_n856), .B2(G124), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n789), .C2(new_n785), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1190), .A2(new_n1191), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n771), .B1(new_n1194), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n863), .A2(new_n218), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1184), .A2(new_n764), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1183), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n901), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT119), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1183), .A2(new_n892), .A3(G330), .A4(new_n900), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n932), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n920), .B(new_n921), .C1(new_n1110), .C2(new_n930), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1216), .A2(new_n1212), .A3(new_n1213), .A4(new_n1211), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1209), .B1(new_n1218), .B2(new_n1005), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1160), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1216), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n932), .A2(new_n1213), .A3(new_n1211), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(KEYINPUT57), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n715), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1169), .B1(new_n1146), .B2(new_n1159), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT57), .B1(new_n1226), .B2(new_n1218), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1219), .B1(new_n1225), .B2(new_n1227), .ZN(G375));
  AOI22_X1  g1028(.A1(G137), .A2(new_n797), .B1(new_n858), .B2(G58), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n813), .A2(G132), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(new_n851), .C2(new_n801), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G159), .B2(new_n800), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n260), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G128), .B2(new_n856), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n218), .B2(new_n792), .C1(new_n805), .C2(new_n1117), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1016), .B1(new_n514), .B2(new_n801), .C1(new_n458), .C2(new_n805), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G283), .B2(new_n797), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n799), .A2(new_n212), .B1(new_n792), .B2(new_n393), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n260), .B(new_n1238), .C1(G294), .C2(new_n813), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1237), .B(new_n1239), .C1(new_n840), .C2(new_n788), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT121), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1035), .B1(new_n1235), .B2(new_n1241), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n765), .B(new_n1242), .C1(new_n207), .C2(new_n863), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT122), .Z(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n766), .B2(new_n1134), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT120), .B1(new_n1159), .B2(new_n1004), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT120), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1154), .A2(KEYINPUT115), .B1(new_n903), .B2(new_n873), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n913), .B1(new_n1248), .B2(new_n1157), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1247), .B(new_n1005), .C1(new_n1249), .C2(new_n1150), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1245), .B1(new_n1246), .B2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1166), .A2(new_n1160), .A3(new_n1167), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1170), .A2(new_n975), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1251), .A2(new_n1253), .ZN(G381));
  INV_X1    g1054(.A(KEYINPUT123), .ZN(new_n1255));
  INV_X1    g1055(.A(G387), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1104), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1258), .A3(new_n1083), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1259), .A2(G384), .A3(G381), .ZN(new_n1260));
  OR2_X1    g1060(.A1(G375), .A2(G378), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1042), .A2(new_n827), .A3(new_n1071), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1255), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1259), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(G381), .A2(G384), .ZN(new_n1266));
  AND4_X1   g1066(.A1(new_n1255), .A2(new_n1265), .A3(new_n1266), .A4(new_n1263), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1264), .A2(new_n1267), .ZN(G407));
  OR2_X1    g1068(.A1(new_n1261), .A2(G343), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G213), .B(new_n1269), .C1(new_n1264), .C2(new_n1267), .ZN(G409));
  NAND2_X1  g1070(.A1(G375), .A2(G378), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n685), .A2(G213), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1252), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1159), .A2(KEYINPUT60), .A3(new_n1160), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1170), .A3(new_n1275), .A4(new_n715), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1276), .A2(new_n1251), .A3(G384), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G384), .B1(new_n1276), .B2(new_n1251), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1226), .A2(new_n1218), .A3(new_n975), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(KEYINPUT124), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1222), .A2(new_n1005), .A3(new_n1223), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1282), .A2(new_n1208), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1226), .A2(new_n1218), .A3(new_n1284), .A4(new_n975), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1281), .A2(new_n1172), .A3(new_n1283), .A4(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1271), .A2(new_n1272), .A3(new_n1279), .A4(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(G375), .A2(G378), .B1(G213), .B2(new_n685), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1289), .A2(new_n1286), .A3(new_n1279), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1278), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1276), .A2(new_n1251), .A3(G384), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n685), .A2(G213), .A3(G2897), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1295), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1289), .A2(new_n1286), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT61), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G390), .A2(G387), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G393), .A2(G396), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1262), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT126), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1307), .A3(new_n1262), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1303), .A2(new_n1309), .A3(new_n1259), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1308), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n1303), .B2(new_n1259), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1292), .B(new_n1302), .C1(new_n1310), .C2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1289), .A2(new_n1314), .A3(new_n1286), .A4(new_n1279), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT62), .B1(new_n1315), .B2(KEYINPUT127), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1271), .A2(new_n1272), .A3(new_n1286), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1318), .B2(new_n1299), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1314), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1287), .A2(new_n1321), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1316), .A2(new_n1319), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1303), .A2(new_n1259), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1308), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1303), .A2(new_n1259), .A3(new_n1309), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1313), .B1(new_n1323), .B2(new_n1327), .ZN(G405));
  AOI211_X1 g1128(.A(new_n1278), .B(new_n1277), .C1(new_n1261), .C2(new_n1271), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1261), .A2(new_n1271), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1330), .A2(new_n1279), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(new_n1326), .A3(new_n1325), .ZN(new_n1333));
  OAI22_X1  g1133(.A1(new_n1310), .A2(new_n1312), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(G402));
endmodule


