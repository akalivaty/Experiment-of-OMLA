//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(new_n203), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT64), .Z(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n214), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n213), .B(new_n217), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G250), .B(G257), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G264), .B(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n230), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  AND2_X1   g0044(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n245));
  NOR2_X1   g0045(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(new_n232), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT72), .ZN(new_n251));
  AND2_X1   g0051(.A1(new_n248), .A2(G1698), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n252), .A2(G238), .B1(new_n255), .B2(G107), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G1), .A2(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT67), .B(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT68), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n266), .B1(new_n258), .B2(new_n259), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT67), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n272), .A3(new_n263), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n267), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT68), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G244), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n274), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n260), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n261), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G179), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI221_X1 g0084(.A(new_n277), .B1(new_n278), .B2(new_n280), .C1(new_n257), .C2(new_n260), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n289), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n211), .A2(G33), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT15), .B(G87), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n210), .ZN(new_n296));
  INV_X1    g0096(.A(G77), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n274), .A2(G13), .A3(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT70), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n300), .A2(new_n274), .A3(G13), .A4(G20), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n294), .A2(new_n296), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n301), .ZN(new_n304));
  INV_X1    g0104(.A(new_n296), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n211), .A2(G1), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n306), .A2(new_n297), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n284), .A2(new_n287), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n285), .A2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n309), .B(new_n303), .C1(new_n285), .C2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n317));
  INV_X1    g0117(.A(G150), .ZN(new_n318));
  INV_X1    g0118(.A(G33), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n211), .A2(new_n319), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n317), .B1(new_n318), .B2(new_n320), .C1(new_n292), .C2(new_n288), .ZN(new_n321));
  INV_X1    g0121(.A(G50), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n321), .A2(new_n296), .B1(new_n302), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n306), .ZN(new_n324));
  INV_X1    g0124(.A(new_n307), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(G50), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n326), .A3(KEYINPUT9), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT73), .ZN(new_n328));
  INV_X1    g0128(.A(new_n260), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT69), .B(G1698), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n255), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n331), .A2(G222), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n248), .A2(G1698), .ZN(new_n333));
  INV_X1    g0133(.A(G223), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n333), .A2(new_n334), .B1(new_n297), .B2(new_n248), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n329), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n280), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G226), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n277), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G190), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n323), .A2(new_n326), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT9), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n339), .A2(G200), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n328), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT10), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT10), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n328), .A2(new_n347), .A3(new_n341), .A4(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT71), .B1(new_n340), .B2(G169), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(G179), .B2(new_n339), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n340), .A2(KEYINPUT71), .A3(new_n283), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n342), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n248), .A2(G226), .A3(G1698), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G87), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n355), .B(new_n356), .C1(new_n249), .C2(new_n334), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n329), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n337), .A2(G232), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n265), .B1(new_n264), .B2(new_n267), .ZN(new_n361));
  AND4_X1   g0161(.A1(new_n265), .A2(new_n273), .A3(new_n267), .A4(new_n274), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G169), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n268), .A2(new_n276), .B1(G232), .B2(new_n337), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(G179), .A3(new_n358), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n248), .B2(G20), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n202), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT76), .B1(new_n320), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT76), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n290), .A2(new_n375), .A3(G159), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g0177(.A(G58), .B(G68), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n368), .B1(new_n372), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n255), .B2(new_n211), .ZN(new_n382));
  NOR4_X1   g0182(.A1(new_n253), .A2(new_n254), .A3(new_n369), .A4(G20), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n374), .A2(new_n376), .B1(new_n378), .B2(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n386), .A3(new_n296), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n288), .A2(new_n307), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n324), .A2(new_n388), .B1(new_n302), .B2(new_n288), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n367), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT18), .ZN(new_n392));
  INV_X1    g0192(.A(new_n390), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n365), .A2(G190), .A3(new_n358), .ZN(new_n394));
  OAI21_X1  g0194(.A(G200), .B1(new_n359), .B2(new_n363), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n393), .A2(KEYINPUT17), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n387), .A3(new_n389), .A4(new_n394), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n367), .A2(new_n400), .A3(new_n390), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n392), .A2(new_n396), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n316), .A2(new_n354), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n304), .A2(G68), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT12), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n306), .A2(new_n202), .A3(new_n307), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n292), .A2(new_n297), .B1(new_n211), .B2(G68), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT74), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n408), .A2(new_n409), .B1(new_n322), .B2(new_n320), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n408), .A2(new_n409), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n296), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT11), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n412), .A2(new_n413), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n407), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT75), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT14), .ZN(new_n419));
  INV_X1    g0219(.A(G238), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n280), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n268), .B2(new_n276), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  OR2_X1    g0223(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n424));
  NAND2_X1  g0224(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(G226), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G232), .A2(G1698), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n255), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G97), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n329), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n422), .A2(new_n423), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n423), .B1(new_n422), .B2(new_n431), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n419), .B(G169), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n361), .A2(new_n362), .B1(new_n420), .B2(new_n280), .ZN(new_n435));
  INV_X1    g0235(.A(new_n431), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n422), .A2(new_n423), .A3(new_n431), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(G179), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n419), .B1(new_n441), .B2(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n418), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(G169), .B1(new_n432), .B2(new_n433), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n445), .A2(KEYINPUT75), .A3(new_n439), .A4(new_n434), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n417), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(G200), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n437), .A2(G190), .A3(new_n438), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n417), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n403), .A2(new_n452), .ZN(new_n453));
  OR3_X1    g0253(.A1(new_n211), .A2(KEYINPUT23), .A3(G107), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G116), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT84), .ZN(new_n457));
  OAI221_X1 g0257(.A(new_n454), .B1(G20), .B2(new_n455), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n456), .A2(new_n457), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT24), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n248), .A2(new_n211), .A3(G87), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT22), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT22), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n248), .A2(new_n464), .A3(new_n211), .A4(G87), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n460), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n461), .B1(new_n460), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n296), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n306), .B1(new_n274), .B2(G33), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G107), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n304), .A2(G107), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT25), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n247), .A2(new_n248), .A3(G250), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT85), .A2(G294), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT85), .A2(G294), .ZN(new_n478));
  OAI21_X1  g0278(.A(G33), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n329), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n262), .A2(KEYINPUT5), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n274), .B(G45), .C1(new_n483), .C2(G41), .ZN(new_n484));
  OAI211_X1 g0284(.A(G264), .B(new_n260), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT86), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n270), .A2(new_n272), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n484), .B1(new_n488), .B2(new_n483), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n267), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT86), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n481), .A2(new_n491), .A3(new_n485), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n487), .A2(G179), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT87), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n481), .A2(new_n490), .A3(new_n485), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G169), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n493), .B2(new_n494), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n474), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n474), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n502));
  INV_X1    g0302(.A(G200), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n497), .A2(G190), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G244), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT79), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT79), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n248), .A2(new_n511), .A3(G244), .A4(G1698), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n455), .B1(new_n249), .B2(new_n420), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT80), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n455), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n331), .B2(G238), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT80), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n510), .A2(new_n512), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n515), .A2(new_n329), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n274), .A2(new_n266), .A3(G45), .ZN(new_n522));
  INV_X1    g0322(.A(G250), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n263), .B2(G1), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n260), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(G169), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n525), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n517), .A2(new_n519), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n260), .B1(new_n528), .B2(KEYINPUT80), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n527), .B1(new_n529), .B2(new_n520), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n526), .B1(new_n283), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n293), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n470), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n211), .B1(new_n429), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G87), .B2(new_n206), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n211), .B(G68), .C1(new_n253), .C2(new_n254), .ZN(new_n537));
  INV_X1    g0337(.A(G97), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n534), .B1(new_n292), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n296), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n302), .A2(new_n293), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n541), .A2(KEYINPUT81), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT81), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n533), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT82), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT82), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n547), .B(new_n533), .C1(new_n543), .C2(new_n544), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n521), .A2(new_n525), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G200), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n274), .A2(G33), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n304), .A2(new_n305), .A3(G87), .A4(new_n552), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT83), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n543), .B2(new_n544), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n530), .B2(G190), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n531), .A2(new_n549), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G257), .ZN(new_n558));
  OR2_X1    g0358(.A1(KEYINPUT3), .A2(G33), .ZN(new_n559));
  NAND2_X1  g0359(.A1(KEYINPUT3), .A2(G33), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n247), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n248), .A2(G264), .A3(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n255), .A2(G303), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n329), .ZN(new_n566));
  OAI211_X1 g0366(.A(G270), .B(new_n260), .C1(new_n482), .C2(new_n484), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n490), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  INV_X1    g0369(.A(G116), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n302), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n304), .A2(new_n305), .A3(G116), .A4(new_n552), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n295), .A2(new_n210), .B1(G20), .B2(new_n570), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G283), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n211), .C1(G33), .C2(new_n538), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT20), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n573), .A2(KEYINPUT20), .A3(new_n575), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n571), .B(new_n572), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n569), .B(new_n579), .C1(new_n568), .C2(new_n314), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n568), .A2(G169), .A3(new_n578), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n567), .A2(new_n490), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n561), .A2(new_n247), .B1(new_n255), .B2(G303), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n260), .B1(new_n585), .B2(new_n563), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G179), .A3(new_n578), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n568), .A2(KEYINPUT21), .A3(G169), .A4(new_n578), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n580), .A2(new_n583), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n324), .A2(G97), .A3(new_n552), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(G97), .B2(new_n304), .ZN(new_n593));
  OAI21_X1  g0393(.A(G107), .B1(new_n382), .B2(new_n383), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT6), .ZN(new_n595));
  AND2_X1   g0395(.A1(G97), .A2(G107), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n205), .ZN(new_n597));
  INV_X1    g0397(.A(G107), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(KEYINPUT6), .A3(G97), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT77), .B1(new_n602), .B2(new_n305), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n305), .B1(new_n594), .B2(new_n601), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT77), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n593), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(G257), .B(new_n260), .C1(new_n482), .C2(new_n484), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n490), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT4), .A4(G244), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(new_n574), .C1(new_n523), .C2(new_n333), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n247), .A2(new_n248), .A3(G244), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT4), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT78), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT78), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(new_n617), .A3(new_n614), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n610), .B1(new_n619), .B2(new_n260), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G200), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n252), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n613), .A2(new_n617), .A3(new_n614), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n617), .B1(new_n613), .B2(new_n614), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n611), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n609), .B1(new_n625), .B2(new_n329), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G190), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n607), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n620), .A2(new_n286), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n626), .A2(new_n283), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n304), .A2(G97), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n470), .B2(G97), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n604), .A2(new_n605), .ZN(new_n633));
  AOI211_X1 g0433(.A(KEYINPUT77), .B(new_n305), .C1(new_n594), .C2(new_n601), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n629), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n557), .A2(new_n591), .A3(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n453), .A2(new_n508), .A3(new_n638), .ZN(G372));
  AND2_X1   g0439(.A1(new_n396), .A2(new_n399), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n311), .A2(new_n451), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n447), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n392), .A2(new_n401), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n349), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n353), .ZN(new_n646));
  INV_X1    g0446(.A(new_n453), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n550), .A2(new_n286), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n530), .A2(new_n283), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n541), .A2(new_n542), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT81), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n541), .A2(KEYINPUT81), .A3(new_n542), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n547), .B1(new_n654), .B2(new_n533), .ZN(new_n655));
  INV_X1    g0455(.A(new_n548), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n648), .B(new_n649), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n556), .A2(new_n551), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n659), .B1(new_n661), .B2(new_n636), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n629), .A2(new_n630), .A3(new_n635), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n557), .A2(KEYINPUT26), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n583), .A2(new_n588), .A3(new_n589), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n500), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT88), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND4_X1   g0470(.A1(new_n636), .A2(new_n657), .A3(new_n628), .A4(new_n660), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n500), .A2(KEYINPUT88), .A3(new_n667), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n507), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n647), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n646), .A2(new_n675), .ZN(G369));
  NAND3_X1  g0476(.A1(new_n274), .A2(new_n211), .A3(G13), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT89), .Z(new_n679));
  INV_X1    g0479(.A(G213), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n677), .B2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G343), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n474), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n500), .A2(new_n507), .A3(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n481), .A2(new_n491), .A3(new_n485), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n491), .B1(new_n481), .B2(new_n485), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(KEYINPUT87), .A3(G179), .A4(new_n490), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n495), .A3(new_n498), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n474), .A3(new_n685), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n684), .A2(new_n579), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n590), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n666), .A2(new_n696), .ZN(new_n698));
  OAI21_X1  g0498(.A(G330), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n666), .A2(new_n684), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n500), .A3(new_n507), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n692), .A2(new_n474), .A3(new_n684), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n700), .A2(new_n704), .ZN(G399));
  INV_X1    g0505(.A(new_n215), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n488), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n208), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT90), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT91), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n690), .A2(new_n714), .A3(new_n525), .A4(new_n521), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n568), .A2(new_n283), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT92), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n521), .A2(new_n487), .A3(new_n492), .A4(new_n525), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n626), .A4(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n716), .A3(new_n626), .A4(new_n715), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT92), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n620), .A2(new_n724), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n717), .A2(KEYINPUT94), .A3(new_n720), .A4(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n720), .A2(new_n716), .A3(new_n715), .A4(new_n726), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT94), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT93), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n568), .A2(new_n283), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n732), .B1(new_n530), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n587), .A2(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n550), .A2(KEYINPUT93), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n626), .B1(new_n490), .B2(new_n690), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n725), .A2(new_n731), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n684), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n500), .A2(new_n507), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n671), .A2(new_n743), .A3(new_n591), .A4(new_n684), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n738), .A2(KEYINPUT95), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT95), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n734), .A2(new_n736), .A3(new_n737), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n725), .A2(new_n731), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n750), .B2(new_n685), .ZN(new_n751));
  OAI21_X1  g0551(.A(G330), .B1(new_n745), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n668), .A2(new_n507), .A3(new_n557), .A4(new_n637), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT26), .B1(new_n557), .B2(new_n663), .ZN(new_n754));
  AND4_X1   g0554(.A1(KEYINPUT26), .A2(new_n657), .A3(new_n663), .A4(new_n660), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n753), .B(new_n657), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(KEYINPUT29), .A3(new_n684), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n685), .B1(new_n665), .B2(new_n673), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n758), .B2(KEYINPUT29), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n752), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n713), .B1(new_n760), .B2(G1), .ZN(G364));
  NAND2_X1  g0561(.A1(new_n211), .A2(G13), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n274), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n707), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n697), .A2(new_n698), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(new_n767), .B2(G330), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n767), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT96), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n210), .B1(G20), .B2(new_n286), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n314), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n211), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n538), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G190), .A2(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G20), .A3(new_n283), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G159), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n774), .B1(KEYINPUT32), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n211), .A2(new_n283), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G190), .A3(new_n503), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n255), .B1(new_n782), .B2(G58), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n780), .A2(new_n775), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n779), .B(new_n783), .C1(new_n297), .C2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n211), .A2(new_n503), .A3(G179), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n780), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G190), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G87), .A2(new_n788), .B1(new_n790), .B2(G68), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n789), .A2(new_n314), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n791), .B1(KEYINPUT32), .B2(new_n778), .C1(new_n322), .C2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n786), .A2(new_n314), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT99), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT99), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n785), .B(new_n794), .C1(G107), .C2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n782), .A2(G322), .B1(G329), .B2(new_n777), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n801), .B(new_n255), .C1(new_n802), .C2(new_n784), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G303), .A2(new_n788), .B1(new_n792), .B2(G326), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n477), .A2(new_n478), .ZN(new_n805));
  INV_X1    g0605(.A(new_n790), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT33), .B(G317), .Z(new_n807));
  OAI221_X1 g0607(.A(new_n804), .B1(new_n805), .B2(new_n773), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n803), .B(new_n808), .C1(G283), .C2(new_n799), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n771), .B1(new_n800), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G13), .A2(G33), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n771), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT98), .Z(new_n815));
  INV_X1    g0615(.A(new_n243), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n706), .A2(new_n248), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(new_n263), .B2(new_n209), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n816), .A2(G45), .B1(new_n819), .B2(KEYINPUT97), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(KEYINPUT97), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n706), .A2(new_n255), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n822), .A2(G355), .B1(new_n570), .B2(new_n706), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n810), .B(new_n766), .C1(new_n815), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT100), .ZN(new_n826));
  INV_X1    g0626(.A(new_n813), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n767), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n770), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  OR2_X1    g0631(.A1(new_n771), .A2(new_n811), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n766), .B1(G77), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT101), .ZN(new_n834));
  INV_X1    g0634(.A(G283), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n806), .A2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n774), .B(new_n836), .C1(G303), .C2(new_n792), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n255), .B1(new_n787), .B2(new_n598), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n799), .A2(G87), .ZN(new_n840));
  INV_X1    g0640(.A(G294), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n781), .A2(new_n841), .B1(new_n784), .B2(new_n570), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G311), .B2(new_n777), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n837), .A2(new_n839), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n784), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n782), .A2(G143), .B1(new_n845), .B2(G159), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n806), .B2(new_n318), .C1(new_n847), .C2(new_n793), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT34), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n799), .A2(G68), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n255), .B1(new_n777), .B2(G132), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n201), .B2(new_n773), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G50), .B2(new_n788), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n851), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n844), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n834), .B1(new_n857), .B2(new_n771), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n284), .A2(new_n287), .A3(new_n310), .A4(new_n684), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n685), .A2(new_n310), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n313), .B2(new_n315), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n860), .B1(new_n862), .B2(new_n311), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n858), .B1(new_n863), .B2(new_n812), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n758), .B(new_n863), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n766), .B1(new_n865), .B2(new_n752), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n752), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(G384));
  OR2_X1    g0669(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n600), .A2(KEYINPUT35), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(G116), .A3(new_n212), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT36), .Z(new_n873));
  OAI211_X1 g0673(.A(new_n209), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n322), .A2(G68), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n274), .B(G13), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n310), .B1(new_n282), .B2(G190), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n878), .A2(new_n312), .B1(new_n310), .B2(new_n685), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n284), .A2(new_n287), .A3(new_n310), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n859), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n417), .A2(new_n684), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n452), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n447), .B2(new_n451), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT40), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n390), .A2(new_n683), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n643), .B2(new_n640), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n391), .A2(new_n397), .A3(new_n889), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n891), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n888), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n387), .A2(KEYINPUT103), .A3(new_n389), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT103), .B1(new_n387), .B2(new_n389), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n683), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n402), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n397), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n390), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n895), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n901), .B1(new_n904), .B2(new_n367), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n892), .B1(new_n905), .B2(new_n898), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n391), .A2(new_n892), .A3(new_n397), .A4(new_n889), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(KEYINPUT38), .B(new_n900), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n887), .B1(new_n894), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n750), .A2(new_n741), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n744), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n886), .B(new_n910), .C1(new_n912), .C2(new_n751), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT105), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n727), .A2(new_n730), .B1(new_n746), .B2(new_n748), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n684), .B1(new_n916), .B2(new_n725), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n911), .B(new_n744), .C1(KEYINPUT31), .C2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n918), .A2(KEYINPUT105), .A3(new_n886), .A4(new_n910), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n909), .A2(KEYINPUT104), .ZN(new_n921));
  INV_X1    g0721(.A(new_n900), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n367), .B1(new_n896), .B2(new_n897), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n898), .A2(new_n923), .A3(new_n397), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n908), .B1(new_n924), .B2(KEYINPUT37), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n888), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n907), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT104), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT38), .A4(new_n900), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n921), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(new_n886), .C1(new_n912), .C2(new_n751), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n887), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n750), .A2(new_n685), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n740), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n638), .A2(new_n508), .A3(new_n685), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n750), .B2(new_n741), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n453), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n920), .A2(new_n933), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(new_n920), .B2(new_n933), .ZN(new_n940));
  INV_X1    g0740(.A(G330), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT106), .Z(new_n943));
  OAI21_X1  g0743(.A(new_n657), .B1(new_n754), .B2(new_n755), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n557), .A2(new_n507), .A3(new_n637), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n669), .B(new_n666), .C1(new_n692), .C2(new_n474), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT88), .B1(new_n500), .B2(new_n667), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n684), .B(new_n863), .C1(new_n944), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n859), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n443), .A2(new_n446), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n416), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n883), .B1(new_n952), .B2(new_n450), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n447), .A2(new_n451), .A3(new_n882), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n950), .A2(new_n956), .A3(new_n931), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n643), .A2(new_n683), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n894), .A2(new_n909), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT39), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(KEYINPUT39), .B2(new_n931), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n447), .A2(new_n684), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n957), .B(new_n958), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n647), .B(new_n757), .C1(KEYINPUT29), .C2(new_n758), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n646), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n963), .B(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n943), .A2(new_n967), .B1(new_n274), .B2(new_n763), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n943), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n877), .B1(new_n968), .B2(new_n969), .ZN(G367));
  NOR2_X1   g0770(.A1(new_n230), .A2(new_n818), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n814), .B1(new_n215), .B2(new_n293), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n766), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n799), .A2(G77), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n784), .A2(new_n322), .B1(new_n776), .B2(new_n847), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n255), .B(new_n975), .C1(G150), .C2(new_n782), .ZN(new_n976));
  INV_X1    g0776(.A(new_n773), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G68), .A2(new_n977), .B1(new_n790), .B2(G159), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G58), .A2(new_n788), .B1(new_n792), .B2(G143), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n974), .A2(new_n976), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n799), .A2(G97), .ZN(new_n981));
  INV_X1    g0781(.A(new_n805), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G107), .A2(new_n977), .B1(new_n790), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(new_n802), .C2(new_n793), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n788), .A2(KEYINPUT46), .A3(G116), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n248), .B1(new_n782), .B2(G303), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n845), .A2(G283), .B1(new_n777), .B2(G317), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT46), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n787), .B2(new_n570), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n985), .A2(new_n986), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n980), .B1(new_n984), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT47), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n973), .B1(new_n992), .B2(new_n771), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n684), .B1(new_n654), .B2(new_n554), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT107), .B1(new_n658), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n661), .B2(new_n994), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n658), .A2(KEYINPUT107), .A3(new_n994), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n993), .B1(new_n998), .B2(new_n827), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT111), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n694), .B2(new_n701), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n699), .A2(KEYINPUT112), .B1(new_n743), .B2(new_n701), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n701), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n687), .A2(KEYINPUT111), .A3(new_n693), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n699), .A2(KEYINPUT112), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1006), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1008), .A2(new_n1001), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(new_n752), .A3(new_n759), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT113), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n752), .A3(KEYINPUT113), .A4(new_n759), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n628), .B(new_n636), .C1(new_n607), .C2(new_n684), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n663), .A2(new_n685), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n703), .B2(new_n702), .ZN(new_n1018));
  XOR2_X1   g0818(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1017), .A2(new_n702), .A3(new_n703), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT45), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n700), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT45), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1023), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n700), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1027), .A2(new_n1028), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1013), .A2(new_n1014), .A3(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(KEYINPUT114), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT114), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1033), .B1(new_n1035), .B2(new_n1014), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n760), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n707), .B(KEYINPUT41), .Z(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n765), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT42), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1017), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n702), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1017), .A2(KEYINPUT42), .A3(new_n743), .A4(new_n701), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n636), .B1(new_n1015), .B2(new_n500), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1043), .A2(new_n1044), .B1(new_n684), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT108), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n1048), .A3(KEYINPUT43), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT43), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1046), .B2(KEYINPUT108), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1047), .A2(new_n998), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n998), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT109), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1028), .A2(new_n1042), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n998), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT109), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n1061), .A3(new_n1053), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1057), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1058), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n999), .B1(new_n1040), .B2(new_n1066), .ZN(G387));
  NAND2_X1  g0867(.A1(new_n695), .A2(new_n813), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n822), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1069), .A2(new_n709), .B1(G107), .B2(new_n215), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n235), .A2(new_n263), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n709), .ZN(new_n1072));
  AOI211_X1 g0872(.A(G45), .B(new_n1072), .C1(G68), .C2(G77), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n288), .A2(G50), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT50), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n818), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1070), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n766), .B1(new_n1077), .B2(new_n815), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n781), .A2(new_n322), .B1(new_n784), .B2(new_n202), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n255), .B(new_n1079), .C1(G150), .C2(new_n777), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n532), .A2(new_n977), .B1(new_n792), .B2(G159), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G77), .A2(new_n788), .B1(new_n790), .B2(new_n289), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n981), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n248), .B1(new_n777), .B2(G326), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n782), .A2(G317), .B1(new_n845), .B2(G303), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n792), .A2(G322), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n802), .C2(new_n806), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n788), .A2(new_n982), .B1(new_n977), .B2(G283), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT49), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1084), .B1(new_n570), .B2(new_n798), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1083), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1078), .B1(new_n1096), .B2(new_n771), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1010), .A2(new_n765), .B1(new_n1068), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1011), .A2(new_n707), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n760), .B2(new_n1010), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1098), .B1(new_n1101), .B2(new_n1102), .ZN(G393));
  NAND2_X1  g0903(.A1(new_n1030), .A2(new_n765), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n240), .A2(new_n818), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n814), .B1(new_n538), .B2(new_n215), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n766), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n799), .A2(G107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n255), .B1(new_n784), .B2(new_n841), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G322), .B2(new_n777), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n977), .A2(G116), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G283), .A2(new_n788), .B1(new_n790), .B2(G303), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G317), .A2(new_n792), .B1(new_n782), .B2(G311), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT52), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G150), .A2(new_n792), .B1(new_n782), .B2(G159), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n840), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n788), .A2(G68), .B1(new_n977), .B2(G77), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n777), .A2(G143), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n255), .B1(new_n845), .B2(new_n289), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n790), .A2(G50), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1113), .A2(new_n1115), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1107), .B1(new_n1126), .B2(new_n771), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1017), .B2(new_n827), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1104), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1031), .A2(KEYINPUT114), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1035), .A2(new_n1033), .A3(new_n1014), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n708), .B1(new_n1034), .B2(new_n1011), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(G390));
  NOR2_X1   g0935(.A1(new_n881), .A2(new_n941), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n918), .A2(new_n956), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1136), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n936), .B1(new_n739), .B2(new_n741), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n935), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1137), .B1(new_n1140), .B2(new_n956), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n950), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n862), .A2(new_n311), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n756), .A2(new_n684), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n859), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n918), .A2(new_n1136), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n955), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1140), .A2(new_n956), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1142), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n647), .A2(new_n918), .A3(G330), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT117), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n938), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n965), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n685), .B1(new_n665), .B2(new_n753), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n860), .B1(new_n1157), .B2(new_n1143), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n959), .B(new_n962), .C1(new_n1158), .C2(new_n955), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n962), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n950), .B2(new_n956), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n931), .A2(KEYINPUT39), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(KEYINPUT39), .B2(new_n959), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1159), .B(new_n1148), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n959), .A2(new_n962), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1145), .B2(new_n956), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n860), .B1(new_n758), .B2(new_n863), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n962), .B1(new_n1167), .B2(new_n955), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n1168), .B2(new_n961), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1164), .B1(new_n1169), .B2(new_n1137), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1156), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1159), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1172), .A2(new_n918), .A3(new_n956), .A4(new_n1136), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1173), .A2(new_n1150), .A3(new_n1155), .A4(new_n1164), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1171), .A2(new_n1174), .A3(new_n707), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n766), .B1(new_n289), .B2(new_n832), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n781), .A2(new_n570), .B1(new_n784), .B2(new_n538), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n248), .B(new_n1177), .C1(G294), .C2(new_n777), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n788), .A2(G87), .B1(new_n977), .B2(G77), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G107), .A2(new_n790), .B1(new_n792), .B2(G283), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n852), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT120), .Z(new_n1182));
  OAI21_X1  g0982(.A(new_n248), .B1(new_n798), .B2(new_n322), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT119), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n782), .A2(G132), .B1(G125), .B2(new_n777), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n373), .B2(new_n773), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G128), .B2(new_n792), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n788), .A2(G150), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT53), .Z(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n790), .A2(G137), .B1(new_n845), .B2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT118), .Z(new_n1195));
  NAND4_X1  g0995(.A1(new_n1186), .A2(new_n1189), .A3(new_n1191), .A4(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1182), .B1(new_n1185), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1176), .B1(new_n1197), .B2(new_n771), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1163), .B2(new_n812), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1170), .B2(new_n764), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT121), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1173), .A2(new_n765), .A3(new_n1164), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT121), .B1(new_n1203), .B2(new_n1199), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1175), .B1(new_n1202), .B2(new_n1204), .ZN(G378));
  NAND2_X1  g1005(.A1(new_n683), .A2(new_n342), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n354), .B(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1207), .B(new_n1208), .Z(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n811), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n766), .B1(G50), .B2(new_n832), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n322), .B1(G33), .B2(G41), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n255), .B2(new_n262), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n798), .A2(new_n201), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n255), .B(new_n262), .C1(new_n787), .C2(new_n297), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT122), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G68), .A2(new_n977), .B1(new_n792), .B2(G116), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n538), .B2(new_n806), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n782), .A2(G107), .B1(G283), .B2(new_n777), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n293), .B2(new_n784), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1214), .A2(new_n1216), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1213), .B1(new_n1221), .B2(KEYINPUT58), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G33), .B(G41), .C1(new_n777), .C2(G124), .ZN(new_n1223));
  INV_X1    g1023(.A(G128), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n781), .A2(new_n1224), .B1(new_n784), .B2(new_n847), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n788), .A2(new_n1193), .B1(new_n790), .B2(G132), .ZN(new_n1226));
  INV_X1    g1026(.A(G125), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n793), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1225), .B(new_n1228), .C1(G150), .C2(new_n977), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT59), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1223), .B1(new_n373), .B2(new_n798), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1229), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1222), .B1(KEYINPUT58), .B2(new_n1221), .C1(new_n1231), .C2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1211), .B1(new_n1234), .B2(new_n771), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1210), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n941), .B1(new_n932), .B2(new_n887), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1209), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n920), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n920), .B2(new_n1237), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n963), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n863), .B1(new_n953), .B2(new_n954), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n935), .B2(new_n937), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT105), .B1(new_n1243), .B2(new_n910), .ZN(new_n1244));
  AND4_X1   g1044(.A1(KEYINPUT105), .A2(new_n918), .A3(new_n886), .A4(new_n910), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1237), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1209), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n963), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n920), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1241), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1236), .B1(new_n1251), .B2(new_n765), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1141), .A2(new_n950), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1155), .B1(new_n1170), .B2(new_n1253), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1239), .A2(new_n1240), .A3(new_n963), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1248), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1256));
  OAI211_X1 g1056(.A(KEYINPUT57), .B(new_n1254), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n707), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT57), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1252), .B1(new_n1258), .B2(new_n1259), .ZN(G375));
  NAND2_X1  g1060(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n646), .A3(new_n964), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1253), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1038), .B(KEYINPUT123), .Z(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1156), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n955), .A2(new_n811), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n766), .B1(G68), .B2(new_n832), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n781), .A2(new_n835), .B1(new_n784), .B2(new_n598), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n248), .B(new_n1268), .C1(G303), .C2(new_n777), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n532), .A2(new_n977), .B1(new_n790), .B2(G116), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G97), .A2(new_n788), .B1(new_n792), .B2(G294), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n974), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G50), .A2(new_n977), .B1(new_n790), .B2(new_n1193), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(G159), .A2(new_n788), .B1(new_n792), .B2(G132), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n255), .B1(new_n777), .B2(G128), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n782), .A2(G137), .B1(new_n845), .B2(G150), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1272), .B1(new_n1214), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1267), .B1(new_n1278), .B2(new_n771), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1150), .A2(new_n765), .B1(new_n1266), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1265), .A2(new_n1280), .ZN(G381));
  NOR4_X1   g1081(.A1(G381), .A2(G396), .A3(G393), .A4(G384), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1282), .A2(new_n1134), .ZN(new_n1283));
  INV_X1    g1083(.A(G375), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n999), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n760), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n764), .B1(new_n1287), .B2(new_n1038), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1285), .B1(new_n1288), .B2(new_n1065), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1175), .A2(new_n1203), .A3(new_n1199), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1283), .A2(new_n1284), .A3(new_n1289), .A4(new_n1290), .ZN(G407));
  NOR2_X1   g1091(.A1(new_n680), .A2(G343), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1284), .A2(new_n1290), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(G407), .A2(G213), .A3(new_n1293), .ZN(G409));
  XNOR2_X1  g1094(.A(G393), .B(new_n830), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1289), .A2(G390), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1285), .B(new_n1134), .C1(new_n1288), .C2(new_n1065), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(new_n1134), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1289), .A2(G390), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1295), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G378), .B(new_n1252), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1251), .A2(new_n1254), .A3(new_n1264), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1252), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1290), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1292), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1262), .A2(new_n1253), .A3(KEYINPUT60), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n707), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1156), .A2(KEYINPUT60), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1263), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G384), .B1(new_n1317), .B2(new_n1280), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(G384), .B(new_n1280), .C1(new_n1322), .C2(new_n1313), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1311), .B1(new_n1318), .B2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1280), .B1(new_n1322), .B2(new_n1313), .ZN(new_n1326));
  INV_X1    g1126(.A(G384), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(KEYINPUT125), .A3(new_n1323), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1325), .A2(KEYINPUT62), .A3(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1310), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1308), .A2(KEYINPUT124), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1328), .A2(KEYINPUT125), .A3(new_n1323), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT125), .B1(new_n1328), .B2(new_n1323), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT124), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1304), .A2(new_n1307), .A3(new_n1336), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1332), .A2(new_n1309), .A3(new_n1335), .A4(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1331), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1318), .A2(new_n1324), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1292), .A2(G2897), .ZN(new_n1342));
  OR2_X1    g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1325), .A2(new_n1329), .A3(new_n1342), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1310), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT61), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1303), .B1(new_n1340), .B2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1299), .A2(new_n1302), .A3(new_n1346), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(KEYINPUT126), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT126), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1299), .A2(new_n1302), .A3(new_n1351), .A4(new_n1346), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1350), .A2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT63), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1338), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1332), .A2(new_n1309), .A3(new_n1337), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1356), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1335), .A2(KEYINPUT63), .A3(new_n1309), .A4(new_n1308), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1353), .A2(new_n1355), .A3(new_n1357), .A4(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1348), .A2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(G375), .A2(new_n1290), .ZN(new_n1361));
  OR2_X1    g1161(.A1(new_n1361), .A2(KEYINPUT127), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1335), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1361), .A2(KEYINPUT127), .A3(new_n1304), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1362), .A2(new_n1363), .A3(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1341), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1367), .B1(new_n1362), .B2(new_n1364), .ZN(new_n1368));
  OAI211_X1 g1168(.A(new_n1302), .B(new_n1299), .C1(new_n1366), .C2(new_n1368), .ZN(new_n1369));
  AND2_X1   g1169(.A1(new_n1362), .A2(new_n1364), .ZN(new_n1370));
  OAI211_X1 g1170(.A(new_n1303), .B(new_n1365), .C1(new_n1370), .C2(new_n1367), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1369), .A2(new_n1371), .ZN(G402));
endmodule


