//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(KEYINPUT28), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n202), .B(new_n203), .C1(new_n205), .C2(KEYINPUT28), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT26), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n207), .A2(new_n208), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(G183gat), .A3(G190gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT23), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(KEYINPUT24), .ZN(new_n224));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n222), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n216), .B1(KEYINPUT23), .B2(new_n213), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n229), .B(new_n222), .C1(new_n224), .C2(new_n225), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n231), .B(new_n230), .C1(new_n226), .C2(new_n227), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n234), .B1(new_n233), .B2(new_n235), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n220), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G134gat), .ZN(new_n239));
  INV_X1    g038(.A(G120gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G113gat), .ZN(new_n241));
  INV_X1    g040(.A(G113gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G120gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT1), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G127gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n247), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n239), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n245), .ZN(new_n250));
  OAI21_X1  g049(.A(G127gat), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(G134gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n255), .B(new_n220), .C1(new_n236), .C2(new_n237), .ZN(new_n256));
  INV_X1    g055(.A(G227gat), .ZN(new_n257));
  INV_X1    g056(.A(G233gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT34), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT34), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n254), .A2(new_n256), .A3(new_n263), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G15gat), .B(G43gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT67), .ZN(new_n267));
  XNOR2_X1  g066(.A(G71gat), .B(G99gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(KEYINPUT24), .A3(new_n219), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n213), .A2(KEYINPUT23), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n211), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n272), .A2(new_n274), .A3(new_n222), .A4(new_n223), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n231), .B2(new_n230), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n228), .A2(new_n232), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT65), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n255), .B1(new_n280), .B2(new_n220), .ZN(new_n281));
  INV_X1    g080(.A(new_n219), .ZN(new_n282));
  AOI221_X4 g081(.A(new_n282), .B1(new_n217), .B2(new_n212), .C1(new_n207), .C2(new_n208), .ZN(new_n283));
  AOI211_X1 g082(.A(new_n253), .B(new_n283), .C1(new_n278), .C2(new_n279), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n259), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT33), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n270), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n254), .A2(new_n256), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT33), .B1(new_n289), .B2(new_n259), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n262), .B(new_n264), .C1(new_n290), .C2(new_n270), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n288), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n288), .B2(new_n291), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT68), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G228gat), .A2(G233gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT75), .ZN(new_n299));
  XOR2_X1   g098(.A(G211gat), .B(G218gat), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n301), .A2(KEYINPUT69), .ZN(new_n302));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303));
  INV_X1    g102(.A(G211gat), .ZN(new_n304));
  INV_X1    g103(.A(G218gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n303), .B1(KEYINPUT22), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n302), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310));
  INV_X1    g109(.A(G155gat), .ZN(new_n311));
  INV_X1    g110(.A(G162gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n311), .B2(new_n312), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT71), .B1(new_n315), .B2(G141gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n317));
  INV_X1    g116(.A(G141gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(G148gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n318), .A2(G148gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n315), .A2(G141gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n310), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(G155gat), .B(G162gat), .Z(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n322), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT29), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n309), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(new_n327), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT29), .B1(new_n307), .B2(new_n301), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n333), .B1(new_n301), .B2(new_n307), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n334), .B2(new_n323), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n299), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n323), .B1(new_n308), .B2(KEYINPUT29), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n331), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n309), .B2(new_n329), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n336), .B1(new_n339), .B2(new_n298), .ZN(new_n340));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT31), .B(G50gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(G22gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(G22gat), .B2(new_n343), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n340), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n295), .A2(new_n297), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n323), .B1(new_n322), .B2(new_n327), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT72), .B1(new_n328), .B2(new_n350), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n350), .A2(KEYINPUT72), .ZN(new_n352));
  INV_X1    g151(.A(new_n252), .ZN(new_n353));
  AOI21_X1  g152(.A(G134gat), .B1(new_n250), .B2(new_n251), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT73), .B1(new_n249), .B2(new_n252), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n351), .B(new_n352), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT4), .B1(new_n253), .B2(new_n331), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n332), .A2(new_n249), .A3(new_n360), .A4(new_n252), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n363), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n355), .B1(new_n353), .B2(new_n354), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n249), .A2(KEYINPUT73), .A3(new_n252), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n332), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n253), .A2(new_n331), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT5), .ZN(new_n372));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT0), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(G57gat), .ZN(new_n375));
  INV_X1    g174(.A(G85gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n372), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n380), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n379), .B1(new_n364), .B2(new_n370), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n377), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT6), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n372), .A2(KEYINPUT6), .A3(new_n378), .A4(new_n380), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT74), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n381), .A2(new_n384), .A3(KEYINPUT74), .A4(new_n385), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n280), .A2(new_n220), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n233), .A2(new_n235), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n220), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n393), .A2(KEYINPUT29), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n309), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n396), .A2(new_n392), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n238), .B2(new_n397), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n401), .B2(new_n309), .ZN(new_n402));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G64gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n404), .B(G92gat), .Z(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(KEYINPUT30), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n402), .B2(new_n405), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT70), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n406), .B(KEYINPUT70), .C1(new_n402), .C2(new_n405), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT30), .B1(new_n402), .B2(new_n405), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT35), .B1(new_n349), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n293), .A2(new_n294), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(new_n347), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n384), .A2(new_n385), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT79), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n381), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n382), .A2(new_n383), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT79), .B1(new_n424), .B2(new_n378), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n421), .B(KEYINPUT80), .C1(new_n423), .C2(new_n425), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n387), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT35), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n407), .A2(new_n411), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n420), .A2(new_n430), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(KEYINPUT83), .B(KEYINPUT35), .C1(new_n349), .C2(new_n414), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n358), .A2(new_n362), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n365), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n368), .A2(new_n369), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n437), .B(KEYINPUT39), .C1(new_n438), .C2(new_n365), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n437), .A2(KEYINPUT39), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n440), .A2(KEYINPUT77), .A3(new_n377), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT77), .B1(new_n440), .B2(new_n377), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT40), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT78), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(KEYINPUT78), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n446), .B(new_n439), .C1(new_n441), .C2(new_n442), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n423), .A2(new_n425), .ZN(new_n448));
  INV_X1    g247(.A(new_n432), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n445), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n394), .A2(new_n308), .A3(new_n398), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n238), .A2(new_n397), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n309), .B1(new_n453), .B2(new_n400), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n394), .A2(new_n455), .A3(new_n308), .A4(new_n398), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT37), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT38), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n405), .B1(new_n402), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n402), .A2(new_n405), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT38), .B1(new_n457), .B2(KEYINPUT37), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n459), .B1(new_n466), .B2(new_n462), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(new_n428), .A3(new_n387), .A4(new_n429), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n402), .A2(new_n461), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n460), .B1(new_n470), .B2(new_n462), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n348), .B(new_n450), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n389), .A2(new_n390), .B1(new_n408), .B2(new_n407), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n348), .B1(new_n473), .B2(new_n413), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n295), .B2(new_n297), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT36), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n435), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT84), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n435), .A2(new_n482), .A3(new_n479), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n484));
  INV_X1    g283(.A(G29gat), .ZN(new_n485));
  INV_X1    g284(.A(G36gat), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT14), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G43gat), .B(G50gat), .Z(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(KEYINPUT85), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(new_n489), .A3(new_n488), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n497));
  INV_X1    g296(.A(new_n494), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n496), .B(new_n497), .C1(KEYINPUT15), .C2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(KEYINPUT15), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(new_n492), .B2(new_n494), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT86), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n484), .B1(new_n504), .B2(KEYINPUT17), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT16), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(G1gat), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n508), .B(KEYINPUT88), .C1(G1gat), .C2(new_n506), .ZN(new_n509));
  INV_X1    g308(.A(G8gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT17), .B1(new_n500), .B2(new_n502), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT87), .A4(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n505), .A2(new_n511), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n504), .ZN(new_n517));
  INV_X1    g316(.A(new_n511), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT18), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT89), .B1(new_n504), .B2(new_n511), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n516), .B(KEYINPUT13), .Z(new_n525));
  NAND3_X1  g324(.A1(new_n517), .A2(KEYINPUT89), .A3(new_n518), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n515), .A2(KEYINPUT18), .A3(new_n516), .A4(new_n519), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G197gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT11), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(new_n209), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT12), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n522), .A2(new_n534), .A3(new_n527), .A4(new_n528), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n481), .A2(new_n483), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G99gat), .ZN(new_n544));
  INV_X1    g343(.A(G106gat), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT8), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT95), .B(G92gat), .Z(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(G85gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT96), .ZN(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G99gat), .B(G106gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n505), .A2(new_n512), .A3(new_n514), .A4(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G190gat), .B(G218gat), .Z(new_n556));
  INV_X1    g355(.A(new_n554), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n517), .ZN(new_n558));
  NAND3_X1  g357(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n555), .A2(new_n556), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT97), .ZN(new_n561));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT94), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n569));
  INV_X1    g368(.A(new_n556), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(KEYINPUT97), .A3(new_n560), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n566), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT98), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT98), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n568), .A2(new_n572), .A3(new_n576), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n571), .A2(new_n564), .A3(new_n560), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT21), .ZN(new_n582));
  XNOR2_X1  g381(.A(G57gat), .B(G64gat), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  OAI21_X1  g386(.A(new_n511), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT93), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n582), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n589), .B(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT91), .B(KEYINPUT92), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n595), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n581), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(G230gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(new_n258), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n549), .A2(KEYINPUT99), .A3(new_n551), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT99), .B1(new_n549), .B2(new_n551), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n553), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT100), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n552), .A2(new_n553), .ZN(new_n610));
  INV_X1    g409(.A(new_n587), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n612), .B(new_n553), .C1(new_n606), .C2(new_n607), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n609), .A2(new_n610), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n554), .A2(new_n587), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n557), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n605), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n605), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n620), .B1(new_n614), .B2(new_n616), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT101), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(new_n210), .ZN(new_n625));
  INV_X1    g424(.A(G204gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n622), .A2(KEYINPUT102), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n628), .B1(new_n622), .B2(KEYINPUT102), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n603), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n543), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n391), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g435(.A1(new_n543), .A2(new_n432), .A3(new_n632), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n507), .A2(new_n510), .ZN(new_n638));
  NAND2_X1  g437(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n640), .A2(new_n642), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT42), .B1(new_n637), .B2(new_n510), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT103), .B1(new_n645), .B2(new_n640), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(G1325gat));
  AOI21_X1  g446(.A(G15gat), .B1(new_n633), .B2(new_n418), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n476), .A2(new_n477), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n650), .A2(G15gat), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n648), .B1(new_n633), .B2(new_n651), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n633), .A2(new_n347), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT43), .B(G22gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NAND4_X1  g454(.A1(new_n481), .A2(new_n483), .A3(new_n541), .A4(new_n581), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n602), .A2(new_n631), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n485), .A3(new_n634), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n659), .A2(KEYINPUT45), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(KEYINPUT45), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n579), .B1(new_n575), .B2(new_n577), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n481), .A2(new_n483), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n480), .A2(new_n581), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n663), .ZN(new_n667));
  INV_X1    g466(.A(new_n538), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n657), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT104), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n665), .A2(new_n667), .A3(new_n672), .A4(new_n669), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n391), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OAI22_X1  g473(.A1(new_n660), .A2(new_n661), .B1(new_n674), .B2(new_n485), .ZN(G1328gat));
  NAND3_X1  g474(.A1(new_n658), .A2(new_n486), .A3(new_n449), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(KEYINPUT46), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(KEYINPUT46), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n432), .B1(new_n671), .B2(new_n673), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n677), .B(new_n678), .C1(new_n486), .C2(new_n679), .ZN(G1329gat));
  OAI21_X1  g479(.A(G43gat), .B1(new_n670), .B2(new_n649), .ZN(new_n681));
  INV_X1    g480(.A(G43gat), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n658), .A2(new_n682), .A3(new_n418), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n683), .A3(KEYINPUT47), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n671), .A2(new_n673), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n682), .B1(new_n686), .B2(new_n650), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(KEYINPUT105), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI211_X1 g488(.A(KEYINPUT105), .B(new_n682), .C1(new_n686), .C2(new_n650), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n684), .B1(new_n689), .B2(new_n690), .ZN(G1330gat));
  INV_X1    g490(.A(new_n657), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n542), .A2(KEYINPUT106), .A3(new_n581), .A4(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(G50gat), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n656), .B2(new_n657), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n693), .A2(new_n694), .A3(new_n696), .A4(new_n347), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT48), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n665), .A2(new_n667), .A3(new_n347), .A4(new_n669), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(G50gat), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n697), .A2(KEYINPUT107), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT107), .B1(new_n697), .B2(new_n700), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n694), .B1(new_n686), .B2(new_n347), .ZN(new_n704));
  INV_X1    g503(.A(new_n697), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n698), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(G1331gat));
  INV_X1    g506(.A(new_n631), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n603), .A2(new_n668), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT108), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n480), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n634), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g513(.A(new_n432), .B(KEYINPUT109), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT49), .B(G64gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n715), .ZN(new_n718));
  OAI22_X1  g517(.A1(new_n711), .A2(new_n718), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT110), .Z(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n711), .B2(new_n649), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n711), .A2(G71gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n419), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1334gat));
  NAND2_X1  g525(.A1(new_n712), .A2(new_n347), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n601), .A2(new_n538), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n480), .A2(new_n581), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT112), .Z(new_n733));
  NOR2_X1   g532(.A1(new_n631), .A2(new_n391), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n376), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n665), .A2(new_n667), .A3(new_n729), .ZN(new_n736));
  INV_X1    g535(.A(new_n734), .ZN(new_n737));
  OAI21_X1  g536(.A(G85gat), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(G1336gat));
  NAND4_X1  g538(.A1(new_n665), .A2(new_n667), .A3(new_n708), .A4(new_n729), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n740), .A2(KEYINPUT116), .A3(new_n718), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT116), .B1(new_n740), .B2(new_n718), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(new_n547), .A3(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n631), .A2(new_n718), .A3(G92gat), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT52), .B1(new_n732), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT113), .B1(new_n731), .B2(KEYINPUT114), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n730), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT114), .B1(new_n749), .B2(KEYINPUT113), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n744), .B(new_n748), .C1(new_n750), .C2(KEYINPUT51), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n547), .B1(new_n740), .B2(new_n432), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n753), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT115), .B1(new_n753), .B2(KEYINPUT52), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n746), .B1(new_n754), .B2(new_n755), .ZN(G1337gat));
  NAND4_X1  g555(.A1(new_n733), .A2(new_n544), .A3(new_n418), .A4(new_n708), .ZN(new_n757));
  OAI21_X1  g556(.A(G99gat), .B1(new_n740), .B2(new_n649), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1338gat));
  OR2_X1    g558(.A1(new_n740), .A2(new_n348), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G106gat), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n631), .A2(G106gat), .A3(new_n348), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT53), .B1(new_n732), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n750), .A2(KEYINPUT51), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n730), .B2(new_n747), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n766), .A2(new_n762), .B1(G106gat), .B2(new_n760), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n764), .B1(new_n767), .B2(new_n768), .ZN(G1339gat));
  NAND2_X1  g568(.A1(new_n617), .A2(new_n618), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n620), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n617), .A2(new_n605), .A3(new_n618), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(KEYINPUT54), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n627), .B1(new_n619), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n622), .A2(new_n627), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n773), .A2(KEYINPUT55), .A3(new_n775), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n778), .A2(new_n538), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n516), .B1(new_n515), .B2(new_n519), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n525), .B1(new_n524), .B2(new_n526), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n533), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT117), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n786), .B(new_n533), .C1(new_n782), .C2(new_n783), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n537), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n629), .A3(new_n630), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n581), .B1(new_n781), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n662), .A2(new_n792), .A3(new_n788), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n602), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NOR4_X1   g593(.A1(new_n581), .A2(new_n708), .A3(new_n602), .A4(new_n538), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n715), .A2(new_n391), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n420), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n242), .B1(new_n801), .B2(new_n541), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT118), .ZN(new_n803));
  INV_X1    g602(.A(new_n799), .ZN(new_n804));
  INV_X1    g603(.A(new_n349), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n806), .A2(G113gat), .A3(new_n668), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n803), .A2(new_n807), .ZN(G1340gat));
  INV_X1    g607(.A(new_n801), .ZN(new_n809));
  OAI21_X1  g608(.A(G120gat), .B1(new_n809), .B2(new_n631), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n708), .A2(new_n240), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n806), .B2(new_n811), .ZN(G1341gat));
  NAND3_X1  g611(.A1(new_n801), .A2(G127gat), .A3(new_n601), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n801), .A2(KEYINPUT119), .A3(G127gat), .A4(new_n601), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n245), .B1(new_n806), .B2(new_n602), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n815), .A2(new_n817), .A3(KEYINPUT120), .A4(new_n816), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1342gat));
  OR3_X1    g621(.A1(new_n662), .A2(new_n792), .A3(new_n788), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n781), .A2(new_n790), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n662), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n795), .B1(new_n826), .B2(new_n602), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n391), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n828), .A2(new_n432), .A3(new_n805), .A4(new_n581), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT56), .B1(new_n829), .B2(G134gat), .ZN(new_n830));
  OAI21_X1  g629(.A(G134gat), .B1(new_n809), .B2(new_n662), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n829), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n830), .B(new_n831), .C1(new_n834), .C2(new_n835), .ZN(G1343gat));
  AOI21_X1  g635(.A(new_n348), .B1(new_n794), .B2(new_n796), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT122), .B1(new_n837), .B2(KEYINPUT57), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n839), .B(new_n840), .C1(new_n827), .C2(new_n348), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n790), .B1(new_n540), .B2(new_n792), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n662), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n601), .B1(new_n843), .B2(new_n823), .ZN(new_n844));
  OAI211_X1 g643(.A(KEYINPUT57), .B(new_n347), .C1(new_n844), .C2(new_n795), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n838), .A2(new_n841), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n649), .A2(new_n798), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n541), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(G141gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n827), .A2(new_n348), .A3(new_n847), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n851), .A2(new_n318), .A3(new_n541), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n852), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n846), .A2(new_n538), .A3(new_n848), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT58), .A3(G141gat), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n855), .A2(new_n856), .B1(new_n857), .B2(new_n859), .ZN(G1344gat));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n848), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n861), .B(G148gat), .C1(new_n862), .C2(new_n631), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT57), .B1(new_n827), .B2(new_n348), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n632), .A2(new_n541), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n840), .B(new_n347), .C1(new_n844), .C2(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n864), .A2(new_n866), .A3(new_n708), .A4(new_n848), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G148gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT59), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n315), .A3(new_n708), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1345gat));
  AOI21_X1  g671(.A(G155gat), .B1(new_n851), .B2(new_n601), .ZN(new_n873));
  INV_X1    g672(.A(new_n862), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n601), .A2(G155gat), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT124), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(G1346gat));
  OAI21_X1  g676(.A(G162gat), .B1(new_n862), .B2(new_n662), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n828), .A2(new_n432), .A3(new_n581), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n650), .A2(new_n348), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n312), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n878), .B1(new_n879), .B2(new_n881), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n827), .A2(new_n634), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n805), .A2(new_n715), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT125), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n884), .A2(KEYINPUT125), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n209), .A3(new_n538), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n634), .A2(new_n432), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n797), .A2(new_n420), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G169gat), .B1(new_n890), .B2(new_n540), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(G1348gat));
  NOR3_X1   g691(.A1(new_n890), .A2(new_n210), .A3(new_n631), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n887), .A2(new_n708), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n210), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n887), .A2(new_n202), .A3(new_n601), .ZN(new_n896));
  OAI21_X1  g695(.A(G183gat), .B1(new_n890), .B2(new_n602), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n890), .B2(new_n662), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT61), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n887), .A2(new_n203), .A3(new_n581), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1351gat));
  NAND3_X1  g702(.A1(new_n883), .A2(new_n715), .A3(new_n880), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(G197gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n906), .A3(new_n538), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n864), .A2(new_n866), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n649), .A2(new_n889), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(new_n541), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n907), .B1(new_n911), .B2(new_n906), .ZN(G1352gat));
  NOR3_X1   g711(.A1(new_n904), .A2(G204gat), .A3(new_n631), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n908), .A2(new_n708), .A3(new_n909), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n915), .B(new_n916), .C1(new_n626), .C2(new_n917), .ZN(G1353gat));
  NAND3_X1  g717(.A1(new_n905), .A2(new_n304), .A3(new_n601), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n908), .A2(new_n601), .A3(new_n909), .ZN(new_n920));
  AND3_X1   g719(.A1(new_n920), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT63), .B1(new_n920), .B2(G211gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(G1354gat));
  AOI21_X1  g722(.A(G218gat), .B1(new_n905), .B2(new_n581), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n662), .A2(new_n305), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT126), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n910), .B2(new_n926), .ZN(G1355gat));
endmodule


