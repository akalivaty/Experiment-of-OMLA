//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(new_n211), .B2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n210), .A2(KEYINPUT64), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n209), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n225), .B(new_n232), .C1(new_n234), .C2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(G223), .B1(new_n262), .B2(G77), .ZN(new_n263));
  INV_X1    g0063(.A(G222), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1698), .B1(new_n257), .B2(new_n258), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  OAI211_X1 g0069(.A(G1), .B(G13), .C1(new_n256), .C2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n267), .A2(new_n268), .B1(G226), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n270), .A2(G274), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT67), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT67), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G45), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n279), .A3(new_n269), .ZN(new_n280));
  AND3_X1   g0080(.A1(new_n280), .A2(KEYINPUT68), .A3(new_n208), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT68), .B1(new_n280), .B2(new_n208), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n275), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT69), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n274), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G58), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT8), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT8), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G58), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n209), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n209), .A2(new_n256), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n296), .A2(new_n298), .B1(new_n300), .B2(G150), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT70), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n301), .A2(new_n302), .B1(G20), .B2(new_n203), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n302), .B2(new_n301), .ZN(new_n304));
  NAND3_X1  g0104(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n233), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n228), .A2(new_n209), .A3(G1), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n306), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n309), .A2(new_n310), .B1(new_n202), .B2(new_n308), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n288), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n291), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n312), .B(KEYINPUT9), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT72), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n318), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n289), .A2(G200), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT10), .B1(new_n288), .B2(G190), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n319), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n321), .B(new_n317), .C1(new_n289), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT10), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n316), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n213), .A2(G20), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n328), .B1(new_n297), .B2(new_n219), .C1(new_n202), .C2(new_n299), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n306), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT11), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n228), .A2(G1), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G20), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT71), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n308), .A2(KEYINPUT71), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n306), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n208), .A2(G20), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n337), .A2(G68), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n331), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT12), .B1(new_n337), .B2(G68), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT74), .ZN(new_n343));
  INV_X1    g0143(.A(new_n332), .ZN(new_n344));
  OR3_X1    g0144(.A1(new_n344), .A2(KEYINPUT12), .A3(new_n328), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n341), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n273), .A2(G238), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n283), .A2(new_n348), .ZN(new_n349));
  OR2_X1    g0149(.A1(G226), .A2(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G232), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G1698), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n350), .B(new_n352), .C1(new_n260), .C2(new_n261), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT73), .B1(new_n355), .B2(new_n268), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n357), .B(new_n270), .C1(new_n353), .C2(new_n354), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT13), .B1(new_n349), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n280), .A2(new_n208), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT68), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n280), .A2(KEYINPUT68), .A3(new_n208), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n275), .B1(G238), .B2(new_n273), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n355), .A2(new_n268), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n357), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n355), .A2(KEYINPUT73), .A3(new_n268), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n360), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(G169), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n360), .A2(new_n372), .A3(G179), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n373), .B2(G169), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n347), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n373), .A2(G200), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n360), .A2(new_n372), .A3(G190), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n346), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n265), .A2(G232), .B1(new_n262), .B2(G107), .ZN(new_n384));
  INV_X1    g0184(.A(new_n259), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n214), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n268), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n283), .C1(new_n220), .C2(new_n272), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n290), .ZN(new_n389));
  INV_X1    g0189(.A(new_n296), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n390), .A2(new_n299), .B1(new_n209), .B2(new_n219), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT15), .B(G87), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n297), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n306), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n337), .A2(G77), .A3(new_n338), .A4(new_n339), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n394), .B(new_n395), .C1(G77), .C2(new_n337), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n388), .A2(G179), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n388), .B2(G200), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n388), .A2(new_n324), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n397), .A2(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n327), .A2(new_n383), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n272), .A2(new_n351), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n283), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT78), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n265), .A2(new_n406), .A3(G223), .ZN(new_n407));
  OAI211_X1 g0207(.A(G223), .B(new_n254), .C1(new_n260), .C2(new_n261), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT78), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n259), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n270), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(G169), .B1(new_n405), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n403), .B1(new_n365), .B2(new_n275), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n406), .B1(new_n265), .B2(G223), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n408), .A2(KEYINPUT78), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n411), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n268), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(G179), .A3(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n413), .A2(new_n419), .A3(KEYINPUT79), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT79), .B1(new_n413), .B2(new_n419), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n309), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n296), .A2(new_n339), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n423), .A2(new_n424), .B1(new_n333), .B2(new_n296), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT77), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n260), .B2(new_n261), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n257), .A2(KEYINPUT75), .A3(new_n258), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n209), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT7), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n258), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G68), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n292), .A2(new_n213), .ZN(new_n437));
  OAI21_X1  g0237(.A(G20), .B1(new_n437), .B2(new_n201), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n300), .A2(G159), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT16), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n338), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n257), .A2(new_n209), .A3(new_n258), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n432), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(KEYINPUT76), .A3(new_n434), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n262), .A2(new_n445), .A3(KEYINPUT7), .A4(new_n209), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(G68), .A3(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n438), .A2(new_n439), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT16), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n427), .B1(new_n441), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n434), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n431), .B2(new_n432), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n440), .B1(new_n454), .B2(new_n213), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n306), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT16), .B1(new_n447), .B2(new_n448), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT77), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n426), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT18), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n422), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n405), .A2(new_n412), .A3(new_n313), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n290), .B1(new_n414), .B2(new_n418), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n413), .A2(new_n419), .A3(KEYINPUT79), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n451), .A2(new_n427), .A3(new_n306), .A4(new_n455), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT77), .B1(new_n456), .B2(new_n457), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n425), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT18), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G200), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n405), .B2(new_n412), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n414), .A2(new_n324), .A3(new_n418), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n426), .B(new_n475), .C1(new_n452), .C2(new_n458), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT17), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(KEYINPUT17), .A3(new_n475), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n461), .A2(new_n471), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n402), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n265), .A2(KEYINPUT4), .A3(G244), .ZN(new_n482));
  OAI211_X1 g0282(.A(G244), .B(new_n254), .C1(new_n260), .C2(new_n261), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n259), .A2(G250), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n482), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n268), .ZN(new_n489));
  XNOR2_X1  g0289(.A(KEYINPUT5), .B(G41), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n276), .A2(G1), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(G257), .A3(new_n270), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n490), .A2(new_n270), .A3(G274), .A4(new_n491), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n489), .A2(new_n496), .A3(new_n313), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(new_n268), .B2(new_n488), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(G169), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n308), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n208), .A2(G33), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n309), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n503), .B2(new_n500), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n444), .A2(G107), .A3(new_n446), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n221), .A2(KEYINPUT6), .A3(G97), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n500), .A2(new_n221), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n205), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n506), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(G20), .B1(G77), .B2(new_n300), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n504), .B1(new_n511), .B2(new_n306), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n499), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n489), .A2(new_n496), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT81), .B1(new_n514), .B2(new_n324), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT81), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n498), .A2(new_n516), .A3(G190), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(KEYINPUT80), .A3(G200), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT80), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n498), .B2(new_n472), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(new_n522), .A3(new_n512), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n518), .A2(new_n522), .A3(KEYINPUT82), .A4(new_n512), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n513), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT89), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n257), .A2(new_n258), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(G257), .A3(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n531), .C1(new_n266), .C2(new_n216), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n268), .B1(new_n491), .B2(new_n490), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n532), .A2(new_n268), .B1(new_n533), .B2(G264), .ZN(new_n534));
  AOI21_X1  g0334(.A(G200), .B1(new_n534), .B2(new_n494), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n494), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n324), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n529), .A2(new_n209), .A3(G87), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT22), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT22), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n529), .A2(new_n540), .A3(new_n209), .A4(G87), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT24), .ZN(new_n543));
  INV_X1    g0343(.A(G116), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n256), .A2(new_n544), .A3(G20), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n209), .A2(G107), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n546), .A2(KEYINPUT23), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(KEYINPUT23), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n542), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n543), .B1(new_n542), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n306), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT87), .ZN(new_n553));
  OR2_X1    g0353(.A1(new_n553), .A2(KEYINPUT25), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(KEYINPUT25), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n554), .A2(new_n332), .A3(new_n546), .A4(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n332), .A2(new_n546), .ZN(new_n557));
  OAI221_X1 g0357(.A(new_n556), .B1(new_n555), .B2(new_n557), .C1(new_n503), .C2(new_n221), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n528), .B1(new_n537), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n534), .A2(new_n324), .A3(new_n494), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n536), .B2(G200), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(KEYINPUT89), .A3(new_n552), .A4(new_n559), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n534), .A2(new_n494), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G169), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n534), .A2(G179), .A3(new_n494), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT88), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n568), .A2(new_n569), .B1(new_n552), .B2(new_n559), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(KEYINPUT88), .A3(new_n567), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n561), .A2(new_n564), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n529), .A2(G257), .A3(new_n254), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n262), .A2(G303), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n385), .C2(new_n222), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT84), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n268), .ZN(new_n577));
  INV_X1    g0377(.A(new_n492), .ZN(new_n578));
  AOI22_X1  g0378(.A1(G270), .A2(new_n533), .B1(new_n578), .B2(new_n275), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n576), .B1(new_n575), .B2(new_n268), .ZN(new_n581));
  OAI21_X1  g0381(.A(G200), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n337), .A2(G116), .A3(new_n338), .A4(new_n502), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n305), .A2(new_n233), .B1(G20), .B2(new_n544), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n487), .B(new_n209), .C1(G33), .C2(new_n500), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT85), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n584), .A2(new_n585), .B1(new_n586), .B2(KEYINPUT20), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n586), .B2(KEYINPUT20), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT20), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n584), .A2(KEYINPUT85), .A3(new_n585), .A4(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n335), .A2(new_n336), .A3(new_n544), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n583), .A2(new_n588), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n575), .A2(new_n268), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT84), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n577), .A3(new_n579), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n582), .B(new_n593), .C1(new_n324), .C2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n580), .A2(new_n581), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n592), .A2(G169), .ZN(new_n600));
  OAI211_X1 g0400(.A(KEYINPUT86), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n580), .A2(new_n313), .A3(new_n581), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n592), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n598), .A2(KEYINPUT86), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n596), .A2(G169), .A3(new_n604), .A4(new_n592), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n597), .A2(new_n601), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G244), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n607));
  OAI211_X1 g0407(.A(G238), .B(new_n254), .C1(new_n260), .C2(new_n261), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(new_n256), .C2(new_n544), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n268), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n491), .A2(new_n216), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n275), .A2(new_n491), .B1(new_n270), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT83), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n313), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n529), .A2(new_n209), .A3(G68), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT19), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n209), .B1(new_n354), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(G87), .B2(new_n206), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n297), .B2(new_n500), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n618), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n306), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n335), .A2(new_n336), .A3(new_n392), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n625), .C1(new_n392), .C2(new_n503), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n610), .A2(KEYINPUT83), .A3(new_n612), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT83), .B1(new_n610), .B2(new_n612), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n617), .B(new_n626), .C1(new_n629), .C2(G169), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n615), .A2(G190), .A3(new_n616), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n625), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n503), .A2(new_n215), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n631), .B(new_n634), .C1(new_n629), .C2(new_n472), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n606), .A2(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n481), .A2(new_n527), .A3(new_n572), .A4(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n525), .A2(new_n526), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n613), .A2(new_n290), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT90), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT90), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n613), .A2(new_n642), .A3(new_n290), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n617), .A2(new_n641), .A3(new_n626), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n613), .A2(G200), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n631), .A2(new_n634), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n561), .B2(new_n564), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n603), .A2(new_n605), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n568), .A2(new_n560), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n601), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n513), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n639), .A2(new_n648), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n630), .A2(new_n635), .A3(new_n513), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n513), .A2(new_n644), .A3(new_n646), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n644), .B1(new_n656), .B2(KEYINPUT26), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n481), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n413), .A2(new_n419), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n459), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n460), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n459), .A2(new_n661), .A3(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n379), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n397), .A2(new_n398), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n666), .B1(new_n382), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n478), .A2(new_n479), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n323), .A2(new_n326), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n316), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n660), .A2(new_n673), .ZN(G369));
  NAND2_X1  g0474(.A1(new_n649), .A2(new_n601), .ZN(new_n675));
  OR3_X1    g0475(.A1(new_n344), .A2(KEYINPUT27), .A3(G20), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT27), .B1(new_n344), .B2(G20), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(KEYINPUT91), .B(G343), .Z(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n593), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n606), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n560), .A2(new_n680), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n570), .A2(new_n571), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n572), .A2(new_n686), .B1(new_n688), .B2(new_n680), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n572), .A2(new_n675), .A3(new_n681), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n568), .A2(new_n560), .A3(new_n681), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT92), .Z(G399));
  INV_X1    g0495(.A(new_n230), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n697), .A2(new_n208), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n236), .B2(new_n697), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  OAI211_X1 g0502(.A(new_n527), .B(new_n648), .C1(new_n688), .C2(new_n675), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n644), .B1(new_n654), .B2(KEYINPUT26), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(KEYINPUT26), .B2(new_n656), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n680), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n659), .A2(new_n681), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n498), .A2(new_n534), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n602), .A2(KEYINPUT30), .A3(new_n712), .A4(new_n629), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n615), .A2(new_n498), .A3(new_n616), .A4(new_n534), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n595), .A2(G179), .A3(new_n577), .A4(new_n579), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(G179), .B1(new_n610), .B2(new_n612), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n596), .A2(new_n514), .A3(new_n718), .A4(new_n565), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n713), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n720), .B2(new_n680), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(KEYINPUT93), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n527), .A2(new_n572), .A3(new_n637), .A4(new_n681), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT93), .ZN(new_n727));
  OAI21_X1  g0527(.A(G330), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n711), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n702), .B1(new_n730), .B2(G1), .ZN(G364));
  INV_X1    g0531(.A(new_n685), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n228), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n208), .B1(new_n733), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n697), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G330), .B2(new_n684), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n290), .A2(KEYINPUT95), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n209), .B1(KEYINPUT95), .B2(new_n290), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n233), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n209), .A2(G190), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT96), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n744), .A2(KEYINPUT96), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G159), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT32), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n209), .A2(new_n313), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n209), .B1(new_n746), .B2(G190), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n213), .B1(new_n756), .B2(new_n500), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n753), .A2(new_n324), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n757), .B1(G50), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n209), .A2(new_n324), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n313), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n529), .B1(new_n762), .B2(new_n292), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n472), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n744), .A2(new_n761), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n765), .A2(new_n215), .B1(new_n766), .B2(new_n219), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n745), .A2(new_n747), .A3(new_n764), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n763), .B(new_n767), .C1(new_n769), .C2(G107), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n751), .A2(new_n759), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n758), .ZN(new_n772));
  INV_X1    g0572(.A(G326), .ZN(new_n773));
  INV_X1    g0573(.A(G294), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n772), .A2(new_n773), .B1(new_n756), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n775), .B1(new_n754), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n748), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G329), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n769), .A2(G283), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n762), .A2(new_n781), .B1(new_n766), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n765), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n529), .B(new_n783), .C1(G303), .C2(new_n784), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n777), .A2(new_n779), .A3(new_n780), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n743), .B1(new_n771), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n230), .A2(new_n529), .ZN(new_n788));
  INV_X1    g0588(.A(G355), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n788), .A2(new_n789), .B1(G116), .B2(new_n230), .ZN(new_n790));
  INV_X1    g0590(.A(new_n236), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n277), .A2(new_n279), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G45), .B2(new_n252), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n429), .A2(new_n430), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n696), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n790), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT94), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n742), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n736), .B1(new_n797), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n787), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n800), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n684), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n738), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(G396));
  INV_X1    g0608(.A(new_n799), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n742), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n735), .B(new_n697), .C1(new_n219), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n756), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n758), .A2(G303), .B1(G97), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n766), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G107), .A2(new_n784), .B1(new_n814), .B2(G116), .ZN(new_n815));
  INV_X1    g0615(.A(new_n762), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n529), .B1(new_n816), .B2(G294), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n813), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n769), .A2(G87), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n782), .B2(new_n748), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n755), .A2(KEYINPUT97), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n755), .A2(KEYINPUT97), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n818), .B(new_n820), .C1(new_n824), .C2(G283), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n795), .B1(new_n748), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT98), .Z(new_n828));
  NAND2_X1  g0628(.A1(new_n769), .A2(G68), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n829), .B1(new_n202), .B2(new_n765), .C1(new_n292), .C2(new_n756), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G143), .A2(new_n816), .B1(new_n814), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n772), .B2(new_n834), .C1(new_n835), .C2(new_n755), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT34), .Z(new_n837));
  NOR2_X1   g0637(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n825), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT100), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n667), .B2(new_n681), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n397), .A2(KEYINPUT100), .A3(new_n398), .A4(new_n680), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n396), .A2(new_n680), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n401), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n811), .B1(new_n743), .B2(new_n840), .C1(new_n847), .C2(new_n799), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n842), .A2(new_n843), .B1(new_n401), .B2(new_n845), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n709), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n659), .A2(new_n681), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n728), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(new_n736), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT101), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n852), .A2(new_n728), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n854), .A2(KEYINPUT101), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n848), .B1(new_n857), .B2(new_n858), .ZN(G384));
  OR2_X1    g0659(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n509), .A2(KEYINPUT35), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n860), .A2(G116), .A3(new_n234), .A4(new_n861), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT36), .Z(new_n863));
  NOR3_X1   g0663(.A1(new_n791), .A2(new_n219), .A3(new_n437), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(KEYINPUT102), .B1(new_n202), .B2(G68), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(KEYINPUT102), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n208), .A2(G13), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n481), .B1(new_n708), .B2(new_n710), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n673), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT106), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT16), .B1(new_n436), .B2(new_n448), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n426), .B1(new_n872), .B2(new_n456), .ZN(new_n873));
  INV_X1    g0673(.A(new_n678), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n461), .A2(new_n471), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n876), .B2(new_n670), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n459), .B1(new_n422), .B2(new_n874), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT37), .B1(new_n470), .B2(new_n475), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n873), .B1(new_n661), .B2(new_n874), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n476), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n480), .A2(new_n875), .B1(new_n880), .B2(new_n883), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(KEYINPUT38), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n877), .A2(new_n884), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(KEYINPUT104), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT39), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n666), .A2(new_n681), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n459), .A2(new_n874), .ZN(new_n898));
  INV_X1    g0698(.A(new_n670), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(new_n665), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n476), .A2(KEYINPUT105), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n662), .A2(new_n898), .A3(KEYINPUT105), .A4(new_n476), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n903), .A2(new_n904), .B1(new_n879), .B2(new_n878), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n892), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT39), .B1(new_n906), .B2(new_n885), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n895), .A2(new_n897), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT104), .B1(new_n888), .B2(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n891), .A2(new_n892), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT103), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n373), .A2(G169), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT14), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n382), .A2(new_n915), .A3(new_n376), .A4(new_n375), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n346), .A2(new_n681), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n917), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n379), .A2(new_n382), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n379), .A2(new_n913), .A3(new_n382), .A4(new_n919), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n667), .A2(new_n680), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n923), .B1(new_n851), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n912), .A2(new_n926), .A3(new_n893), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n663), .A2(new_n664), .A3(new_n678), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n909), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n871), .B(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n921), .A2(new_n847), .A3(new_n922), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n723), .A2(new_n721), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n725), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n912), .A2(new_n893), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n906), .B2(new_n885), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n935), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(G330), .A3(new_n940), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n402), .A2(new_n480), .A3(new_n934), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(G330), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n936), .A2(new_n937), .B1(new_n935), .B2(new_n939), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n944), .A2(KEYINPUT107), .B1(new_n945), .B2(new_n942), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(KEYINPUT107), .B2(new_n944), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n931), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n208), .B2(new_n733), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n931), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n868), .B1(new_n949), .B2(new_n950), .ZN(G367));
  OAI21_X1  g0751(.A(new_n527), .B1(new_n512), .B2(new_n681), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n513), .A2(new_n680), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n955), .A2(KEYINPUT42), .A3(new_n691), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n687), .B1(new_n525), .B2(new_n526), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n681), .B1(new_n957), .B2(new_n513), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT42), .B1(new_n955), .B2(new_n691), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n680), .B1(new_n632), .B2(new_n633), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n644), .A2(new_n646), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n644), .B2(new_n961), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n960), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n967), .B1(new_n960), .B2(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(new_n690), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(new_n955), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n969), .A2(new_n970), .B1(KEYINPUT110), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT110), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n972), .ZN(new_n976));
  OAI211_X1 g0776(.A(KEYINPUT110), .B(new_n973), .C1(new_n969), .C2(new_n970), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n697), .B(KEYINPUT41), .Z(new_n978));
  AOI21_X1  g0778(.A(new_n954), .B1(new_n692), .B2(new_n691), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT44), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n955), .B2(new_n693), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n954), .A2(KEYINPUT45), .A3(new_n692), .A4(new_n691), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT112), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n982), .A2(new_n983), .B1(new_n984), .B2(new_n690), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n971), .A2(KEYINPUT112), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n980), .A2(new_n987), .A3(new_n985), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n675), .A2(new_n681), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n689), .A2(KEYINPUT111), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n691), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT111), .B1(new_n689), .B2(new_n992), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(new_n732), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n732), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n729), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n991), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n978), .B1(new_n1000), .B2(new_n730), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n976), .B(new_n977), .C1(new_n1001), .C2(new_n735), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n796), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n245), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n801), .B1(new_n230), .B2(new_n392), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n736), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n765), .A2(new_n544), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(KEYINPUT46), .A2(new_n1007), .B1(new_n758), .B2(G311), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(KEYINPUT46), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G107), .B2(new_n812), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(new_n823), .C2(new_n774), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n769), .A2(G97), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n778), .A2(G317), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G303), .A2(new_n816), .B1(new_n814), .B2(G283), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n795), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n762), .A2(new_n835), .B1(new_n766), .B2(new_n202), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n262), .B(new_n1017), .C1(G58), .C2(new_n784), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G77), .A2(new_n769), .B1(new_n778), .B2(G137), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n756), .A2(new_n213), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n758), .B2(G143), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n823), .A2(new_n749), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1011), .A2(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT47), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1006), .B1(new_n1025), .B2(new_n742), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n963), .A2(new_n805), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1002), .A2(new_n1028), .ZN(G387));
  OAI22_X1  g0829(.A1(new_n788), .A2(new_n698), .B1(G107), .B2(new_n230), .ZN(new_n1030));
  XOR2_X1   g0830(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n390), .B2(G50), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n390), .A2(new_n1031), .A3(G50), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n276), .B1(new_n213), .B2(new_n219), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1033), .A2(new_n699), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1003), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n242), .A2(new_n792), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1030), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n392), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n754), .A2(new_n296), .B1(new_n1039), .B2(new_n812), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n795), .C1(new_n749), .C2(new_n772), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n765), .A2(new_n219), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G68), .B2(new_n814), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1012), .B(new_n1043), .C1(new_n202), .C2(new_n762), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1041), .B(new_n1044), .C1(G150), .C2(new_n778), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G317), .A2(new_n816), .B1(new_n814), .B2(G303), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n781), .B2(new_n772), .C1(new_n823), .C2(new_n782), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n784), .A2(G294), .B1(new_n812), .B2(G283), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1015), .B1(new_n768), .B2(new_n544), .C1(new_n773), .C2(new_n748), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1045), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n736), .B1(new_n802), .B2(new_n1038), .C1(new_n1058), .C2(new_n743), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT114), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n689), .B2(new_n800), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n997), .A2(new_n998), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n735), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n730), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n697), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1062), .A2(new_n730), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(G393));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n989), .A3(new_n990), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1000), .A2(new_n1068), .A3(new_n697), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1003), .A2(new_n249), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n801), .B1(new_n500), .B2(new_n230), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n784), .A2(G68), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n814), .A2(new_n296), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n812), .A2(G77), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n795), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(G143), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n819), .B1(new_n1076), .B2(new_n748), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1075), .B(new_n1077), .C1(new_n824), .C2(G50), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n758), .A2(G150), .B1(new_n816), .B2(G159), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT51), .Z(new_n1080));
  AOI21_X1  g0880(.A(new_n529), .B1(new_n784), .B2(G283), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n544), .B2(new_n756), .C1(new_n774), .C2(new_n766), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n221), .A2(new_n768), .B1(new_n748), .B2(new_n781), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(new_n824), .C2(G303), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n758), .A2(G317), .B1(new_n816), .B2(G311), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT52), .Z(new_n1086));
  AOI22_X1  g0886(.A1(new_n1078), .A2(new_n1080), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n736), .B1(new_n1070), .B2(new_n1071), .C1(new_n1087), .C2(new_n743), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n955), .B2(new_n800), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n991), .B2(new_n735), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1069), .A2(new_n1090), .ZN(G390));
  INV_X1    g0891(.A(KEYINPUT39), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n912), .B2(new_n893), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n907), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1094), .A2(new_n799), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n810), .ZN(new_n1096));
  INV_X1    g0896(.A(G283), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n772), .A2(new_n1097), .B1(new_n766), .B2(new_n500), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n824), .B2(G107), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT119), .Z(new_n1100));
  OAI221_X1 g0900(.A(new_n262), .B1(new_n762), .B2(new_n544), .C1(new_n215), .C2(new_n765), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n829), .B1(new_n774), .B2(new_n748), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(G77), .C2(new_n812), .ZN(new_n1103));
  OR3_X1    g0903(.A1(new_n765), .A2(KEYINPUT53), .A3(new_n835), .ZN(new_n1104));
  OAI21_X1  g0904(.A(KEYINPUT53), .B1(new_n765), .B2(new_n835), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(new_n749), .C2(new_n756), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G132), .A2(new_n816), .B1(new_n814), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(G125), .ZN(new_n1110));
  INV_X1    g0910(.A(G128), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n748), .C1(new_n1111), .C2(new_n772), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1106), .B(new_n1112), .C1(new_n824), .C2(G137), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n529), .B1(new_n768), .B2(new_n202), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT118), .Z(new_n1115));
  AOI22_X1  g0915(.A1(new_n1100), .A2(new_n1103), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n736), .B1(new_n296), .B2(new_n1096), .C1(new_n1116), .C2(new_n743), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1095), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT116), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n935), .A2(new_n1119), .A3(G330), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n725), .A2(new_n933), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1121), .A2(new_n847), .A3(new_n921), .A4(new_n922), .ZN(new_n1122));
  INV_X1    g0922(.A(G330), .ZN(new_n1123));
  OAI21_X1  g0923(.A(KEYINPUT116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n926), .A2(new_n897), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n1093), .B2(new_n907), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n923), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n680), .B(new_n849), .C1(new_n705), .C2(new_n703), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n924), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT115), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n896), .B(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n885), .B2(new_n906), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1126), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT117), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n926), .A2(new_n897), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n895), .B2(new_n908), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n728), .A2(new_n849), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1129), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1137), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1131), .A2(new_n1134), .B1(new_n1140), .B2(new_n1129), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1128), .A2(KEYINPUT117), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1136), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1118), .B1(new_n1146), .B2(new_n735), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n943), .A2(new_n869), .A3(new_n673), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n923), .B1(new_n728), .B2(new_n849), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1120), .A2(new_n1149), .A3(new_n1124), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n851), .A2(new_n925), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1130), .A2(new_n924), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n847), .A2(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n923), .B1(new_n934), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1141), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1148), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n697), .B1(new_n1146), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1135), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1125), .B1(new_n1139), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1128), .A2(KEYINPUT117), .A3(new_n1144), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT117), .B1(new_n1128), .B2(new_n1144), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1160), .B(new_n1157), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1147), .B1(new_n1158), .B2(new_n1164), .ZN(G378));
  XNOR2_X1  g0965(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n312), .A2(new_n874), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n327), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n327), .A2(new_n1168), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1171), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n1169), .A3(new_n1166), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n809), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n736), .B1(G50), .B2(new_n1096), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n755), .A2(new_n826), .B1(new_n756), .B2(new_n835), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n784), .A2(new_n1108), .B1(new_n816), .B2(G128), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n834), .B2(new_n766), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G125), .C2(new_n758), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n256), .B(new_n269), .C1(new_n768), .C2(new_n749), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G124), .B2(new_n778), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n768), .A2(new_n292), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n762), .A2(new_n221), .B1(new_n766), .B2(new_n392), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1188), .A2(new_n1189), .A3(G41), .A4(new_n1042), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1097), .B2(new_n748), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n755), .A2(new_n500), .B1(new_n772), .B2(new_n544), .ZN(new_n1192));
  NOR4_X1   g0992(.A1(new_n1191), .A2(new_n795), .A3(new_n1020), .A4(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n269), .B1(new_n1015), .B2(new_n256), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n202), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1193), .A2(KEYINPUT58), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1187), .A2(new_n1194), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1177), .B1(new_n1198), .B2(new_n742), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1176), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT120), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n909), .B2(new_n929), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n941), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n945), .A2(new_n1175), .A3(G330), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1204), .A2(new_n1205), .B1(new_n930), .B2(KEYINPUT120), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1200), .B1(new_n1208), .B2(new_n734), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n697), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n941), .A2(new_n1203), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1175), .B1(new_n945), .B2(G330), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n930), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n927), .A2(new_n928), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1094), .B2(new_n897), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1204), .A2(new_n1215), .A3(new_n1205), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1213), .A2(KEYINPUT57), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1148), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1163), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1210), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT57), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1148), .B1(new_n1146), .B2(new_n1157), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1222), .B2(new_n1208), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1209), .B1(new_n1220), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(G375));
  INV_X1    g1025(.A(new_n1157), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n978), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1152), .A2(new_n1148), .A3(new_n1156), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n262), .B1(new_n762), .B2(new_n1097), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n772), .A2(new_n774), .B1(new_n756), .B2(new_n392), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(G107), .C2(new_n814), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n219), .B2(new_n768), .C1(new_n544), .C2(new_n823), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n778), .A2(G303), .B1(G97), .B2(new_n784), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT122), .Z(new_n1235));
  NOR2_X1   g1035(.A1(new_n766), .A2(new_n835), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n834), .A2(new_n762), .B1(new_n765), .B2(new_n749), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1188), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1111), .B2(new_n748), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1015), .B1(G132), .B2(new_n758), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n202), .B2(new_n756), .C1(new_n823), .C2(new_n1107), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1233), .A2(new_n1235), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n742), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n736), .C1(G68), .C2(new_n1096), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n923), .B2(new_n809), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n734), .B(KEYINPUT121), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1229), .A2(new_n1248), .ZN(G381));
  OR2_X1    g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1250), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G378), .A2(new_n1251), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1052(.A(G378), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n679), .A2(G213), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1224), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G407), .A2(G213), .A3(new_n1256), .ZN(G409));
  XNOR2_X1  g1057(.A(G393), .B(new_n807), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1000), .A2(new_n730), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n735), .B1(new_n1260), .B2(new_n1227), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n976), .A2(new_n977), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1028), .B(G390), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G390), .B1(new_n1002), .B2(new_n1028), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1259), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G390), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1260), .A2(new_n1227), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1262), .B1(new_n1268), .B2(new_n734), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1028), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1267), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n1258), .A3(new_n1263), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1266), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1213), .A2(new_n1216), .A3(new_n1247), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1200), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1275), .A2(KEYINPUT124), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n1211), .A2(new_n1212), .B1(new_n1215), .B2(new_n1201), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1219), .A2(new_n1279), .A3(new_n1227), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1275), .A2(KEYINPUT124), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1276), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1253), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT123), .B1(new_n1224), .B2(G378), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1279), .A2(new_n735), .B1(new_n1176), .B2(new_n1199), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1213), .A2(KEYINPUT57), .A3(new_n1216), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n697), .B1(new_n1222), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT57), .B1(new_n1219), .B2(new_n1279), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1285), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT123), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1283), .B1(new_n1284), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  AND2_X1   g1093(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1228), .B1(new_n1157), .B2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1152), .A2(new_n1148), .A3(KEYINPUT60), .A4(new_n1156), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n697), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1248), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1294), .B1(new_n1300), .B2(new_n1248), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1292), .A2(new_n1293), .A3(new_n1254), .A4(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1255), .A2(G2897), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1304), .B(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1311), .A2(KEYINPUT123), .A3(G378), .A4(new_n1285), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1310), .A2(new_n1312), .B1(new_n1253), .B2(new_n1282), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1309), .B1(new_n1313), .B2(new_n1255), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1305), .A2(new_n1306), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1255), .B1(new_n1316), .B2(new_n1283), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1293), .B1(new_n1317), .B2(new_n1304), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1273), .B1(new_n1315), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1304), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1317), .A2(KEYINPUT63), .A3(new_n1304), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1266), .A2(new_n1306), .A3(new_n1272), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(KEYINPUT126), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1322), .A2(new_n1314), .A3(new_n1323), .A4(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1319), .A2(new_n1326), .ZN(G405));
  NAND2_X1  g1127(.A1(G375), .A2(new_n1253), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1273), .A2(new_n1316), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1273), .B1(new_n1316), .B2(new_n1328), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  OR3_X1    g1131(.A1(new_n1302), .A2(KEYINPUT127), .A3(new_n1303), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1331), .B(new_n1333), .ZN(G402));
endmodule


