//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n477), .B2(new_n471), .ZN(new_n478));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  OAI21_X1  g055(.A(G125), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n483), .A2(new_n484), .A3(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n475), .B1(new_n478), .B2(new_n485), .ZN(G160));
  AOI21_X1  g061(.A(new_n471), .B1(new_n464), .B2(new_n465), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(G136), .B2(new_n466), .ZN(G162));
  NAND2_X1  g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n464), .B2(new_n465), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n471), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n466), .B2(G138), .ZN(new_n500));
  OAI211_X1 g075(.A(G138), .B(new_n471), .C1(new_n479), .C2(new_n480), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n506), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n514), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n512), .A2(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(new_n515), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n507), .A2(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n509), .A2(KEYINPUT72), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT72), .B1(new_n509), .B2(new_n528), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n525), .B(new_n527), .C1(new_n529), .C2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n515), .A2(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n518), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n509), .A2(G64), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n511), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n535), .A2(new_n538), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n508), .ZN(new_n541));
  AOI21_X1  g116(.A(G543), .B1(KEYINPUT71), .B2(KEYINPUT5), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n511), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n547), .B1(new_n546), .B2(new_n545), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n526), .A2(G81), .B1(new_n515), .B2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(G91), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT74), .B1(new_n518), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n526), .A2(new_n559), .A3(G91), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n515), .A2(new_n563), .A3(G53), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n558), .A2(new_n560), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n567), .B1(new_n541), .B2(new_n542), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n507), .A2(KEYINPUT76), .A3(new_n508), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT75), .Z(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n565), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(new_n538), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n526), .A2(G90), .B1(new_n515), .B2(G52), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(KEYINPUT77), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n578), .B1(new_n535), .B2(new_n538), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G301));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND2_X1  g157(.A1(new_n526), .A2(G87), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n515), .A2(G49), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  AOI22_X1  g161(.A1(new_n526), .A2(G86), .B1(new_n515), .B2(G48), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT78), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n507), .B2(new_n508), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n543), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n515), .A2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n526), .A2(G85), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n597), .A2(KEYINPUT79), .A3(new_n598), .A4(new_n599), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G301), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n518), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n526), .A2(G92), .A3(new_n607), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n610), .A2(new_n611), .B1(G54), .B2(new_n515), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n568), .B2(new_n569), .ZN(new_n614));
  AND2_X1   g189(.A1(G79), .A2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(G651), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n606), .B1(new_n619), .B2(new_n605), .ZN(G284));
  AOI21_X1  g195(.A(new_n606), .B1(new_n619), .B2(new_n605), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n565), .A2(new_n573), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  OAI21_X1  g202(.A(KEYINPUT82), .B1(new_n551), .B2(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n619), .A2(new_n626), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  MUX2_X1   g205(.A(KEYINPUT82), .B(new_n628), .S(new_n630), .Z(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n473), .A2(new_n476), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n487), .A2(G123), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n466), .A2(G135), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n471), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G2096), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n637), .A2(new_n638), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2443), .B(G2446), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2451), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2454), .Z(new_n659));
  XOR2_X1   g234(.A(new_n655), .B(new_n659), .Z(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G14), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n636), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n644), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n684), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  OAI221_X1 g265(.A(new_n686), .B1(new_n684), .B2(new_n682), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G21), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G168), .B2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(G1966), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G29), .A2(G35), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G162), .B2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n704), .B1(G2090), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT24), .ZN(new_n710));
  INV_X1    g285(.A(G34), .ZN(new_n711));
  AOI21_X1  g286(.A(G29), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n710), .B2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(G160), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(G2084), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n700), .A2(G5), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G171), .B2(new_n700), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1961), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n709), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(G2084), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n708), .A2(G2090), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n714), .A2(G26), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT93), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n487), .A2(G128), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT92), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(G116), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G2105), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G140), .B2(new_n466), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(G29), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2067), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n720), .A2(new_n721), .A3(new_n722), .A4(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n700), .A2(KEYINPUT89), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n700), .A2(KEYINPUT89), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n551), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G19), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n742), .A2(G1341), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(G1341), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  INV_X1    g320(.A(G28), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(KEYINPUT30), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT95), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n643), .B2(new_n714), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n714), .A2(G33), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT25), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(new_n471), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n754), .B(new_n756), .C1(G139), .C2(new_n466), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n752), .B1(new_n757), .B2(new_n714), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(G2072), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n714), .A2(G27), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G164), .B2(new_n714), .ZN(new_n761));
  INV_X1    g336(.A(G2078), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n759), .B(new_n763), .C1(G2072), .C2(new_n758), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n735), .A2(new_n743), .A3(new_n744), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n739), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT97), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G16), .B2(G299), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n714), .A2(G32), .ZN(new_n771));
  AOI22_X1  g346(.A1(G141), .A2(new_n466), .B1(new_n473), .B2(G105), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n487), .A2(G129), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT26), .Z(new_n775));
  NAND3_X1  g350(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n771), .B1(new_n781), .B2(new_n714), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT27), .Z(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G1996), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n770), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  MUX2_X1   g362(.A(G24), .B(G290), .S(new_n738), .Z(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1986), .Z(new_n789));
  MUX2_X1   g364(.A(G6), .B(G305), .S(G16), .Z(new_n790));
  XOR2_X1   g365(.A(KEYINPUT32), .B(G1981), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G23), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT90), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G288), .B2(new_n700), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT33), .B(G1976), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n738), .A2(G22), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n738), .ZN(new_n799));
  INV_X1    g374(.A(G1971), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n792), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n714), .A2(G25), .ZN(new_n805));
  OR2_X1    g380(.A1(G95), .A2(G2105), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n806), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT88), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n487), .A2(G119), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n466), .A2(G131), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n805), .B1(new_n812), .B2(new_n714), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G1991), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n813), .B(new_n814), .Z(new_n815));
  NAND4_X1  g390(.A1(new_n789), .A2(new_n803), .A3(new_n804), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT36), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n700), .A2(G4), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n619), .B2(new_n700), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT91), .B(G1348), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n765), .A2(new_n787), .A3(new_n817), .A4(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  NAND2_X1  g398(.A1(new_n619), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n511), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n515), .A2(G55), .ZN(new_n828));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n518), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n550), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n548), .A2(new_n549), .A3(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n825), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT98), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n832), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(G162), .B(new_n643), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G160), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n494), .B2(new_n497), .ZN(new_n849));
  OAI211_X1 g424(.A(G126), .B(G2105), .C1(new_n479), .C2(new_n480), .ZN(new_n850));
  INV_X1    g425(.A(G114), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT99), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n849), .B(new_n854), .C1(new_n500), .C2(new_n502), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n781), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n780), .A2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n732), .B(KEYINPUT100), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n757), .A2(KEYINPUT101), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n857), .A2(new_n860), .A3(new_n858), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(KEYINPUT101), .A3(new_n757), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n634), .B(new_n812), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n466), .A2(G142), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n487), .A2(G130), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n471), .A2(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n867), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n757), .A2(KEYINPUT101), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n862), .A2(new_n874), .A3(new_n863), .A4(new_n864), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n866), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n873), .B1(new_n866), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n847), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n846), .A3(new_n876), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(new_n832), .A2(new_n605), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n833), .A2(new_n834), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n629), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n617), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n623), .A2(new_n617), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n888), .B2(G299), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(KEYINPUT102), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n623), .A2(new_n898), .A3(new_n617), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n897), .A2(new_n889), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n896), .B1(new_n900), .B2(KEYINPUT41), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n893), .B1(new_n887), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(G305), .ZN(new_n903));
  XNOR2_X1  g478(.A(G166), .B(G288), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT42), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n902), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n885), .B1(new_n907), .B2(new_n605), .ZN(G295));
  OAI21_X1  g483(.A(new_n885), .B1(new_n907), .B2(new_n605), .ZN(G331));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n580), .A2(G168), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n529), .A2(new_n530), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n527), .A2(new_n524), .A3(new_n522), .ZN(new_n915));
  AOI21_X1  g490(.A(G171), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n911), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(G286), .B1(new_n579), .B2(new_n577), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n919), .A2(KEYINPUT103), .A3(new_n916), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n886), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n917), .A3(new_n911), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT103), .B1(new_n919), .B2(new_n916), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n835), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(KEYINPUT104), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n922), .A2(new_n923), .A3(new_n835), .A4(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n892), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n891), .A2(new_n894), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n897), .A2(new_n899), .A3(new_n895), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n921), .A2(new_n924), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n905), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n901), .A2(new_n925), .A3(new_n927), .ZN(new_n933));
  INV_X1    g508(.A(new_n905), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n921), .A2(new_n891), .A3(new_n924), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n882), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT105), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n932), .A2(new_n939), .A3(new_n936), .A4(new_n882), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n910), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n882), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT44), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n942), .B2(new_n943), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(KEYINPUT43), .B2(new_n937), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n950), .ZN(G397));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n855), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n467), .A2(new_n474), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n484), .B1(new_n483), .B2(G2105), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT69), .B(new_n471), .C1(new_n481), .C2(new_n482), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n956), .B(G40), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n780), .B(new_n785), .ZN(new_n961));
  INV_X1    g536(.A(G2067), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n732), .B(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n812), .B(new_n814), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(G290), .B(G1986), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  NOR2_X1   g544(.A1(G288), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n973), .B(G8), .C1(new_n953), .C2(new_n959), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(G160), .A2(G40), .A3(new_n952), .A4(new_n855), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n976), .B2(G8), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n971), .B(new_n972), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1981), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n526), .A2(G86), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n515), .A2(G48), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n592), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT49), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n979), .B1(new_n587), .B2(new_n592), .ZN(new_n987));
  OAI22_X1  g562(.A1(new_n986), .A2(new_n987), .B1(new_n983), .B2(new_n984), .ZN(new_n988));
  INV_X1    g563(.A(new_n987), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n989), .A2(KEYINPUT111), .A3(KEYINPUT49), .A4(new_n982), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n975), .B2(new_n977), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n978), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(G8), .B1(new_n953), .B2(new_n959), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT110), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n970), .B1(new_n995), .B2(new_n974), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT55), .B(G8), .C1(new_n512), .C2(new_n520), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(G166), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT108), .B(new_n1003), .C1(G166), .C2(new_n1004), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n954), .A2(G1384), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n855), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n855), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n503), .A2(new_n952), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n959), .B1(new_n954), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(G1971), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n1020));
  INV_X1    g595(.A(G40), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n1021), .B(new_n475), .C1(new_n478), .C2(new_n485), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n503), .A2(new_n1023), .A3(new_n952), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G2090), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1019), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1010), .B1(new_n1029), .B2(new_n1004), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1009), .A2(KEYINPUT109), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1017), .A2(new_n954), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n855), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1022), .B(new_n1032), .C1(new_n1033), .C2(new_n1013), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n800), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n855), .A2(new_n1023), .A3(new_n952), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n1022), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1035), .B1(G2090), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1002), .A2(new_n1040), .A3(new_n1008), .A4(new_n1007), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1031), .A2(new_n1039), .A3(G8), .A4(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n999), .A2(new_n1030), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1016), .A2(new_n762), .A3(new_n1018), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  INV_X1    g620(.A(G1961), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1044), .A2(new_n1045), .B1(new_n1046), .B2(new_n1038), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n762), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n1048), .B(new_n475), .C1(G2105), .C2(new_n483), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1016), .A2(new_n955), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(G301), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1045), .B1(new_n1034), .B2(G2078), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1012), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n466), .A2(new_n499), .A3(G138), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1053), .B1(new_n1056), .B2(new_n498), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n959), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1058), .A2(new_n955), .A3(KEYINPUT53), .A4(new_n762), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1052), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n580), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT54), .B1(new_n1051), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1043), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(G160), .B(G40), .C1(G164), .C2(new_n1053), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT45), .B1(new_n855), .B2(new_n952), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n703), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT115), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1036), .A2(new_n1022), .A3(new_n1037), .ZN(new_n1069));
  INV_X1    g644(.A(G2084), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(new_n703), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1068), .A2(new_n1071), .A3(G168), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G8), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1966), .B1(new_n1058), .B2(new_n955), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1072), .A2(new_n1076), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1077));
  AOI21_X1  g652(.A(G168), .B1(new_n1077), .B2(new_n1068), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT51), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1074), .A2(new_n1080), .A3(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1052), .A2(new_n1060), .A3(new_n1050), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1084), .B(KEYINPUT54), .C1(new_n580), .C2(new_n1061), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1085), .A2(KEYINPUT125), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(KEYINPUT125), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1064), .B(new_n1082), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1956), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1024), .A2(G40), .A3(G160), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1023), .B1(new_n855), .B2(new_n952), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT56), .B(G2072), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1034), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT118), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1098), .B(new_n1099), .C1(new_n565), .C2(new_n573), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1016), .A2(new_n1018), .A3(new_n1093), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n1092), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1096), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1101), .A3(new_n1092), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1103), .A2(new_n1101), .A3(KEYINPUT122), .A4(new_n1092), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1106), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1108), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1101), .B1(new_n1103), .B2(new_n1092), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT58), .B(G1341), .Z(new_n1118));
  NAND2_X1  g693(.A1(new_n976), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT119), .B(G1996), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1034), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1120), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1018), .B(new_n1124), .C1(new_n1013), .C2(new_n1033), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT120), .A3(new_n1119), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1117), .B1(new_n1127), .B2(new_n551), .ZN(new_n1128));
  AOI211_X1 g703(.A(KEYINPUT59), .B(new_n550), .C1(new_n1123), .C2(new_n1126), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1112), .B(new_n1116), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT123), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1125), .A2(KEYINPUT120), .A3(new_n1119), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT120), .B1(new_n1125), .B2(new_n1119), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n551), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1127), .A2(new_n1117), .A3(new_n551), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n1112), .A4(new_n1116), .ZN(new_n1139));
  INV_X1    g714(.A(G1348), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1038), .A2(new_n1140), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n976), .A2(G2067), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(KEYINPUT124), .ZN(new_n1146));
  INV_X1    g721(.A(new_n619), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1146), .A2(new_n1147), .B1(new_n1144), .B2(new_n1143), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1145), .A2(KEYINPUT124), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n619), .B1(new_n1145), .B2(KEYINPUT124), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1131), .A2(new_n1139), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1143), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1106), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1108), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1088), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  AND4_X1   g731(.A1(G8), .A2(new_n1031), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n993), .A2(new_n998), .A3(KEYINPUT112), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT112), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n995), .A2(new_n974), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n996), .A2(new_n972), .B1(new_n1160), .B2(new_n991), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n975), .A2(new_n977), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT52), .B1(new_n1162), .B2(new_n970), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1159), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1157), .B1(new_n1158), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n992), .ZN(new_n1166));
  OR2_X1    g741(.A1(G288), .A2(G1976), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n982), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1162), .B(KEYINPUT113), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1165), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(G301), .B1(new_n1047), .B2(new_n1059), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n999), .A2(new_n1030), .A3(new_n1042), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1082), .B2(KEYINPUT62), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1079), .A2(new_n1175), .A3(new_n1081), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1171), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1077), .A2(new_n1068), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(G8), .A3(G168), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1178), .B1(new_n1043), .B2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1157), .A2(new_n1180), .A3(new_n1178), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1009), .B1(new_n1039), .B2(G8), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT112), .B1(new_n993), .B2(new_n998), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1161), .A2(new_n1163), .A3(new_n1159), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1182), .B1(new_n1186), .B2(KEYINPUT116), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT116), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n1188), .B(new_n1183), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1181), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1177), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n968), .B1(new_n1156), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n960), .A2(new_n785), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT46), .ZN(new_n1194));
  INV_X1    g769(.A(new_n960), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n963), .A2(new_n781), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT47), .Z(new_n1198));
  OR2_X1    g773(.A1(new_n1198), .A2(KEYINPUT126), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(KEYINPUT126), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n808), .A2(new_n814), .A3(new_n811), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n964), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n727), .A2(new_n962), .A3(new_n731), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1195), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n966), .A2(new_n960), .ZN(new_n1205));
  NOR3_X1   g780(.A1(new_n1195), .A2(G1986), .A3(G290), .ZN(new_n1206));
  XNOR2_X1  g781(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1206), .B(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1204), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  AND3_X1   g784(.A1(new_n1199), .A2(new_n1200), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1192), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g786(.A1(new_n462), .A2(G227), .ZN(new_n1213));
  AND2_X1   g787(.A1(new_n698), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g788(.A(G401), .ZN(new_n1215));
  NAND4_X1  g789(.A1(new_n1214), .A2(new_n1215), .A3(new_n948), .A4(new_n883), .ZN(G225));
  INV_X1    g790(.A(G225), .ZN(G308));
endmodule


