

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U321 ( .A(n346), .B(n328), .ZN(n332) );
  XNOR2_X1 U322 ( .A(n327), .B(KEYINPUT11), .ZN(n328) );
  XNOR2_X1 U323 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U324 ( .A(n367), .B(n340), .ZN(n341) );
  XOR2_X1 U325 ( .A(n353), .B(n352), .Z(n289) );
  INV_X1 U326 ( .A(KEYINPUT25), .ZN(n452) );
  XNOR2_X1 U327 ( .A(n452), .B(KEYINPUT94), .ZN(n453) );
  INV_X1 U328 ( .A(KEYINPUT73), .ZN(n343) );
  XNOR2_X1 U329 ( .A(n454), .B(n453), .ZN(n457) );
  XNOR2_X1 U330 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U331 ( .A(n404), .B(KEYINPUT54), .ZN(n405) );
  XOR2_X1 U332 ( .A(G106GAT), .B(G92GAT), .Z(n326) );
  XNOR2_X1 U333 ( .A(n424), .B(KEYINPUT55), .ZN(n425) );
  XNOR2_X1 U334 ( .A(n388), .B(G36GAT), .ZN(n392) );
  XNOR2_X1 U335 ( .A(n354), .B(n289), .ZN(n355) );
  XNOR2_X1 U336 ( .A(n426), .B(n425), .ZN(n444) );
  XNOR2_X1 U337 ( .A(n392), .B(n412), .ZN(n397) );
  XNOR2_X1 U338 ( .A(n356), .B(n355), .ZN(n360) );
  XNOR2_X1 U339 ( .A(n342), .B(n341), .ZN(n561) );
  XNOR2_X1 U340 ( .A(n403), .B(n402), .ZN(n518) );
  XNOR2_X1 U341 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n475) );
  XNOR2_X1 U342 ( .A(n472), .B(G43GAT), .ZN(n473) );
  XNOR2_X1 U343 ( .A(n476), .B(n475), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n474), .B(n473), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT88), .B(KEYINPUT1), .Z(n291) );
  XNOR2_X1 U346 ( .A(KEYINPUT89), .B(KEYINPUT4), .ZN(n290) );
  XNOR2_X1 U347 ( .A(n291), .B(n290), .ZN(n307) );
  XOR2_X1 U348 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n293) );
  XNOR2_X1 U349 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n292) );
  XNOR2_X1 U350 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U351 ( .A(n294), .B(G85GAT), .Z(n296) );
  XOR2_X1 U352 ( .A(KEYINPUT0), .B(G127GAT), .Z(n432) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(n432), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n301) );
  XOR2_X1 U355 ( .A(G134GAT), .B(G162GAT), .Z(n339) );
  XNOR2_X1 U356 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n297), .B(KEYINPUT2), .ZN(n413) );
  XOR2_X1 U358 ( .A(n339), .B(n413), .Z(n299) );
  NAND2_X1 U359 ( .A1(G225GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U360 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U361 ( .A(n301), .B(n300), .Z(n305) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(G141GAT), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n302), .B(G113GAT), .ZN(n372) );
  XNOR2_X1 U364 ( .A(G120GAT), .B(G57GAT), .ZN(n303) );
  XNOR2_X1 U365 ( .A(n303), .B(G148GAT), .ZN(n358) );
  XNOR2_X1 U366 ( .A(n372), .B(n358), .ZN(n304) );
  XNOR2_X1 U367 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U368 ( .A(n307), .B(n306), .Z(n460) );
  XNOR2_X1 U369 ( .A(KEYINPUT90), .B(n460), .ZN(n516) );
  XOR2_X1 U370 ( .A(G64GAT), .B(G211GAT), .Z(n309) );
  XNOR2_X1 U371 ( .A(G8GAT), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U372 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U373 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n311) );
  XNOR2_X1 U374 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n310) );
  XNOR2_X1 U375 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U376 ( .A(n313), .B(n312), .ZN(n324) );
  XOR2_X1 U377 ( .A(G22GAT), .B(G15GAT), .Z(n370) );
  XOR2_X1 U378 ( .A(G155GAT), .B(G57GAT), .Z(n315) );
  XNOR2_X1 U379 ( .A(G1GAT), .B(G127GAT), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U381 ( .A(n370), .B(n316), .Z(n318) );
  NAND2_X1 U382 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U384 ( .A(n319), .B(KEYINPUT81), .Z(n322) );
  XNOR2_X1 U385 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n320) );
  XNOR2_X1 U386 ( .A(n320), .B(G78GAT), .ZN(n357) );
  XNOR2_X1 U387 ( .A(n357), .B(KEYINPUT14), .ZN(n321) );
  XNOR2_X1 U388 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U389 ( .A(n324), .B(n323), .Z(n577) );
  INV_X1 U390 ( .A(n577), .ZN(n557) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .ZN(n325) );
  XNOR2_X1 U392 ( .A(n326), .B(n325), .ZN(n346) );
  AND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  XOR2_X1 U394 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n330) );
  XNOR2_X1 U395 ( .A(KEYINPUT77), .B(KEYINPUT76), .ZN(n329) );
  XNOR2_X1 U396 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U397 ( .A(n332), .B(n331), .Z(n342) );
  XOR2_X1 U398 ( .A(G29GAT), .B(G36GAT), .Z(n334) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(G43GAT), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U401 ( .A(KEYINPUT7), .B(KEYINPUT70), .Z(n336) );
  XNOR2_X1 U402 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U404 ( .A(n338), .B(n337), .Z(n367) );
  XOR2_X1 U405 ( .A(G190GAT), .B(G218GAT), .Z(n393) );
  XNOR2_X1 U406 ( .A(n339), .B(n393), .ZN(n340) );
  NAND2_X1 U407 ( .A1(n557), .A2(n561), .ZN(n377) );
  NAND2_X1 U408 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  NAND2_X1 U409 ( .A1(n347), .A2(KEYINPUT31), .ZN(n351) );
  INV_X1 U410 ( .A(n347), .ZN(n349) );
  INV_X1 U411 ( .A(KEYINPUT31), .ZN(n348) );
  NAND2_X1 U412 ( .A1(n349), .A2(n348), .ZN(n350) );
  NAND2_X1 U413 ( .A1(n351), .A2(n350), .ZN(n356) );
  XOR2_X1 U414 ( .A(G176GAT), .B(G64GAT), .Z(n387) );
  XOR2_X1 U415 ( .A(G204GAT), .B(n387), .Z(n354) );
  XOR2_X1 U416 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n353) );
  XNOR2_X1 U417 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n573) );
  XNOR2_X1 U420 ( .A(n573), .B(KEYINPUT41), .ZN(n552) );
  XOR2_X1 U421 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n362) );
  NAND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U424 ( .A(n363), .B(KEYINPUT66), .Z(n369) );
  XOR2_X1 U425 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n365) );
  XNOR2_X1 U426 ( .A(G197GAT), .B(KEYINPUT67), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U429 ( .A(n369), .B(n368), .ZN(n371) );
  XOR2_X1 U430 ( .A(n371), .B(n370), .Z(n374) );
  XOR2_X1 U431 ( .A(G169GAT), .B(G8GAT), .Z(n401) );
  XNOR2_X1 U432 ( .A(n372), .B(n401), .ZN(n373) );
  XNOR2_X1 U433 ( .A(n374), .B(n373), .ZN(n569) );
  NOR2_X1 U434 ( .A1(n552), .A2(n569), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n375), .B(KEYINPUT46), .ZN(n376) );
  NOR2_X1 U436 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n378), .B(KEYINPUT47), .ZN(n385) );
  INV_X1 U438 ( .A(KEYINPUT36), .ZN(n380) );
  INV_X1 U439 ( .A(KEYINPUT78), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n379), .B(n561), .ZN(n542) );
  XNOR2_X1 U441 ( .A(n380), .B(n542), .ZN(n449) );
  NOR2_X1 U442 ( .A1(n557), .A2(n449), .ZN(n381) );
  XOR2_X1 U443 ( .A(KEYINPUT45), .B(n381), .Z(n382) );
  NOR2_X1 U444 ( .A1(n573), .A2(n382), .ZN(n383) );
  XNOR2_X1 U445 ( .A(n569), .B(KEYINPUT72), .ZN(n531) );
  NAND2_X1 U446 ( .A1(n383), .A2(n531), .ZN(n384) );
  NAND2_X1 U447 ( .A1(n385), .A2(n384), .ZN(n386) );
  XNOR2_X1 U448 ( .A(KEYINPUT48), .B(n386), .ZN(n527) );
  XOR2_X1 U449 ( .A(n387), .B(G92GAT), .Z(n388) );
  XOR2_X1 U450 ( .A(KEYINPUT85), .B(G211GAT), .Z(n390) );
  XNOR2_X1 U451 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U453 ( .A(G197GAT), .B(n391), .Z(n412) );
  XOR2_X1 U454 ( .A(KEYINPUT91), .B(n393), .Z(n395) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U457 ( .A(n397), .B(n396), .Z(n403) );
  XOR2_X1 U458 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n399) );
  XNOR2_X1 U459 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U461 ( .A(KEYINPUT19), .B(n400), .Z(n439) );
  XNOR2_X1 U462 ( .A(n401), .B(n439), .ZN(n402) );
  NAND2_X1 U463 ( .A1(n527), .A2(n518), .ZN(n406) );
  XOR2_X1 U464 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n404) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n407) );
  NOR2_X1 U466 ( .A1(n516), .A2(n407), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n408), .B(KEYINPUT64), .ZN(n568) );
  XOR2_X1 U468 ( .A(G78GAT), .B(G148GAT), .Z(n410) );
  XNOR2_X1 U469 ( .A(G141GAT), .B(G22GAT), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n423) );
  XOR2_X1 U472 ( .A(G106GAT), .B(G218GAT), .Z(n415) );
  XNOR2_X1 U473 ( .A(G50GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U475 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n417) );
  NAND2_X1 U476 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U478 ( .A(n419), .B(n418), .Z(n421) );
  XNOR2_X1 U479 ( .A(G162GAT), .B(KEYINPUT22), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n461) );
  NAND2_X1 U482 ( .A1(n568), .A2(n461), .ZN(n426) );
  XOR2_X1 U483 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n424) );
  XOR2_X1 U484 ( .A(G71GAT), .B(G176GAT), .Z(n428) );
  XNOR2_X1 U485 ( .A(G169GAT), .B(G15GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n443) );
  XOR2_X1 U487 ( .A(G120GAT), .B(G99GAT), .Z(n430) );
  XNOR2_X1 U488 ( .A(G113GAT), .B(G190GAT), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U490 ( .A(n431), .B(G134GAT), .Z(n434) );
  XNOR2_X1 U491 ( .A(G43GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U493 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n436) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U496 ( .A(n438), .B(n437), .Z(n441) );
  XNOR2_X1 U497 ( .A(n439), .B(KEYINPUT83), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U499 ( .A(n443), .B(n442), .Z(n530) );
  INV_X1 U500 ( .A(n530), .ZN(n520) );
  NAND2_X1 U501 ( .A1(n444), .A2(n520), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n445), .B(KEYINPUT125), .ZN(n565) );
  INV_X1 U503 ( .A(n552), .ZN(n534) );
  NAND2_X1 U504 ( .A1(n565), .A2(n534), .ZN(n448) );
  XOR2_X1 U505 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n446) );
  XNOR2_X1 U506 ( .A(n446), .B(G176GAT), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(G1349GAT) );
  XOR2_X1 U508 ( .A(KEYINPUT38), .B(KEYINPUT102), .Z(n471) );
  NOR2_X1 U509 ( .A1(n573), .A2(n531), .ZN(n480) );
  NAND2_X1 U510 ( .A1(n518), .A2(n520), .ZN(n450) );
  XOR2_X1 U511 ( .A(KEYINPUT93), .B(n450), .Z(n451) );
  NAND2_X1 U512 ( .A1(n451), .A2(n461), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n518), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U514 ( .A1(n520), .A2(n461), .ZN(n455) );
  XOR2_X1 U515 ( .A(n455), .B(KEYINPUT26), .Z(n547) );
  INV_X1 U516 ( .A(n547), .ZN(n567) );
  NAND2_X1 U517 ( .A1(n463), .A2(n567), .ZN(n456) );
  NAND2_X1 U518 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U519 ( .A(KEYINPUT95), .B(n458), .ZN(n459) );
  NOR2_X1 U520 ( .A1(n460), .A2(n459), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n461), .B(KEYINPUT65), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT28), .ZN(n523) );
  NAND2_X1 U523 ( .A1(n516), .A2(n463), .ZN(n546) );
  NOR2_X1 U524 ( .A1(n523), .A2(n546), .ZN(n528) );
  XOR2_X1 U525 ( .A(n528), .B(KEYINPUT92), .Z(n464) );
  NOR2_X1 U526 ( .A1(n520), .A2(n464), .ZN(n465) );
  NOR2_X1 U527 ( .A1(n466), .A2(n465), .ZN(n479) );
  NOR2_X1 U528 ( .A1(n449), .A2(n479), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n557), .A2(n467), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT101), .B(n468), .ZN(n469) );
  XOR2_X1 U531 ( .A(KEYINPUT37), .B(n469), .Z(n513) );
  NAND2_X1 U532 ( .A1(n480), .A2(n513), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n471), .B(n470), .ZN(n498) );
  NAND2_X1 U534 ( .A1(n498), .A2(n520), .ZN(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n472) );
  NAND2_X1 U536 ( .A1(n542), .A2(n565), .ZN(n476) );
  NOR2_X1 U537 ( .A1(n557), .A2(n542), .ZN(n477) );
  XOR2_X1 U538 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  NOR2_X1 U539 ( .A1(n479), .A2(n478), .ZN(n501) );
  AND2_X1 U540 ( .A1(n480), .A2(n501), .ZN(n489) );
  NAND2_X1 U541 ( .A1(n516), .A2(n489), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(KEYINPUT34), .ZN(n482) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U544 ( .A1(n489), .A2(n518), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n483), .B(KEYINPUT96), .ZN(n484) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(n484), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n486) );
  NAND2_X1 U548 ( .A1(n489), .A2(n520), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(n488) );
  XOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT97), .Z(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  XOR2_X1 U552 ( .A(G22GAT), .B(KEYINPUT99), .Z(n491) );
  NAND2_X1 U553 ( .A1(n489), .A2(n523), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT100), .B(KEYINPUT103), .Z(n493) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(n495) );
  NAND2_X1 U558 ( .A1(n516), .A2(n498), .ZN(n494) );
  XOR2_X1 U559 ( .A(n495), .B(n494), .Z(G1328GAT) );
  NAND2_X1 U560 ( .A1(n498), .A2(n518), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n496), .B(KEYINPUT104), .ZN(n497) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n498), .A2(n523), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U565 ( .A1(n534), .A2(n569), .ZN(n500) );
  XOR2_X1 U566 ( .A(KEYINPUT106), .B(n500), .Z(n514) );
  AND2_X1 U567 ( .A1(n501), .A2(n514), .ZN(n508) );
  NAND2_X1 U568 ( .A1(n508), .A2(n516), .ZN(n502) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n502), .ZN(n503) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n505) );
  NAND2_X1 U572 ( .A1(n508), .A2(n518), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U574 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n520), .A2(n508), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U578 ( .A1(n508), .A2(n523), .ZN(n509) );
  XNOR2_X1 U579 ( .A(n510), .B(n509), .ZN(n512) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT110), .Z(n511) );
  XNOR2_X1 U581 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(KEYINPUT111), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n516), .A2(n524), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n517), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n524), .A2(n518), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n520), .A2(n524), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n521), .B(KEYINPUT112), .ZN(n522) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n522), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT113), .Z(n533) );
  NAND2_X1 U595 ( .A1(n527), .A2(n528), .ZN(n529) );
  NOR2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n543) );
  INV_X1 U597 ( .A(n531), .ZN(n563) );
  NAND2_X1 U598 ( .A1(n543), .A2(n563), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n536) );
  NAND2_X1 U601 ( .A1(n543), .A2(n534), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT114), .Z(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n540) );
  NAND2_X1 U606 ( .A1(n543), .A2(n577), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n527), .A2(n548), .ZN(n560) );
  NOR2_X1 U614 ( .A1(n569), .A2(n560), .ZN(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  NOR2_X1 U618 ( .A1(n560), .A2(n552), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n560), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(n558), .Z(n559) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NAND2_X1 U628 ( .A1(n565), .A2(n563), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n577), .A2(n565), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n581) );
  NOR2_X1 U633 ( .A1(n569), .A2(n581), .ZN(n571) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  INV_X1 U638 ( .A(n581), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n576), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n449), .A2(n581), .ZN(n582) );
  XOR2_X1 U647 ( .A(n583), .B(n582), .Z(G1355GAT) );
endmodule

