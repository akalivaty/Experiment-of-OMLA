//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT29), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n205));
  INV_X1    g004(.A(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT73), .A2(G197gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(KEYINPUT73), .A2(G197gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n211));
  INV_X1    g010(.A(G197gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(G204gat), .A3(new_n207), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n205), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G211gat), .B(G218gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n204), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  AOI211_X1 g017(.A(new_n205), .B(new_n216), .C1(new_n210), .C2(new_n214), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n203), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G141gat), .B(G148gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(KEYINPUT2), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G148gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT78), .B(G141gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G148gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n221), .B1(new_n230), .B2(new_n222), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n225), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n220), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n216), .A2(KEYINPUT74), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n215), .B(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n203), .B(new_n225), .C1(new_n229), .C2(new_n231), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n204), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G228gat), .A2(G233gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT86), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n210), .A2(new_n214), .ZN(new_n243));
  INV_X1    g042(.A(new_n205), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n234), .ZN(new_n246));
  INV_X1    g045(.A(new_n234), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n215), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT29), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n232), .B1(new_n249), .B2(KEYINPUT3), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n240), .B1(new_n235), .B2(new_n237), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G22gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n242), .A2(new_n252), .A3(KEYINPUT87), .A4(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G78gat), .B(G106gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G50gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n250), .A2(new_n251), .ZN(new_n260));
  INV_X1    g059(.A(new_n241), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n261), .B1(new_n233), .B2(new_n238), .ZN(new_n262));
  OAI21_X1  g061(.A(G22gat), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT87), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n252), .A3(new_n253), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT88), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n239), .A2(new_n241), .B1(new_n250), .B2(new_n251), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n258), .B1(new_n270), .B2(new_n253), .ZN(new_n271));
  OAI211_X1 g070(.A(KEYINPUT88), .B(G22gat), .C1(new_n260), .C2(new_n262), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n267), .A2(new_n273), .A3(KEYINPUT89), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT89), .B1(new_n267), .B2(new_n273), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT23), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(G169gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n279));
  INV_X1    g078(.A(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT65), .ZN(new_n284));
  OR2_X1    g083(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(G190gat), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n277), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n278), .A2(new_n281), .A3(new_n293), .A4(new_n282), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n284), .A2(new_n287), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND4_X1   g096(.A1(new_n287), .A2(new_n288), .A3(new_n290), .A4(new_n291), .ZN(new_n298));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n296), .B1(new_n299), .B2(KEYINPUT23), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(KEYINPUT26), .ZN(new_n303));
  INV_X1    g102(.A(G183gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n304), .B2(new_n289), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT26), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(new_n299), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(new_n289), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n312), .B2(new_n289), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n316));
  OAI22_X1  g115(.A1(KEYINPUT67), .A2(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n304), .A2(KEYINPUT27), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G183gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n320), .A3(new_n289), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n316), .B1(new_n321), .B2(KEYINPUT67), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT67), .B1(new_n321), .B2(KEYINPUT66), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n310), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n322), .A2(new_n323), .ZN(new_n327));
  AOI211_X1 g126(.A(KEYINPUT67), .B(new_n316), .C1(new_n321), .C2(KEYINPUT66), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n309), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n302), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G134gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G127gat), .ZN(new_n334));
  INV_X1    g133(.A(G127gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G134gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n337), .B1(new_n338), .B2(KEYINPUT1), .ZN(new_n339));
  INV_X1    g138(.A(G120gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G113gat), .ZN(new_n341));
  INV_X1    g140(.A(G113gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n295), .A2(new_n296), .B1(new_n298), .B2(new_n300), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n329), .A2(new_n330), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n339), .A2(new_n347), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n349), .A2(new_n350), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT72), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT34), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI211_X1 g160(.A(KEYINPUT72), .B(KEYINPUT34), .C1(new_n357), .C2(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(KEYINPUT72), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n350), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n354), .A2(new_n355), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n348), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n370));
  XNOR2_X1  g169(.A(G15gat), .B(G43gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n369), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n370), .B(new_n374), .C1(new_n375), .C2(KEYINPUT33), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n349), .A2(new_n356), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(new_n366), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n373), .A2(KEYINPUT69), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n373), .A2(KEYINPUT69), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(KEYINPUT33), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT70), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n369), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n382), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n376), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n369), .A2(KEYINPUT32), .A3(new_n382), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT70), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n384), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n359), .A2(new_n360), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n363), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n391), .B(new_n376), .C1(new_n393), .C2(new_n361), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n276), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n396));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n302), .A2(new_n329), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n204), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n399), .B(new_n235), .C1(new_n354), .C2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  AOI21_X1  g203(.A(KEYINPUT29), .B1(new_n302), .B2(new_n329), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n405), .A2(new_n406), .A3(new_n398), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n204), .B1(new_n325), .B2(new_n351), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT75), .B1(new_n408), .B2(new_n397), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n246), .A2(new_n248), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n354), .B2(new_n397), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n401), .B(new_n404), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n401), .B1(new_n410), .B2(new_n412), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT76), .B(new_n401), .C1(new_n410), .C2(new_n412), .ZN(new_n419));
  INV_X1    g218(.A(new_n404), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT77), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT77), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n418), .A2(new_n423), .A3(new_n419), .A4(new_n420), .ZN(new_n424));
  AOI211_X1 g223(.A(new_n396), .B(new_n415), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n424), .ZN(new_n426));
  INV_X1    g225(.A(new_n415), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT90), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n202), .B(new_n395), .C1(new_n425), .C2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430));
  XOR2_X1   g229(.A(G1gat), .B(G29gat), .Z(new_n431));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n232), .A2(new_n348), .A3(KEYINPUT79), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n226), .A2(KEYINPUT78), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT78), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G141gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n441), .A3(G148gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n227), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n222), .A2(new_n230), .ZN(new_n445));
  INV_X1    g244(.A(G155gat), .ZN(new_n446));
  INV_X1    g245(.A(G162gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(G148gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(G141gat), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n230), .B1(new_n227), .B2(new_n450), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n444), .A2(new_n448), .B1(new_n451), .B2(new_n223), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n438), .B1(new_n355), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT4), .B1(new_n437), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n232), .A2(new_n348), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(KEYINPUT4), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT81), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT4), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT79), .B1(new_n232), .B2(new_n348), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n355), .A2(new_n452), .A3(new_n438), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT81), .B1(new_n463), .B2(new_n456), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n348), .A3(new_n236), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g266(.A1(G225gat), .A2(G233gat), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n459), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT82), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n459), .A2(new_n464), .A3(new_n469), .A4(KEYINPUT82), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n461), .B(new_n462), .C1(new_n452), .C2(new_n355), .ZN(new_n475));
  INV_X1    g274(.A(new_n468), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n467), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(new_n460), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n455), .A2(KEYINPUT4), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n468), .A4(new_n466), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n436), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n430), .B1(new_n482), .B2(KEYINPUT6), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n481), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n472), .B2(new_n473), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n487));
  NOR4_X1   g286(.A1(new_n486), .A2(KEYINPUT83), .A3(new_n487), .A4(new_n436), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(KEYINPUT94), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(new_n483), .B2(new_n488), .ZN(new_n492));
  INV_X1    g291(.A(new_n482), .ZN(new_n493));
  AOI211_X1 g292(.A(new_n435), .B(new_n485), .C1(new_n472), .C2(new_n473), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n495), .A3(new_n487), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n487), .B1(new_n486), .B2(new_n436), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(new_n494), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT93), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n490), .A2(new_n492), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT95), .B1(new_n429), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n426), .A2(new_n427), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n500), .A2(new_n483), .A3(new_n488), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT84), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n484), .A2(new_n496), .A3(new_n489), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n415), .B1(new_n422), .B2(new_n424), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT84), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n510), .A3(new_n395), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n512));
  INV_X1    g311(.A(new_n428), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(KEYINPUT90), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI211_X1 g314(.A(KEYINPUT35), .B(new_n276), .C1(new_n394), .C2(new_n387), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n490), .A2(new_n492), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n501), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT95), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n515), .A2(new_n516), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n512), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n387), .A2(new_n394), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n387), .A2(new_n394), .A3(KEYINPUT36), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n506), .A2(new_n510), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n528), .B2(new_n276), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n459), .A2(new_n464), .A3(new_n466), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n530), .A2(KEYINPUT91), .A3(new_n476), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT91), .B1(new_n530), .B2(new_n476), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(KEYINPUT39), .C1(new_n476), .C2(new_n475), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT39), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n531), .B2(new_n532), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n536), .A2(new_n537), .A3(new_n436), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n536), .B2(new_n436), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n534), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT40), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n482), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g341(.A(KEYINPUT40), .B(new_n534), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n513), .A2(new_n542), .A3(new_n543), .A4(new_n514), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT38), .ZN(new_n545));
  AOI211_X1 g344(.A(new_n411), .B(new_n410), .C1(new_n332), .C2(new_n398), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n399), .B1(new_n354), .B2(new_n400), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT37), .B1(new_n547), .B2(new_n235), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n545), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n420), .B1(new_n416), .B2(KEYINPUT37), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n413), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n418), .A2(KEYINPUT37), .A3(new_n419), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n552), .B(new_n420), .C1(KEYINPUT37), .C2(new_n416), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n551), .B1(new_n553), .B2(KEYINPUT38), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n502), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n276), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n544), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n529), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n522), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G29gat), .A2(G36gat), .ZN(new_n560));
  OR3_X1    g359(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT97), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n563));
  NOR3_X1   g362(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT97), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n560), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G50gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G43gat), .ZN(new_n569));
  INV_X1    g368(.A(G43gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G50gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT96), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(new_n571), .A3(KEYINPUT96), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n567), .A2(KEYINPUT15), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n560), .B(KEYINPUT99), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n577), .B1(new_n561), .B2(new_n563), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT15), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n571), .A2(KEYINPUT98), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(new_n569), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n571), .A2(KEYINPUT98), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n574), .A2(KEYINPUT15), .A3(new_n575), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n578), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n576), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT17), .ZN(new_n587));
  NAND2_X1  g386(.A1(G85gat), .A2(G92gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT7), .ZN(new_n589));
  NOR2_X1   g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(KEYINPUT8), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G99gat), .B(G106gat), .Z(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT103), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n593), .A2(new_n594), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT104), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n596), .B(new_n597), .Z(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n602), .A2(new_n586), .B1(KEYINPUT41), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G190gat), .B(G218gat), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n606), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n601), .A2(new_n608), .A3(new_n604), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n607), .A2(new_n613), .A3(new_n609), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G57gat), .B(G64gat), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n618), .A2(KEYINPUT101), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G71gat), .B(G78gat), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G127gat), .ZN(new_n630));
  XOR2_X1   g429(.A(G183gat), .B(G211gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G15gat), .B(G22gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT16), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(G1gat), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(G1gat), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G8gat), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n626), .B2(new_n625), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT102), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(new_n446), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n632), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n617), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n602), .A2(new_n625), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n597), .A2(KEYINPUT105), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n647), .A2(new_n595), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n595), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n623), .B(new_n624), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n623), .A4(new_n624), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n646), .A2(new_n650), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT106), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n661), .B(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n637), .A2(new_n586), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n587), .B2(new_n638), .ZN(new_n667));
  NAND2_X1  g466(.A1(G229gat), .A2(G233gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT18), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(KEYINPUT100), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n637), .B(new_n586), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n668), .B(KEYINPUT13), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(KEYINPUT100), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n667), .A2(new_n668), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n671), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G113gat), .B(G141gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G197gat), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT11), .B(G169gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT12), .Z(new_n682));
  OR2_X1    g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n645), .A2(new_n665), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n559), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n507), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(G1gat), .Z(G1324gat));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n688), .A2(new_n515), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT16), .B(G8gat), .Z(new_n693));
  AOI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G8gat), .B1(new_n688), .B2(new_n515), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n696));
  MUX2_X1   g495(.A(KEYINPUT107), .B(new_n696), .S(new_n693), .Z(new_n697));
  AOI22_X1  g496(.A1(new_n694), .A2(new_n695), .B1(new_n692), .B2(new_n697), .ZN(G1325gat));
  INV_X1    g497(.A(new_n527), .ZN(new_n699));
  OAI21_X1  g498(.A(G15gat), .B1(new_n688), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n523), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(G15gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n688), .B2(new_n702), .ZN(G1326gat));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n556), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  AOI21_X1  g505(.A(new_n617), .B1(new_n522), .B2(new_n558), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n665), .A2(new_n686), .A3(new_n644), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G29gat), .A3(new_n507), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT45), .Z(new_n711));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n617), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n615), .A2(KEYINPUT108), .A3(new_n616), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n559), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n707), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n708), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n507), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n711), .A2(new_n721), .ZN(G1328gat));
  NOR3_X1   g521(.A1(new_n709), .A2(G36gat), .A3(new_n515), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n720), .B2(new_n515), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1329gat));
  OAI21_X1  g526(.A(new_n570), .B1(new_n709), .B2(new_n701), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n527), .A2(G43gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n720), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n556), .A2(new_n568), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n719), .A2(new_n708), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n556), .B1(new_n709), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n707), .A2(KEYINPUT110), .A3(new_n708), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n732), .B(new_n734), .C1(new_n738), .C2(G50gat), .ZN(new_n739));
  AOI21_X1  g538(.A(G50gat), .B1(new_n736), .B2(new_n737), .ZN(new_n740));
  INV_X1    g539(.A(new_n734), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT48), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(G1331gat));
  NAND2_X1  g542(.A1(new_n665), .A2(new_n686), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n645), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n559), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n505), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g548(.A1(new_n746), .A2(new_n515), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  AND2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n752), .B2(new_n755), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(G1333gat));
  OR3_X1    g558(.A1(new_n746), .A2(G71gat), .A3(new_n701), .ZN(new_n760));
  OAI21_X1  g559(.A(G71gat), .B1(new_n746), .B2(new_n699), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n276), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n744), .A2(new_n644), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT112), .Z(new_n767));
  INV_X1    g566(.A(new_n617), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n718), .B1(new_n559), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n716), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n522), .B2(new_n558), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n505), .B(new_n767), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G85gat), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT51), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n644), .A2(new_n685), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n774), .A2(KEYINPUT51), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n707), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n665), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n779), .A2(G85gat), .A3(new_n507), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n559), .A2(new_n768), .A3(new_n776), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n778), .B(new_n780), .C1(new_n781), .C2(new_n775), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n773), .A2(KEYINPUT114), .A3(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(new_n515), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n788), .B(new_n767), .C1(new_n769), .C2(new_n771), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G92gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n515), .A2(G92gat), .A3(new_n779), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n778), .B(new_n791), .C1(new_n781), .C2(new_n775), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n790), .B2(new_n792), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(G1337gat));
  NAND3_X1  g595(.A1(new_n719), .A2(new_n527), .A3(new_n767), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G99gat), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n779), .A2(new_n701), .A3(G99gat), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n778), .B(new_n799), .C1(new_n781), .C2(new_n775), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1338gat));
  OAI211_X1 g600(.A(new_n276), .B(new_n767), .C1(new_n769), .C2(new_n771), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n719), .A2(KEYINPUT117), .A3(new_n276), .A4(new_n767), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(G106gat), .A3(new_n805), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n779), .A2(G106gat), .A3(new_n556), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT116), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n778), .B(new_n808), .C1(new_n781), .C2(new_n775), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n802), .A2(G106gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n809), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(G1339gat));
  INV_X1    g615(.A(new_n644), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n653), .A2(new_n658), .A3(new_n654), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n657), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n658), .B1(new_n653), .B2(new_n654), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n664), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n657), .A2(new_n659), .A3(new_n664), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n667), .A2(new_n668), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n672), .A2(new_n673), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n681), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n683), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n819), .A2(new_n822), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI211_X1 g632(.A(KEYINPUT118), .B(KEYINPUT55), .C1(new_n819), .C2(new_n822), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n825), .B(new_n829), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n715), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n825), .B(new_n685), .C1(new_n833), .C2(new_n834), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n665), .A2(new_n829), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n837), .A2(new_n838), .B1(new_n713), .B2(new_n714), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n817), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n645), .A2(new_n665), .A3(new_n685), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n276), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(new_n505), .A3(new_n515), .A4(new_n523), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n686), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(new_n342), .ZN(G1340gat));
  OAI21_X1  g646(.A(G120gat), .B1(new_n845), .B2(new_n779), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n665), .A2(new_n340), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT119), .Z(new_n850));
  OAI21_X1  g649(.A(new_n848), .B1(new_n845), .B2(new_n850), .ZN(G1341gat));
  NOR2_X1   g650(.A1(new_n845), .A2(new_n817), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(new_n335), .ZN(G1342gat));
  NOR2_X1   g652(.A1(new_n788), .A2(new_n617), .ZN(new_n854));
  AOI211_X1 g653(.A(new_n507), .B(new_n701), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n844), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n856), .B(new_n857), .Z(G1343gat));
  INV_X1    g657(.A(new_n228), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n788), .A2(new_n507), .A3(new_n527), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n842), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n861), .B2(new_n276), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n556), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n831), .A2(new_n832), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n825), .A2(new_n685), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n768), .B1(new_n838), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n817), .B1(new_n836), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n869), .B2(new_n842), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n860), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n859), .B1(new_n871), .B2(new_n686), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT120), .B1(new_n843), .B2(new_n507), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n527), .A2(new_n556), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n507), .B1(new_n840), .B2(new_n842), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n685), .A2(new_n226), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT121), .Z(new_n880));
  NAND4_X1  g679(.A1(new_n873), .A2(new_n878), .A3(new_n515), .A4(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n872), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n872), .B2(new_n881), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(G1344gat));
  INV_X1    g684(.A(new_n860), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n863), .B1(new_n843), .B2(new_n556), .ZN(new_n887));
  INV_X1    g686(.A(new_n870), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n665), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n835), .A2(new_n617), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n817), .B1(new_n868), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n842), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n276), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n865), .B1(new_n840), .B2(new_n842), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n665), .A3(new_n860), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n873), .A2(new_n878), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n788), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n890), .B1(new_n901), .B2(new_n665), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n891), .B(new_n899), .C1(new_n902), .C2(G148gat), .ZN(G1345gat));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n446), .A3(new_n644), .ZN(new_n904));
  OAI21_X1  g703(.A(G155gat), .B1(new_n871), .B2(new_n817), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  INV_X1    g706(.A(new_n715), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n447), .B1(new_n889), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n854), .A2(new_n447), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n900), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n907), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G162gat), .B1(new_n871), .B2(new_n715), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n913), .B(KEYINPUT123), .C1(new_n900), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1347gat));
  NAND2_X1  g714(.A1(new_n788), .A2(new_n507), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(new_n276), .A3(new_n701), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n861), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(G169gat), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n918), .A2(new_n919), .A3(new_n686), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n861), .A2(new_n507), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n515), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n861), .A2(KEYINPUT124), .A3(new_n507), .ZN(new_n924));
  AND3_X1   g723(.A1(new_n923), .A2(new_n395), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n685), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n920), .B1(new_n926), .B2(new_n919), .ZN(G1348gat));
  AOI21_X1  g726(.A(G176gat), .B1(new_n925), .B2(new_n665), .ZN(new_n928));
  INV_X1    g727(.A(new_n918), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n779), .B1(new_n281), .B2(new_n282), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(G1349gat));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n929), .A2(new_n932), .A3(new_n644), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT125), .B1(new_n918), .B2(new_n817), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(G183gat), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n644), .A2(new_n312), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n923), .A2(new_n395), .A3(new_n924), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n937), .A3(KEYINPUT126), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT60), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n935), .A2(new_n937), .A3(KEYINPUT126), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n289), .A3(new_n908), .ZN(new_n943));
  OAI21_X1  g742(.A(G190gat), .B1(new_n918), .B2(new_n617), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1351gat));
  AND2_X1   g745(.A1(new_n923), .A2(new_n924), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n685), .A3(new_n874), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n916), .A2(new_n527), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n897), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n686), .A2(new_n212), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n948), .A2(new_n212), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  NAND3_X1  g751(.A1(new_n923), .A2(new_n874), .A3(new_n924), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n665), .A2(new_n206), .ZN(new_n954));
  OR3_X1    g753(.A1(new_n953), .A2(KEYINPUT62), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n897), .A2(new_n665), .A3(new_n949), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G204gat), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT62), .B1(new_n953), .B2(new_n954), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(G1353gat));
  NOR2_X1   g758(.A1(new_n817), .A2(G211gat), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n947), .A2(KEYINPUT127), .A3(new_n874), .A4(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962));
  INV_X1    g761(.A(new_n960), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n953), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n644), .B(new_n949), .C1(new_n895), .C2(new_n896), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G211gat), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n965), .A2(new_n969), .ZN(G1354gat));
  INV_X1    g769(.A(G218gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n971), .B1(new_n950), .B2(new_n768), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n953), .A2(G218gat), .A3(new_n715), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n972), .A2(new_n973), .ZN(G1355gat));
endmodule


