

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n702, n703, n704, n705, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799;

  INV_X1 U369 ( .A(n678), .ZN(n347) );
  INV_X1 U370 ( .A(KEYINPUT60), .ZN(n349) );
  INV_X1 U371 ( .A(KEYINPUT56), .ZN(n351) );
  NOR2_X1 U372 ( .A1(n626), .A2(n624), .ZN(n519) );
  XNOR2_X1 U373 ( .A(G137), .B(G128), .ZN(n505) );
  XNOR2_X1 U374 ( .A(n464), .B(KEYINPUT33), .ZN(n731) );
  NAND2_X1 U375 ( .A1(n731), .A2(n552), .ZN(n463) );
  XOR2_X2 U376 ( .A(n695), .B(n694), .Z(n696) );
  NAND2_X2 U377 ( .A1(n643), .A2(n724), .ZN(n543) );
  XNOR2_X2 U378 ( .A(n472), .B(n541), .ZN(n643) );
  XNOR2_X1 U379 ( .A(n348), .B(n347), .ZN(G57) );
  NAND2_X1 U380 ( .A1(n357), .A2(n354), .ZN(n348) );
  XNOR2_X1 U381 ( .A(n350), .B(n349), .ZN(G60) );
  NAND2_X1 U382 ( .A1(n355), .A2(n354), .ZN(n350) );
  XNOR2_X1 U383 ( .A(n352), .B(n351), .ZN(G51) );
  NAND2_X1 U384 ( .A1(n359), .A2(n354), .ZN(n352) );
  XNOR2_X1 U385 ( .A(G131), .B(G101), .ZN(n525) );
  XNOR2_X1 U386 ( .A(G113), .B(G143), .ZN(n556) );
  INV_X1 U387 ( .A(G953), .ZN(n780) );
  XOR2_X1 U388 ( .A(G122), .B(KEYINPUT125), .Z(n353) );
  AND2_X2 U389 ( .A1(n409), .A2(n407), .ZN(n406) );
  AND2_X2 U390 ( .A1(n411), .A2(n475), .ZN(n474) );
  AND2_X1 U391 ( .A1(n373), .A2(n367), .ZN(n366) );
  NAND2_X1 U392 ( .A1(n372), .A2(n371), .ZN(n370) );
  AND2_X1 U393 ( .A1(n685), .A2(n371), .ZN(n364) );
  NOR2_X1 U394 ( .A1(n453), .A2(n476), .ZN(n655) );
  BUF_X1 U395 ( .A(G116), .Z(n690) );
  INV_X1 U396 ( .A(KEYINPUT103), .ZN(n521) );
  INV_X1 U397 ( .A(KEYINPUT4), .ZN(n452) );
  INV_X1 U398 ( .A(KEYINPUT120), .ZN(n377) );
  NAND2_X1 U399 ( .A1(n385), .A2(n354), .ZN(n378) );
  XNOR2_X1 U400 ( .A(n386), .B(n696), .ZN(n385) );
  AND2_X1 U401 ( .A1(n439), .A2(n440), .ZN(n479) );
  AND2_X1 U402 ( .A1(n422), .A2(n539), .ZN(n465) );
  AND2_X1 U403 ( .A1(n456), .A2(n455), .ZN(n709) );
  NAND2_X1 U404 ( .A1(n366), .A2(n363), .ZN(n610) );
  NAND2_X1 U405 ( .A1(n429), .A2(n428), .ZN(n457) );
  XNOR2_X1 U406 ( .A(n430), .B(KEYINPUT46), .ZN(n429) );
  NAND2_X1 U407 ( .A1(n370), .A2(n368), .ZN(n367) );
  NAND2_X1 U408 ( .A1(n365), .A2(n364), .ZN(n363) );
  XNOR2_X1 U409 ( .A(n669), .B(KEYINPUT106), .ZN(n799) );
  NOR2_X1 U410 ( .A1(n798), .A2(n796), .ZN(n430) );
  XNOR2_X1 U411 ( .A(n447), .B(n661), .ZN(n796) );
  XNOR2_X1 U412 ( .A(n656), .B(KEYINPUT39), .ZN(n670) );
  NOR2_X1 U413 ( .A1(n635), .A2(n636), .ZN(n663) );
  XNOR2_X1 U414 ( .A(n454), .B(KEYINPUT30), .ZN(n453) );
  OR2_X1 U415 ( .A1(n607), .A2(KEYINPUT101), .ZN(n369) );
  INV_X1 U416 ( .A(n704), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n568), .B(n567), .ZN(n606) );
  INV_X1 U418 ( .A(n676), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n702), .B(n703), .ZN(n704) );
  INV_X1 U420 ( .A(n699), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U422 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U423 ( .A1(n623), .A2(n548), .ZN(n549) );
  XNOR2_X1 U424 ( .A(n575), .B(n451), .ZN(n707) );
  NAND2_X1 U425 ( .A1(n419), .A2(n416), .ZN(n554) );
  XNOR2_X1 U426 ( .A(n535), .B(G137), .ZN(n451) );
  XNOR2_X1 U427 ( .A(n387), .B(n388), .ZN(n381) );
  XNOR2_X1 U428 ( .A(n537), .B(n491), .ZN(n575) );
  NAND2_X1 U429 ( .A1(n420), .A2(G224), .ZN(n387) );
  XNOR2_X1 U430 ( .A(G122), .B(KEYINPUT100), .ZN(n569) );
  XNOR2_X2 U431 ( .A(G146), .B(G125), .ZN(n536) );
  XNOR2_X1 U432 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n511) );
  XNOR2_X1 U433 ( .A(G119), .B(G116), .ZN(n523) );
  XNOR2_X1 U434 ( .A(G107), .B(G104), .ZN(n361) );
  XNOR2_X2 U435 ( .A(KEYINPUT5), .B(KEYINPUT77), .ZN(n412) );
  NAND2_X1 U436 ( .A1(n666), .A2(n519), .ZN(n391) );
  INV_X1 U437 ( .A(n720), .ZN(n354) );
  XNOR2_X1 U438 ( .A(n700), .B(n356), .ZN(n355) );
  XNOR2_X1 U439 ( .A(n677), .B(n358), .ZN(n357) );
  XNOR2_X1 U440 ( .A(n705), .B(n360), .ZN(n359) );
  XNOR2_X2 U441 ( .A(n362), .B(n361), .ZN(n788) );
  XNOR2_X2 U442 ( .A(n492), .B(G110), .ZN(n362) );
  INV_X1 U443 ( .A(n375), .ZN(n365) );
  NAND2_X1 U444 ( .A1(n685), .A2(n369), .ZN(n368) );
  INV_X1 U445 ( .A(KEYINPUT101), .ZN(n371) );
  INV_X1 U446 ( .A(n685), .ZN(n372) );
  NAND2_X1 U447 ( .A1(n375), .A2(n374), .ZN(n373) );
  AND2_X1 U448 ( .A1(n607), .A2(KEYINPUT101), .ZN(n374) );
  XNOR2_X2 U449 ( .A(n604), .B(KEYINPUT96), .ZN(n375) );
  NAND2_X1 U450 ( .A1(n376), .A2(n402), .ZN(n411) );
  OR2_X1 U451 ( .A1(n395), .A2(n376), .ZN(n473) );
  OR2_X1 U452 ( .A1(n376), .A2(n595), .ZN(n684) );
  OR2_X1 U453 ( .A1(n376), .A2(n609), .ZN(n685) );
  XNOR2_X2 U454 ( .A(n410), .B(KEYINPUT22), .ZN(n376) );
  XNOR2_X1 U455 ( .A(n398), .B(n380), .ZN(n379) );
  XNOR2_X2 U456 ( .A(n739), .B(KEYINPUT6), .ZN(n634) );
  NAND2_X2 U457 ( .A1(n406), .A2(n405), .ZN(n410) );
  XNOR2_X1 U458 ( .A(n378), .B(n377), .ZN(G54) );
  XNOR2_X2 U459 ( .A(n789), .B(n379), .ZN(n389) );
  XNOR2_X1 U460 ( .A(n535), .B(n381), .ZN(n380) );
  XNOR2_X2 U461 ( .A(n534), .B(n533), .ZN(n789) );
  XNOR2_X2 U462 ( .A(n382), .B(n523), .ZN(n534) );
  XNOR2_X2 U463 ( .A(n522), .B(n524), .ZN(n382) );
  AND2_X1 U464 ( .A1(n383), .A2(n354), .ZN(G66) );
  XNOR2_X1 U465 ( .A(n384), .B(n717), .ZN(n383) );
  NAND2_X1 U466 ( .A1(n716), .A2(G217), .ZN(n384) );
  NAND2_X1 U467 ( .A1(n716), .A2(G469), .ZN(n386) );
  NAND2_X2 U468 ( .A1(n444), .A2(n445), .ZN(n716) );
  XNOR2_X2 U469 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n388) );
  NAND2_X1 U470 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X2 U471 ( .A(n389), .B(n469), .ZN(n471) );
  NAND2_X1 U472 ( .A1(n390), .A2(n634), .ZN(n464) );
  XNOR2_X1 U473 ( .A(n599), .B(n521), .ZN(n390) );
  XNOR2_X2 U474 ( .A(n391), .B(n520), .ZN(n599) );
  NAND2_X1 U475 ( .A1(n597), .A2(n392), .ZN(n613) );
  INV_X1 U476 ( .A(KEYINPUT44), .ZN(n392) );
  XNOR2_X1 U477 ( .A(n597), .B(n353), .ZN(G24) );
  XNOR2_X2 U478 ( .A(n587), .B(n393), .ZN(n597) );
  INV_X1 U479 ( .A(n586), .ZN(n393) );
  NAND2_X1 U480 ( .A1(n542), .A2(G214), .ZN(n724) );
  NOR2_X1 U481 ( .A1(n799), .A2(n671), .ZN(n455) );
  XNOR2_X1 U482 ( .A(n457), .B(n403), .ZN(n456) );
  XNOR2_X1 U483 ( .A(n659), .B(n448), .ZN(n755) );
  INV_X1 U484 ( .A(KEYINPUT41), .ZN(n448) );
  INV_X1 U485 ( .A(KEYINPUT90), .ZN(n596) );
  XOR2_X1 U486 ( .A(G131), .B(G140), .Z(n560) );
  NAND2_X1 U487 ( .A1(n641), .A2(n724), .ZN(n454) );
  INV_X1 U488 ( .A(KEYINPUT10), .ZN(n507) );
  NAND2_X1 U489 ( .A1(n655), .A2(n400), .ZN(n656) );
  XNOR2_X1 U490 ( .A(n663), .B(n426), .ZN(n425) );
  INV_X1 U491 ( .A(KEYINPUT109), .ZN(n426) );
  INV_X1 U492 ( .A(G475), .ZN(n566) );
  NOR2_X1 U493 ( .A1(G237), .A2(KEYINPUT79), .ZN(n421) );
  INV_X1 U494 ( .A(G953), .ZN(n420) );
  NAND2_X1 U495 ( .A1(G953), .A2(KEYINPUT79), .ZN(n417) );
  NAND2_X1 U496 ( .A1(n423), .A2(n468), .ZN(n422) );
  INV_X1 U497 ( .A(n709), .ZN(n423) );
  NAND2_X1 U498 ( .A1(KEYINPUT64), .A2(KEYINPUT87), .ZN(n485) );
  AND2_X1 U499 ( .A1(n468), .A2(n485), .ZN(n442) );
  NOR2_X1 U500 ( .A1(n470), .A2(n487), .ZN(n486) );
  INV_X1 U501 ( .A(G237), .ZN(n540) );
  NAND2_X1 U502 ( .A1(n554), .A2(G210), .ZN(n415) );
  INV_X1 U503 ( .A(KEYINPUT88), .ZN(n662) );
  XNOR2_X1 U504 ( .A(n613), .B(KEYINPUT67), .ZN(n615) );
  AND2_X1 U505 ( .A1(n418), .A2(n417), .ZN(n416) );
  NAND2_X1 U506 ( .A1(n421), .A2(n780), .ZN(n419) );
  NAND2_X1 U507 ( .A1(G237), .A2(KEYINPUT79), .ZN(n418) );
  NOR2_X1 U508 ( .A1(n461), .A2(KEYINPUT64), .ZN(n459) );
  NAND2_X1 U509 ( .A1(G234), .A2(G237), .ZN(n545) );
  INV_X1 U510 ( .A(G902), .ZN(n579) );
  AND2_X1 U511 ( .A1(n589), .A2(n408), .ZN(n407) );
  NAND2_X1 U512 ( .A1(n549), .A2(n484), .ZN(n408) );
  XNOR2_X1 U513 ( .A(KEYINPUT16), .B(G122), .ZN(n532) );
  XNOR2_X1 U514 ( .A(G119), .B(G110), .ZN(n501) );
  XNOR2_X1 U515 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n500) );
  XOR2_X1 U516 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n570) );
  INV_X1 U517 ( .A(G134), .ZN(n491) );
  INV_X1 U518 ( .A(KEYINPUT34), .ZN(n553) );
  NAND2_X1 U519 ( .A1(n519), .A2(n477), .ZN(n476) );
  INV_X1 U520 ( .A(n642), .ZN(n477) );
  BUF_X1 U521 ( .A(n601), .Z(n653) );
  XNOR2_X1 U522 ( .A(n565), .B(n564), .ZN(n698) );
  XNOR2_X1 U523 ( .A(n708), .B(n563), .ZN(n564) );
  NOR2_X1 U524 ( .A1(n780), .A2(G952), .ZN(n720) );
  INV_X1 U525 ( .A(KEYINPUT85), .ZN(n462) );
  NAND2_X1 U526 ( .A1(n755), .A2(n660), .ZN(n447) );
  XNOR2_X1 U527 ( .A(n450), .B(n449), .ZN(n798) );
  INV_X1 U528 ( .A(KEYINPUT40), .ZN(n449) );
  XNOR2_X1 U529 ( .A(n424), .B(KEYINPUT36), .ZN(n639) );
  NAND2_X1 U530 ( .A1(n425), .A2(n638), .ZN(n424) );
  NAND2_X1 U531 ( .A1(n592), .A2(n402), .ZN(n475) );
  OR2_X1 U532 ( .A1(n673), .A2(KEYINPUT2), .ZN(n394) );
  INV_X1 U533 ( .A(n549), .ZN(n431) );
  OR2_X1 U534 ( .A1(n592), .A2(n402), .ZN(n395) );
  AND2_X1 U535 ( .A1(n431), .A2(n551), .ZN(n396) );
  INV_X1 U536 ( .A(KEYINPUT64), .ZN(n487) );
  XOR2_X1 U537 ( .A(n498), .B(KEYINPUT1), .Z(n397) );
  XOR2_X1 U538 ( .A(n537), .B(n536), .Z(n398) );
  XOR2_X1 U539 ( .A(KEYINPUT84), .B(n651), .Z(n399) );
  AND2_X1 U540 ( .A1(n725), .A2(n654), .ZN(n400) );
  AND2_X1 U541 ( .A1(n458), .A2(n462), .ZN(n401) );
  XNOR2_X1 U542 ( .A(KEYINPUT82), .B(KEYINPUT32), .ZN(n402) );
  INV_X1 U543 ( .A(n539), .ZN(n470) );
  INV_X1 U544 ( .A(n394), .ZN(n461) );
  INV_X1 U545 ( .A(KEYINPUT87), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n662), .B(KEYINPUT48), .ZN(n403) );
  AND2_X1 U547 ( .A1(n487), .A2(n488), .ZN(n404) );
  OR2_X1 U548 ( .A1(n432), .A2(n551), .ZN(n405) );
  NAND2_X1 U549 ( .A1(n432), .A2(n396), .ZN(n409) );
  NAND2_X1 U550 ( .A1(n474), .A2(n473), .ZN(n691) );
  XNOR2_X1 U551 ( .A(n412), .B(KEYINPUT95), .ZN(n413) );
  XNOR2_X1 U552 ( .A(n413), .B(n525), .ZN(n414) );
  XNOR2_X1 U553 ( .A(n414), .B(n415), .ZN(n526) );
  NOR2_X1 U554 ( .A1(n777), .A2(n427), .ZN(n428) );
  NAND2_X1 U555 ( .A1(n652), .A2(n399), .ZN(n427) );
  XNOR2_X1 U556 ( .A(n637), .B(n433), .ZN(n432) );
  INV_X1 U557 ( .A(n544), .ZN(n433) );
  INV_X1 U558 ( .A(n519), .ZN(n733) );
  XNOR2_X2 U559 ( .A(n601), .B(n397), .ZN(n666) );
  NAND2_X1 U560 ( .A1(n781), .A2(n709), .ZN(n458) );
  BUF_X1 U561 ( .A(n599), .Z(n434) );
  NOR2_X2 U562 ( .A1(n436), .A2(n549), .ZN(n435) );
  XNOR2_X1 U563 ( .A(n637), .B(n544), .ZN(n436) );
  INV_X1 U564 ( .A(n458), .ZN(n460) );
  BUF_X1 U565 ( .A(n788), .Z(n437) );
  NAND2_X1 U566 ( .A1(n474), .A2(n473), .ZN(n438) );
  NAND2_X1 U567 ( .A1(n467), .A2(n468), .ZN(n466) );
  NAND2_X1 U568 ( .A1(n458), .A2(n442), .ZN(n439) );
  OR2_X1 U569 ( .A1(n441), .A2(n486), .ZN(n440) );
  INV_X1 U570 ( .A(n485), .ZN(n441) );
  BUF_X1 U571 ( .A(n731), .Z(n756) );
  XNOR2_X1 U572 ( .A(n435), .B(n484), .ZN(n443) );
  XNOR2_X2 U573 ( .A(n543), .B(KEYINPUT91), .ZN(n637) );
  INV_X1 U574 ( .A(KEYINPUT2), .ZN(n468) );
  AND2_X2 U575 ( .A1(n480), .A2(n481), .ZN(n444) );
  NAND2_X1 U576 ( .A1(n479), .A2(n478), .ZN(n445) );
  NAND2_X1 U577 ( .A1(n460), .A2(n394), .ZN(n478) );
  XNOR2_X2 U578 ( .A(n446), .B(n596), .ZN(n614) );
  NAND2_X1 U579 ( .A1(n691), .A2(n684), .ZN(n446) );
  NAND2_X1 U580 ( .A1(n670), .A2(n773), .ZN(n450) );
  XNOR2_X2 U581 ( .A(n452), .B(KEYINPUT68), .ZN(n535) );
  XNOR2_X2 U582 ( .A(G143), .B(G128), .ZN(n537) );
  NAND2_X1 U583 ( .A1(n460), .A2(n459), .ZN(n480) );
  XNOR2_X1 U584 ( .A(n463), .B(n553), .ZN(n584) );
  NAND2_X1 U585 ( .A1(n466), .A2(n465), .ZN(n482) );
  INV_X1 U586 ( .A(n781), .ZN(n467) );
  INV_X1 U587 ( .A(n471), .ZN(n702) );
  INV_X1 U588 ( .A(n538), .ZN(n469) );
  XNOR2_X2 U589 ( .A(n618), .B(KEYINPUT45), .ZN(n781) );
  NAND2_X1 U590 ( .A1(n482), .A2(n404), .ZN(n481) );
  NAND2_X1 U591 ( .A1(n483), .A2(KEYINPUT44), .ZN(n611) );
  NAND2_X1 U592 ( .A1(n614), .A2(n597), .ZN(n483) );
  INV_X1 U593 ( .A(n551), .ZN(n484) );
  NAND2_X1 U594 ( .A1(n688), .A2(n765), .ZN(n604) );
  XNOR2_X2 U595 ( .A(n489), .B(n600), .ZN(n688) );
  NAND2_X1 U596 ( .A1(n443), .A2(n490), .ZN(n489) );
  INV_X1 U597 ( .A(n744), .ZN(n490) );
  BUF_X1 U598 ( .A(n534), .Z(n527) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n593) );
  XNOR2_X1 U600 ( .A(n566), .B(KEYINPUT13), .ZN(n567) );
  XNOR2_X1 U601 ( .A(n707), .B(G146), .ZN(n528) );
  XNOR2_X2 U602 ( .A(G101), .B(KEYINPUT78), .ZN(n492) );
  XNOR2_X2 U603 ( .A(n788), .B(KEYINPUT73), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n780), .A2(G227), .ZN(n493) );
  XNOR2_X1 U605 ( .A(n560), .B(n493), .ZN(n494) );
  XNOR2_X1 U606 ( .A(n538), .B(n494), .ZN(n495) );
  XNOR2_X1 U607 ( .A(n495), .B(n528), .ZN(n693) );
  NAND2_X1 U608 ( .A1(n693), .A2(n579), .ZN(n497) );
  INV_X1 U609 ( .A(G469), .ZN(n496) );
  XNOR2_X2 U610 ( .A(n497), .B(n496), .ZN(n601) );
  INV_X1 U611 ( .A(KEYINPUT65), .ZN(n498) );
  NAND2_X1 U612 ( .A1(n780), .A2(G234), .ZN(n499) );
  XNOR2_X1 U613 ( .A(n500), .B(n499), .ZN(n574) );
  NAND2_X1 U614 ( .A1(n574), .A2(G221), .ZN(n504) );
  XOR2_X1 U615 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n502) );
  XNOR2_X1 U616 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U617 ( .A(n504), .B(n503), .ZN(n510) );
  XOR2_X1 U618 ( .A(KEYINPUT94), .B(G140), .Z(n506) );
  XNOR2_X1 U619 ( .A(n506), .B(n505), .ZN(n508) );
  XNOR2_X1 U620 ( .A(n536), .B(n507), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n508), .B(n559), .ZN(n509) );
  XNOR2_X1 U622 ( .A(n510), .B(n509), .ZN(n717) );
  NAND2_X1 U623 ( .A1(n717), .A2(n579), .ZN(n515) );
  XNOR2_X1 U624 ( .A(n511), .B(G902), .ZN(n672) );
  NAND2_X1 U625 ( .A1(G234), .A2(n672), .ZN(n512) );
  XNOR2_X1 U626 ( .A(n512), .B(KEYINPUT20), .ZN(n516) );
  NAND2_X1 U627 ( .A1(G217), .A2(n516), .ZN(n513) );
  XNOR2_X1 U628 ( .A(n513), .B(KEYINPUT25), .ZN(n514) );
  XNOR2_X1 U629 ( .A(n515), .B(n514), .ZN(n626) );
  NAND2_X1 U630 ( .A1(n516), .A2(G221), .ZN(n518) );
  INV_X1 U631 ( .A(KEYINPUT21), .ZN(n517) );
  XNOR2_X1 U632 ( .A(n518), .B(n517), .ZN(n736) );
  INV_X1 U633 ( .A(n736), .ZN(n624) );
  INV_X1 U634 ( .A(KEYINPUT76), .ZN(n520) );
  XNOR2_X2 U635 ( .A(G113), .B(KEYINPUT71), .ZN(n522) );
  XNOR2_X2 U636 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n524) );
  XNOR2_X1 U637 ( .A(n527), .B(n526), .ZN(n529) );
  XNOR2_X1 U638 ( .A(n529), .B(n528), .ZN(n675) );
  NAND2_X1 U639 ( .A1(n675), .A2(n579), .ZN(n531) );
  INV_X1 U640 ( .A(G472), .ZN(n530) );
  BUF_X2 U641 ( .A(n593), .Z(n739) );
  XNOR2_X1 U642 ( .A(n532), .B(KEYINPUT74), .ZN(n533) );
  INV_X1 U643 ( .A(n672), .ZN(n539) );
  NAND2_X1 U644 ( .A1(n579), .A2(n540), .ZN(n542) );
  AND2_X1 U645 ( .A1(n542), .A2(G210), .ZN(n541) );
  XNOR2_X1 U646 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n544) );
  XOR2_X1 U647 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n546) );
  XNOR2_X1 U648 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U649 ( .A1(G952), .A2(n547), .ZN(n752) );
  NOR2_X1 U650 ( .A1(n752), .A2(G953), .ZN(n623) );
  NAND2_X1 U651 ( .A1(G902), .A2(n547), .ZN(n619) );
  XNOR2_X1 U652 ( .A(G898), .B(KEYINPUT93), .ZN(n784) );
  NAND2_X1 U653 ( .A1(G953), .A2(n784), .ZN(n790) );
  NOR2_X1 U654 ( .A1(n619), .A2(n790), .ZN(n548) );
  INV_X1 U655 ( .A(KEYINPUT66), .ZN(n550) );
  XNOR2_X1 U656 ( .A(n550), .B(KEYINPUT0), .ZN(n551) );
  BUF_X1 U657 ( .A(n443), .Z(n552) );
  NAND2_X1 U658 ( .A1(G214), .A2(n554), .ZN(n555) );
  XNOR2_X1 U659 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U660 ( .A(G122), .B(G104), .Z(n557) );
  XNOR2_X1 U661 ( .A(n558), .B(n557), .ZN(n565) );
  XNOR2_X1 U662 ( .A(n560), .B(n559), .ZN(n708) );
  XOR2_X1 U663 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n562) );
  XNOR2_X1 U664 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n561) );
  XNOR2_X1 U665 ( .A(n562), .B(n561), .ZN(n563) );
  NOR2_X1 U666 ( .A1(G902), .A2(n698), .ZN(n568) );
  INV_X1 U667 ( .A(n606), .ZN(n582) );
  XNOR2_X1 U668 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U669 ( .A(n571), .B(KEYINPUT7), .Z(n573) );
  XNOR2_X1 U670 ( .A(n690), .B(G107), .ZN(n572) );
  XNOR2_X1 U671 ( .A(n573), .B(n572), .ZN(n578) );
  AND2_X1 U672 ( .A1(n574), .A2(G217), .ZN(n576) );
  XNOR2_X1 U673 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U674 ( .A(n578), .B(n577), .ZN(n719) );
  NAND2_X1 U675 ( .A1(n719), .A2(n579), .ZN(n581) );
  INV_X1 U676 ( .A(G478), .ZN(n580) );
  XNOR2_X1 U677 ( .A(n581), .B(n580), .ZN(n588) );
  INV_X1 U678 ( .A(n588), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n582), .A2(n605), .ZN(n646) );
  INV_X1 U680 ( .A(n646), .ZN(n583) );
  NAND2_X1 U681 ( .A1(n584), .A2(n583), .ZN(n587) );
  INV_X1 U682 ( .A(KEYINPUT81), .ZN(n585) );
  XNOR2_X1 U683 ( .A(n585), .B(KEYINPUT35), .ZN(n586) );
  NAND2_X1 U684 ( .A1(n606), .A2(n588), .ZN(n727) );
  NOR2_X1 U685 ( .A1(n727), .A2(n624), .ZN(n589) );
  XNOR2_X1 U686 ( .A(n634), .B(KEYINPUT83), .ZN(n591) );
  INV_X1 U687 ( .A(n666), .ZN(n734) );
  INV_X1 U688 ( .A(n626), .ZN(n737) );
  NOR2_X1 U689 ( .A1(n734), .A2(n737), .ZN(n590) );
  NAND2_X1 U690 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U691 ( .A(n593), .B(KEYINPUT102), .ZN(n640) );
  AND2_X1 U692 ( .A1(n640), .A2(n626), .ZN(n594) );
  NAND2_X1 U693 ( .A1(n594), .A2(n734), .ZN(n595) );
  INV_X1 U694 ( .A(n739), .ZN(n598) );
  NAND2_X1 U695 ( .A1(n434), .A2(n598), .ZN(n744) );
  INV_X1 U696 ( .A(KEYINPUT31), .ZN(n600) );
  NAND2_X1 U697 ( .A1(n739), .A2(n519), .ZN(n602) );
  NOR2_X1 U698 ( .A1(n602), .A2(n653), .ZN(n603) );
  NAND2_X1 U699 ( .A1(n552), .A2(n603), .ZN(n765) );
  NOR2_X1 U700 ( .A1(n606), .A2(n605), .ZN(n773) );
  AND2_X1 U701 ( .A1(n606), .A2(n605), .ZN(n769) );
  NOR2_X1 U702 ( .A1(n773), .A2(n769), .ZN(n723) );
  INV_X1 U703 ( .A(n723), .ZN(n607) );
  NOR2_X1 U704 ( .A1(n634), .A2(n626), .ZN(n608) );
  NAND2_X1 U705 ( .A1(n608), .A2(n734), .ZN(n609) );
  NAND2_X1 U706 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U707 ( .A(n612), .B(KEYINPUT89), .ZN(n617) );
  NAND2_X1 U708 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U709 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U710 ( .A1(G900), .A2(n619), .ZN(n620) );
  NAND2_X1 U711 ( .A1(G953), .A2(n620), .ZN(n621) );
  XOR2_X1 U712 ( .A(KEYINPUT104), .B(n621), .Z(n622) );
  NOR2_X1 U713 ( .A1(n623), .A2(n622), .ZN(n642) );
  NOR2_X1 U714 ( .A1(n624), .A2(n642), .ZN(n625) );
  NAND2_X1 U715 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U716 ( .A(KEYINPUT70), .B(n627), .ZN(n636) );
  NOR2_X1 U717 ( .A1(n636), .A2(n640), .ZN(n628) );
  XNOR2_X1 U718 ( .A(n628), .B(KEYINPUT28), .ZN(n630) );
  XNOR2_X1 U719 ( .A(n653), .B(KEYINPUT107), .ZN(n629) );
  NAND2_X1 U720 ( .A1(n630), .A2(n629), .ZN(n657) );
  BUF_X1 U721 ( .A(n436), .Z(n631) );
  NOR2_X1 U722 ( .A1(n657), .A2(n631), .ZN(n774) );
  XOR2_X1 U723 ( .A(KEYINPUT47), .B(n774), .Z(n633) );
  NAND2_X1 U724 ( .A1(n774), .A2(n723), .ZN(n632) );
  NAND2_X1 U725 ( .A1(n633), .A2(n632), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n634), .A2(n773), .ZN(n635) );
  BUF_X1 U727 ( .A(n637), .Z(n638) );
  NOR2_X1 U728 ( .A1(n734), .A2(n639), .ZN(n777) );
  INV_X1 U729 ( .A(n640), .ZN(n641) );
  BUF_X1 U730 ( .A(n643), .Z(n644) );
  INV_X1 U731 ( .A(n644), .ZN(n645) );
  OR2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U733 ( .A1(n647), .A2(n653), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n655), .A2(n648), .ZN(n680) );
  XNOR2_X1 U735 ( .A(n680), .B(KEYINPUT86), .ZN(n650) );
  NAND2_X1 U736 ( .A1(KEYINPUT47), .A2(n723), .ZN(n649) );
  NAND2_X1 U737 ( .A1(n650), .A2(n649), .ZN(n651) );
  INV_X1 U738 ( .A(n653), .ZN(n654) );
  XNOR2_X1 U739 ( .A(n644), .B(KEYINPUT38), .ZN(n658) );
  XOR2_X1 U740 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n661) );
  INV_X1 U741 ( .A(n657), .ZN(n660) );
  INV_X1 U742 ( .A(n658), .ZN(n725) );
  NAND2_X1 U743 ( .A1(n725), .A2(n724), .ZN(n722) );
  NOR2_X1 U744 ( .A1(n727), .A2(n722), .ZN(n659) );
  NAND2_X1 U745 ( .A1(n663), .A2(n724), .ZN(n664) );
  XOR2_X1 U746 ( .A(KEYINPUT105), .B(n664), .Z(n665) );
  NOR2_X1 U747 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n667), .B(KEYINPUT43), .ZN(n668) );
  NOR2_X1 U749 ( .A1(n668), .A2(n644), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n670), .A2(n769), .ZN(n779) );
  INV_X1 U751 ( .A(n779), .ZN(n671) );
  NOR2_X1 U752 ( .A1(n672), .A2(n488), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n716), .A2(G472), .ZN(n677) );
  XOR2_X1 U754 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n674) );
  INV_X1 U755 ( .A(KEYINPUT63), .ZN(n678) );
  XNOR2_X1 U756 ( .A(n680), .B(G143), .ZN(G45) );
  INV_X1 U757 ( .A(n773), .ZN(n686) );
  NOR2_X1 U758 ( .A1(n765), .A2(n686), .ZN(n682) );
  XNOR2_X1 U759 ( .A(G104), .B(KEYINPUT111), .ZN(n681) );
  XNOR2_X1 U760 ( .A(n682), .B(n681), .ZN(G6) );
  XNOR2_X1 U761 ( .A(G110), .B(KEYINPUT112), .ZN(n683) );
  XNOR2_X1 U762 ( .A(n684), .B(n683), .ZN(G12) );
  XNOR2_X1 U763 ( .A(n685), .B(G101), .ZN(G3) );
  NOR2_X1 U764 ( .A1(n688), .A2(n686), .ZN(n687) );
  XOR2_X1 U765 ( .A(G113), .B(n687), .Z(G15) );
  INV_X1 U766 ( .A(n769), .ZN(n764) );
  NOR2_X1 U767 ( .A1(n688), .A2(n764), .ZN(n689) );
  XOR2_X1 U768 ( .A(n690), .B(n689), .Z(G18) );
  XNOR2_X1 U769 ( .A(G119), .B(KEYINPUT126), .ZN(n692) );
  XNOR2_X1 U770 ( .A(n438), .B(n692), .ZN(G21) );
  BUF_X1 U771 ( .A(n693), .Z(n695) );
  XNOR2_X1 U772 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n694) );
  NAND2_X1 U773 ( .A1(n716), .A2(G475), .ZN(n700) );
  XNOR2_X1 U774 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n697) );
  NAND2_X1 U775 ( .A1(n716), .A2(G210), .ZN(n705) );
  XOR2_X1 U776 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n703) );
  XOR2_X1 U777 ( .A(n708), .B(n707), .Z(n711) );
  XOR2_X1 U778 ( .A(n711), .B(n709), .Z(n710) );
  NAND2_X1 U779 ( .A1(n710), .A2(n780), .ZN(n715) );
  XNOR2_X1 U780 ( .A(G227), .B(n711), .ZN(n712) );
  NAND2_X1 U781 ( .A1(G900), .A2(n712), .ZN(n713) );
  NAND2_X1 U782 ( .A1(n713), .A2(G953), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n715), .A2(n714), .ZN(G72) );
  NAND2_X1 U784 ( .A1(n716), .A2(G478), .ZN(n718) );
  XOR2_X1 U785 ( .A(n719), .B(n718), .Z(n721) );
  NOR2_X1 U786 ( .A1(n721), .A2(n720), .ZN(G63) );
  XNOR2_X1 U787 ( .A(n401), .B(KEYINPUT2), .ZN(n761) );
  XOR2_X1 U788 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n751) );
  OR2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n730) );
  NOR2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U792 ( .A(KEYINPUT116), .B(n728), .Z(n729) );
  NAND2_X1 U793 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U794 ( .A1(n732), .A2(n756), .ZN(n749) );
  NAND2_X1 U795 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U796 ( .A(n735), .B(KEYINPUT50), .ZN(n743) );
  NOR2_X1 U797 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U798 ( .A(n738), .B(KEYINPUT49), .ZN(n740) );
  NAND2_X1 U799 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U800 ( .A(KEYINPUT115), .B(n741), .ZN(n742) );
  NAND2_X1 U801 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U802 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U803 ( .A(KEYINPUT51), .B(n746), .Z(n747) );
  NAND2_X1 U804 ( .A1(n755), .A2(n747), .ZN(n748) );
  NAND2_X1 U805 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U806 ( .A(n751), .B(n750), .Z(n753) );
  NOR2_X1 U807 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U808 ( .A1(n754), .A2(G953), .ZN(n759) );
  NAND2_X1 U809 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U810 ( .A(n757), .B(KEYINPUT118), .ZN(n758) );
  NAND2_X1 U811 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n763) );
  XOR2_X1 U813 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n762) );
  XNOR2_X1 U814 ( .A(n763), .B(n762), .ZN(G75) );
  NOR2_X1 U815 ( .A1(n765), .A2(n764), .ZN(n767) );
  XNOR2_X1 U816 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n766) );
  XNOR2_X1 U817 ( .A(n767), .B(n766), .ZN(n768) );
  XNOR2_X1 U818 ( .A(G107), .B(n768), .ZN(G9) );
  XOR2_X1 U819 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n771) );
  NAND2_X1 U820 ( .A1(n774), .A2(n769), .ZN(n770) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(n772) );
  XOR2_X1 U822 ( .A(G128), .B(n772), .Z(G30) );
  NAND2_X1 U823 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U824 ( .A(n775), .B(KEYINPUT114), .ZN(n776) );
  XNOR2_X1 U825 ( .A(G146), .B(n776), .ZN(G48) );
  XNOR2_X1 U826 ( .A(G125), .B(n777), .ZN(n778) );
  XNOR2_X1 U827 ( .A(n778), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U828 ( .A(G134), .B(n779), .ZN(G36) );
  AND2_X1 U829 ( .A1(n781), .A2(n780), .ZN(n786) );
  NAND2_X1 U830 ( .A1(G953), .A2(G224), .ZN(n782) );
  XOR2_X1 U831 ( .A(KEYINPUT61), .B(n782), .Z(n783) );
  NOR2_X1 U832 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U833 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U834 ( .A(n787), .B(KEYINPUT124), .ZN(n795) );
  XOR2_X1 U835 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n793) );
  XNOR2_X1 U836 ( .A(n789), .B(n437), .ZN(n791) );
  NAND2_X1 U837 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U838 ( .A(n793), .B(n792), .ZN(n794) );
  XNOR2_X1 U839 ( .A(n795), .B(n794), .ZN(G69) );
  XNOR2_X1 U840 ( .A(G137), .B(n796), .ZN(n797) );
  XNOR2_X1 U841 ( .A(n797), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U842 ( .A(G131), .B(n798), .Z(G33) );
  XOR2_X1 U843 ( .A(G140), .B(n799), .Z(G42) );
endmodule

