//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(G125), .ZN(new_n194));
  INV_X1    g008(.A(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n197), .B2(new_n191), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT75), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT75), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n202), .A3(new_n199), .ZN(new_n203));
  OAI211_X1 g017(.A(G146), .B(new_n193), .C1(new_n197), .C2(new_n191), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n204), .A2(KEYINPUT74), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(KEYINPUT74), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n201), .B(new_n203), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  XOR2_X1   g021(.A(G119), .B(G128), .Z(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT24), .B(G110), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n211), .B(G119), .C1(KEYINPUT72), .C2(KEYINPUT23), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n213));
  INV_X1    g027(.A(G119), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G128), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT72), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n214), .B2(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G110), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT73), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(KEYINPUT73), .A3(G110), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n210), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n204), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n208), .A2(new_n209), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n218), .B2(G110), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n194), .A2(new_n196), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n199), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n207), .A2(new_n223), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n190), .B1(new_n231), .B2(KEYINPUT77), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n207), .A2(new_n223), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n225), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n190), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G217), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(G234), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G902), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT78), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT78), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n248), .A3(new_n245), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n240), .A2(new_n243), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT25), .ZN(new_n251));
  AOI21_X1  g065(.A(G902), .B1(new_n238), .B2(new_n239), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT25), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n244), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n247), .B(new_n249), .C1(new_n251), .C2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(G472), .A2(G902), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n257));
  INV_X1    g071(.A(G113), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT66), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(KEYINPUT2), .B2(G113), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G116), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G116), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n266), .A3(G119), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT2), .A2(G113), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n263), .A2(G119), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AND4_X1   g084(.A1(new_n262), .A2(new_n267), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n262), .A2(new_n268), .B1(new_n267), .B2(new_n270), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT11), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(G137), .ZN(new_n277));
  INV_X1    g091(.A(G137), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT11), .A3(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(G137), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G131), .ZN(new_n282));
  INV_X1    g096(.A(G131), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n277), .A2(new_n279), .A3(new_n283), .A4(new_n280), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(KEYINPUT65), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(KEYINPUT0), .A2(G128), .ZN(new_n286));
  OR2_X1    g100(.A1(KEYINPUT0), .A2(G128), .ZN(new_n287));
  INV_X1    g101(.A(G143), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(G146), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n199), .A2(G143), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n286), .B(new_n287), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT64), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n288), .B2(G146), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n199), .A2(KEYINPUT64), .A3(G143), .ZN(new_n294));
  INV_X1    g108(.A(new_n286), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n288), .A2(G146), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n293), .A2(new_n294), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n281), .A2(new_n299), .A3(G131), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n285), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT30), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT1), .B1(new_n288), .B2(G146), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n199), .A2(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n296), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n293), .A2(new_n294), .A3(new_n308), .A4(new_n296), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n280), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n276), .A2(G137), .ZN(new_n312));
  OAI21_X1  g126(.A(G131), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n284), .A3(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n301), .A2(new_n302), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n302), .B1(new_n301), .B2(new_n314), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n274), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n301), .A2(new_n273), .A3(new_n314), .ZN(new_n318));
  NOR2_X1   g132(.A1(G237), .A2(G953), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G210), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT27), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT26), .B(G101), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n317), .A2(KEYINPUT31), .A3(new_n318), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n318), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n301), .A2(new_n314), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n274), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n301), .A2(KEYINPUT28), .A3(new_n273), .A4(new_n314), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n323), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT68), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n338), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n328), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n328), .B2(new_n340), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n256), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT70), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n347), .B(new_n256), .C1(new_n342), .C2(new_n343), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n256), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n328), .A2(new_n340), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT69), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n328), .A2(new_n340), .A3(new_n341), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT71), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n332), .A2(new_n355), .A3(new_n318), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n331), .A2(KEYINPUT71), .A3(new_n274), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(KEYINPUT28), .A3(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n358), .A2(KEYINPUT29), .A3(new_n323), .A4(new_n330), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n359), .A2(new_n243), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n317), .A2(new_n318), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n323), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n362), .A2(KEYINPUT29), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n334), .A2(new_n335), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n354), .A2(KEYINPUT32), .B1(G472), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n255), .B1(new_n349), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G478), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(KEYINPUT15), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n288), .A2(G128), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n211), .A2(G143), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT91), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT91), .B1(new_n371), .B2(new_n372), .ZN(new_n374));
  OR3_X1    g188(.A1(new_n373), .A2(new_n374), .A3(new_n276), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n276), .B1(new_n373), .B2(new_n374), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n264), .A2(new_n266), .A3(G122), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n263), .A2(G122), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT14), .A4(G122), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n380), .ZN(new_n383));
  OAI211_X1 g197(.A(G107), .B(new_n382), .C1(new_n383), .C2(KEYINPUT14), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n371), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT13), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n276), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G128), .B(G143), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT13), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n376), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT90), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n383), .A2(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT90), .A3(new_n381), .ZN(new_n398));
  AOI211_X1 g212(.A(KEYINPUT92), .B(new_n392), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n398), .ZN(new_n401));
  INV_X1    g215(.A(new_n392), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n385), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n405), .A2(new_n242), .A3(G953), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n385), .B(new_n406), .C1(new_n399), .C2(new_n403), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n370), .B1(new_n410), .B2(new_n243), .ZN(new_n411));
  AOI211_X1 g225(.A(G902), .B(new_n369), .C1(new_n408), .C2(new_n409), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n198), .A2(new_n202), .A3(new_n199), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n202), .B1(new_n198), .B2(new_n199), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n204), .B(KEYINPUT74), .ZN(new_n417));
  INV_X1    g231(.A(G237), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n188), .A3(G214), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n288), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n319), .A2(G143), .A3(G214), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT17), .A3(G131), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(G131), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n283), .A3(new_n421), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n416), .A2(new_n417), .A3(new_n423), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(KEYINPUT18), .A2(G131), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n422), .B(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n228), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n197), .A2(KEYINPUT86), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(G146), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n229), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n428), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(G113), .B(G122), .Z(new_n438));
  XOR2_X1   g252(.A(KEYINPUT87), .B(G104), .Z(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT89), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n243), .B1(new_n437), .B2(new_n442), .ZN(new_n444));
  OAI21_X1  g258(.A(G475), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n441), .B1(new_n428), .B2(new_n436), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n424), .A2(new_n426), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n432), .A2(KEYINPUT19), .A3(new_n433), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n197), .A2(KEYINPUT19), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n199), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n225), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n440), .B1(new_n430), .B2(new_n435), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(G475), .A2(G902), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT88), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n446), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  NOR4_X1   g273(.A1(new_n447), .A2(new_n454), .A3(KEYINPUT20), .A4(new_n457), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n445), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n243), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(G898), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G952), .ZN(new_n466));
  AOI211_X1 g280(.A(G953), .B(new_n466), .C1(G234), .C2(G237), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n413), .A2(new_n462), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G110), .B(G140), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n188), .A2(G227), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n304), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n309), .ZN(new_n476));
  INV_X1    g290(.A(G104), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT3), .B1(new_n477), .B2(G107), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n379), .A3(G104), .ZN(new_n480));
  INV_X1    g294(.A(G101), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(G107), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n478), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n477), .A2(G107), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n379), .A2(G104), .ZN(new_n485));
  OAI21_X1  g299(.A(G101), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n476), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT10), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n285), .A2(new_n300), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G101), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n483), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n495), .A3(G101), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n298), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n489), .B1(new_n307), .B2(new_n309), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n487), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n490), .A2(new_n491), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n488), .A2(new_n489), .B1(new_n487), .B2(new_n498), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n491), .B1(new_n502), .B2(new_n497), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n473), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT12), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(KEYINPUT12), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n487), .A2(new_n310), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n483), .A2(new_n486), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n309), .B2(new_n475), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n506), .B(new_n508), .C1(new_n512), .C2(new_n491), .ZN(new_n513));
  INV_X1    g327(.A(new_n473), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n488), .B1(new_n310), .B2(new_n487), .ZN(new_n515));
  INV_X1    g329(.A(new_n491), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT12), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n515), .A2(KEYINPUT79), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n513), .A2(new_n514), .A3(new_n500), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n504), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G469), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(new_n243), .ZN(new_n522));
  NAND2_X1  g336(.A1(G469), .A2(G902), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n513), .A2(new_n500), .A3(new_n518), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n473), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n500), .A2(new_n514), .ZN(new_n526));
  INV_X1    g340(.A(new_n503), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(G469), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(G221), .B1(new_n405), .B2(G902), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT80), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(KEYINPUT80), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n267), .A2(KEYINPUT5), .A3(new_n270), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT5), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n258), .B1(new_n269), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n262), .A2(new_n267), .A3(new_n268), .A4(new_n270), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n487), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n496), .B1(new_n271), .B2(new_n272), .ZN(new_n543));
  INV_X1    g357(.A(new_n494), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n546));
  XNOR2_X1  g360(.A(G110), .B(G122), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n545), .A2(KEYINPUT83), .A3(new_n546), .A4(new_n548), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  MUX2_X1   g367(.A(new_n310), .B(new_n298), .S(G125), .Z(new_n554));
  INV_X1    g368(.A(G224), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n555), .A2(G953), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n554), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT82), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n545), .A2(new_n548), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n547), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n561));
  AND4_X1   g375(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT6), .A4(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n546), .B1(new_n545), .B2(new_n548), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n559), .B1(new_n563), .B2(new_n561), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n553), .B(new_n558), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n539), .B(KEYINPUT84), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n566), .A2(new_n537), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n487), .A2(new_n541), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n540), .A2(new_n541), .ZN(new_n569));
  OAI22_X1  g383(.A1(new_n567), .A2(new_n568), .B1(new_n487), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n547), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n554), .A2(KEYINPUT85), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n310), .A2(KEYINPUT85), .A3(G125), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(KEYINPUT7), .B2(new_n557), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n570), .A2(new_n571), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n554), .A2(KEYINPUT7), .A3(new_n557), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n576), .A2(new_n561), .ZN(new_n577));
  AOI21_X1  g391(.A(G902), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n565), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G210), .B1(G237), .B2(G902), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n565), .A2(new_n578), .A3(new_n580), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G214), .B1(G237), .B2(G902), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n586), .B(KEYINPUT81), .Z(new_n587));
  NOR3_X1   g401(.A1(new_n536), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n367), .A2(new_n470), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  OAI21_X1  g404(.A(new_n243), .B1(new_n342), .B2(new_n343), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(new_n345), .A3(new_n348), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n593), .A2(new_n255), .A3(new_n536), .ZN(new_n594));
  INV_X1    g408(.A(new_n586), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n582), .B2(new_n583), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n469), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n392), .B1(new_n396), .B2(new_n398), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n400), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n406), .B1(new_n599), .B2(new_n385), .ZN(new_n600));
  INV_X1    g414(.A(new_n409), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT33), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n408), .A2(new_n603), .A3(new_n409), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(G478), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n368), .A2(new_n243), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n408), .B2(new_n409), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(new_n368), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n461), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n597), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n594), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  OAI21_X1  g428(.A(new_n462), .B1(new_n411), .B2(new_n412), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n597), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n594), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  INV_X1    g433(.A(new_n593), .ZN(new_n620));
  INV_X1    g434(.A(new_n190), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n235), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n245), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n251), .B2(new_n254), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n470), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n620), .A2(new_n588), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT37), .B(G110), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G12));
  NAND4_X1  g443(.A1(new_n534), .A2(new_n596), .A3(new_n625), .A4(new_n535), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n467), .B(KEYINPUT93), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(G900), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(new_n463), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n630), .A2(new_n615), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n349), .A2(new_n366), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  OAI21_X1  g452(.A(new_n461), .B1(new_n411), .B2(new_n412), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n625), .A2(new_n595), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n585), .A2(KEYINPUT38), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n584), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n534), .A2(new_n535), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n634), .B(KEYINPUT39), .Z(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT95), .B(KEYINPUT40), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n644), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT94), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n361), .A2(new_n335), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n356), .A2(new_n357), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n654), .B(new_n243), .C1(new_n323), .C2(new_n655), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n354), .A2(KEYINPUT32), .B1(G472), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n653), .B1(new_n349), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n349), .A2(new_n657), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(KEYINPUT94), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n652), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n652), .B(KEYINPUT96), .C1(new_n658), .C2(new_n660), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  INV_X1    g480(.A(new_n634), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n605), .A2(new_n608), .A3(new_n461), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT97), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n630), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n636), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT98), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n670), .A2(new_n636), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  INV_X1    g490(.A(new_n255), .ZN(new_n677));
  INV_X1    g491(.A(new_n522), .ZN(new_n678));
  INV_X1    g492(.A(new_n531), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n521), .B1(new_n520), .B2(new_n243), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n636), .A2(new_n677), .A3(new_n611), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n636), .A2(new_n677), .A3(new_n616), .A4(new_n681), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NAND2_X1  g500(.A1(new_n596), .A2(new_n681), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n636), .A2(new_n626), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  NAND2_X1  g504(.A1(new_n639), .A2(KEYINPUT102), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n461), .B(new_n692), .C1(new_n411), .C2(new_n412), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n691), .A2(new_n596), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT103), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n691), .A2(new_n596), .A3(new_n696), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT101), .B(G472), .Z(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n591), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n256), .B(KEYINPUT99), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT100), .B1(new_n358), .B2(new_n330), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n323), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT100), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n358), .A2(new_n330), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n703), .B1(new_n708), .B2(new_n328), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n701), .A2(new_n677), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n681), .A2(new_n469), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n698), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  NOR2_X1   g528(.A1(new_n669), .A2(new_n687), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n701), .A2(new_n710), .A3(new_n625), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n715), .A2(new_n717), .A3(KEYINPUT104), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n668), .A2(KEYINPUT97), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n668), .A2(KEYINPUT97), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n688), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n719), .B1(new_n722), .B2(new_n716), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  NAND2_X1  g539(.A1(new_n365), .A2(G472), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n344), .B2(new_n346), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n677), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n731), .B(new_n677), .C1(new_n727), .C2(new_n728), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n524), .A2(new_n473), .B1(new_n526), .B2(new_n527), .ZN(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n735), .B2(G902), .ZN(new_n736));
  AOI211_X1 g550(.A(KEYINPUT105), .B(new_n679), .C1(new_n736), .C2(new_n522), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n530), .B2(new_n531), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n582), .A2(KEYINPUT106), .A3(new_n583), .A4(new_n586), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n740), .A2(new_n743), .A3(new_n747), .A4(new_n744), .ZN(new_n748));
  AOI211_X1 g562(.A(new_n734), .B(new_n669), .C1(new_n746), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n748), .ZN(new_n750));
  INV_X1    g564(.A(new_n669), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n367), .A3(new_n751), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n733), .A2(new_n749), .B1(new_n752), .B2(new_n734), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n283), .ZN(G33));
  NOR2_X1   g568(.A1(new_n615), .A2(new_n634), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n750), .A2(new_n367), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  NAND2_X1  g571(.A1(new_n609), .A2(new_n462), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT43), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n609), .A2(new_n760), .A3(new_n462), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n759), .A2(new_n625), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n593), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n735), .A2(KEYINPUT45), .ZN(new_n766));
  OAI21_X1  g580(.A(G469), .B1(new_n735), .B2(KEYINPUT45), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n523), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n678), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n531), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n646), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n743), .A2(new_n744), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n762), .A2(KEYINPUT44), .A3(new_n593), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n765), .A2(new_n774), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n772), .B(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n636), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n669), .A2(new_n775), .A3(new_n677), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT109), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT109), .B1(new_n783), .B2(new_n784), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n780), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n787), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(KEYINPUT110), .A3(new_n782), .A4(new_n785), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NOR3_X1   g606(.A1(new_n660), .A2(new_n255), .A3(new_n658), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n678), .A2(new_n680), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT111), .Z(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT49), .Z(new_n796));
  AND2_X1   g610(.A1(new_n641), .A2(new_n643), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n797), .A2(new_n587), .A3(new_n679), .A4(new_n758), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n776), .A2(new_n681), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT117), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT117), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n793), .A2(new_n803), .A3(new_n467), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n609), .A2(new_n461), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT118), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n759), .A2(new_n761), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n711), .A3(new_n632), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n681), .A2(new_n595), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT116), .Z(new_n812));
  NOR3_X1   g626(.A1(new_n810), .A2(new_n812), .A3(new_n797), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT50), .Z(new_n814));
  NAND3_X1  g628(.A1(new_n803), .A2(new_n632), .A3(new_n809), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n716), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n795), .A2(new_n531), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n782), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n775), .A3(new_n810), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n814), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n808), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n804), .A2(new_n610), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n810), .A2(new_n687), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n466), .A3(G953), .ZN(new_n826));
  INV_X1    g640(.A(new_n733), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n815), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n828), .A2(KEYINPUT48), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(KEYINPUT48), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n824), .B(new_n826), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n808), .A2(new_n820), .A3(KEYINPUT51), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n823), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n530), .A2(new_n531), .A3(new_n667), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n625), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT113), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n659), .A3(new_n698), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n670), .A2(new_n636), .A3(new_n673), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n673), .B1(new_n670), .B2(new_n636), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT104), .B1(new_n715), .B2(new_n717), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n722), .A2(new_n719), .A3(new_n716), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n637), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT52), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n718), .A2(new_n723), .B1(new_n636), .B2(new_n635), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n675), .A2(new_n846), .A3(new_n847), .A4(new_n838), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n682), .A2(new_n685), .A3(new_n713), .A4(new_n689), .ZN(new_n850));
  INV_X1    g664(.A(new_n587), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n584), .A2(new_n469), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n610), .B2(new_n615), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n620), .A2(new_n677), .A3(new_n645), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n589), .A2(new_n627), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n749), .A2(new_n733), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n752), .A2(new_n734), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n750), .A2(new_n751), .A3(new_n717), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n445), .B(new_n667), .C1(new_n459), .C2(new_n460), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n413), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT112), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT112), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n413), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n864), .A2(new_n625), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n536), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n636), .A2(new_n868), .A3(new_n776), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n756), .A2(new_n860), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n856), .A2(new_n859), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n849), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n849), .B2(new_n871), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n756), .A2(new_n860), .A3(new_n869), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n589), .A2(new_n627), .A3(new_n854), .A4(KEYINPUT53), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n753), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n713), .A2(new_n689), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(KEYINPUT114), .A3(new_n682), .A4(new_n685), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT114), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n850), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n879), .A2(new_n848), .A3(new_n845), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n874), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n876), .A2(KEYINPUT115), .A3(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n887), .A2(KEYINPUT115), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n834), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n799), .B1(new_n890), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n188), .A2(G952), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n243), .B1(new_n874), .B2(new_n885), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(G210), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n553), .B1(new_n562), .B2(new_n564), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(new_n558), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n894), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n896), .B2(new_n899), .ZN(G51));
  NOR2_X1   g715(.A1(new_n766), .A2(new_n767), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n523), .B(KEYINPUT57), .Z(new_n904));
  AND3_X1   g718(.A1(new_n874), .A2(new_n885), .A3(new_n886), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n886), .B1(new_n874), .B2(new_n885), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n903), .B1(new_n907), .B2(new_n520), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT119), .B1(new_n908), .B2(new_n893), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n504), .A2(new_n519), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n874), .A2(new_n885), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT54), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n887), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(new_n914), .B2(new_n904), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n910), .B(new_n894), .C1(new_n915), .C2(new_n903), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n909), .A2(new_n916), .ZN(G54));
  AND2_X1   g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n895), .A2(new_n455), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n455), .B1(new_n895), .B2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n893), .ZN(G60));
  NAND2_X1  g735(.A1(new_n602), .A2(new_n604), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n606), .B(KEYINPUT59), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n914), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n894), .ZN(new_n926));
  INV_X1    g740(.A(new_n922), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n888), .A2(new_n889), .A3(new_n924), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(G63));
  XNOR2_X1  g743(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n242), .A2(new_n243), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n912), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n893), .B1(new_n933), .B2(new_n241), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT61), .B1(new_n934), .B2(KEYINPUT122), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n623), .B(KEYINPUT121), .Z(new_n936));
  NAND3_X1  g750(.A1(new_n912), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n934), .B(new_n937), .C1(KEYINPUT122), .C2(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(G66));
  OAI21_X1  g755(.A(G953), .B1(new_n464), .B2(new_n555), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n856), .B2(G953), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n897), .B1(G898), .B2(new_n188), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  AOI21_X1  g759(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n675), .A2(new_n846), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n665), .A2(KEYINPUT123), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n663), .A2(new_n664), .A3(new_n675), .A4(new_n846), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n955));
  INV_X1    g769(.A(new_n777), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT44), .B1(new_n762), .B2(new_n593), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n773), .A2(new_n646), .A3(new_n776), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n367), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n610), .A2(new_n615), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n645), .A2(new_n961), .A3(new_n646), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n960), .A2(new_n775), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT124), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n963), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n778), .A3(new_n966), .ZN(new_n967));
  AOI22_X1  g781(.A1(new_n964), .A2(new_n967), .B1(new_n788), .B2(new_n790), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n951), .A2(new_n954), .A3(new_n955), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n188), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n315), .A2(new_n316), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n449), .A2(new_n450), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n733), .A2(new_n774), .A3(new_n698), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n778), .A2(new_n756), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n977), .A2(new_n949), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n978), .A2(new_n791), .A3(new_n188), .A4(new_n859), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(G900), .B2(G953), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n979), .A2(KEYINPUT125), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT125), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n947), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n973), .B1(new_n969), .B2(new_n188), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n979), .A2(new_n980), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n947), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(KEYINPUT126), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n982), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n979), .A2(KEYINPUT125), .A3(new_n980), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n946), .B1(new_n992), .B2(new_n985), .ZN(new_n993));
  INV_X1    g807(.A(new_n988), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n989), .A2(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1001));
  INV_X1    g815(.A(new_n324), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n362), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n1000), .B(new_n1003), .C1(new_n1001), .C2(new_n362), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n875), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n978), .A2(new_n791), .A3(new_n859), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1000), .B1(new_n1006), .B2(new_n856), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n361), .A2(new_n335), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n894), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n654), .ZN(new_n1010));
  INV_X1    g824(.A(new_n856), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n999), .B1(new_n969), .B2(new_n1011), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n1005), .B(new_n1009), .C1(new_n1010), .C2(new_n1012), .ZN(G57));
endmodule


