//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  XOR2_X1   g000(.A(G110), .B(G140), .Z(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n188), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(G143), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n198), .A2(new_n199), .A3(G128), .A4(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n196), .A2(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(G128), .B1(new_n202), .B2(new_n199), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT78), .A3(G104), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n208), .B2(G104), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  OAI211_X1 g027(.A(G101), .B(new_n209), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n208), .A3(G104), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(G107), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n215), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n207), .A2(new_n221), .A3(KEYINPUT10), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT64), .B1(new_n196), .B2(G146), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n200), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n203), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n227), .A2(KEYINPUT79), .A3(new_n201), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n202), .B1(new_n195), .B2(new_n197), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n199), .A4(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n223), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(KEYINPUT79), .A3(new_n201), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n234), .A2(new_n221), .A3(KEYINPUT80), .A4(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT10), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n222), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT65), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G134), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n244), .A3(G137), .ZN(new_n245));
  NOR2_X1   g059(.A1(G134), .A2(G137), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n240), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n242), .A2(new_n244), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT11), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n239), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT65), .B(G134), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(new_n240), .A3(new_n249), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n246), .B1(new_n253), .B2(G137), .ZN(new_n255));
  OAI211_X1 g069(.A(G131), .B(new_n254), .C1(new_n255), .C2(new_n240), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n205), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(KEYINPUT0), .B(new_n260), .C1(new_n226), .C2(new_n259), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n200), .B2(new_n204), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n262), .A2(KEYINPUT0), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n215), .A2(new_n217), .A3(new_n219), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G101), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(G101), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n264), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n238), .A2(new_n258), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT82), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n207), .A2(new_n221), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n233), .B2(new_n235), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n273), .ZN(new_n277));
  INV_X1    g091(.A(new_n235), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n214), .A2(new_n220), .ZN(new_n279));
  AND4_X1   g093(.A1(new_n199), .A2(new_n198), .A3(G128), .A4(new_n200), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n280), .B2(new_n230), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT80), .B1(new_n281), .B2(new_n234), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n277), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT82), .A2(KEYINPUT12), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n258), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(KEYINPUT81), .A3(new_n257), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n276), .A2(new_n286), .B1(new_n287), .B2(KEYINPUT12), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n271), .B1(new_n288), .B2(KEYINPUT84), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT82), .B1(new_n283), .B2(KEYINPUT81), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n257), .B1(new_n274), .B2(new_n284), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n274), .A2(new_n275), .A3(new_n258), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT12), .ZN(new_n293));
  OAI22_X1  g107(.A1(new_n290), .A2(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n192), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G469), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n257), .A2(KEYINPUT83), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n238), .A2(new_n300), .A3(new_n270), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n238), .B2(new_n270), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n301), .A2(new_n302), .A3(new_n192), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n297), .A2(new_n298), .A3(new_n299), .A4(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n298), .A2(new_n299), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n192), .B1(new_n288), .B2(new_n271), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n301), .A2(new_n302), .A3(new_n191), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n306), .B1(new_n309), .B2(G469), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT9), .B(G234), .Z(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G221), .B1(new_n313), .B2(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT85), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G210), .B1(G237), .B2(G902), .ZN(new_n319));
  XOR2_X1   g133(.A(G110), .B(G122), .Z(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G116), .ZN(new_n324));
  INV_X1    g138(.A(G116), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT2), .B(G113), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n327), .B(KEYINPUT67), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n269), .A2(new_n267), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n322), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n329), .ZN(new_n334));
  XNOR2_X1  g148(.A(G116), .B(G119), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT67), .ZN(new_n336));
  INV_X1    g150(.A(new_n328), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n338), .A2(KEYINPUT86), .A3(new_n267), .A4(new_n269), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n340));
  INV_X1    g154(.A(G113), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n342), .B1(new_n330), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n334), .A3(new_n221), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n333), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n333), .A2(new_n339), .A3(new_n345), .A4(KEYINPUT87), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n321), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n350), .A2(KEYINPUT6), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n346), .A2(new_n320), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT6), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n261), .A2(G125), .A3(new_n263), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT88), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT89), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(new_n207), .B2(G125), .ZN(new_n358));
  INV_X1    g172(.A(G125), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n201), .A2(new_n206), .A3(KEYINPUT89), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G224), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G953), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n362), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(G902), .B1(new_n354), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n352), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n327), .A2(new_n343), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT90), .ZN(new_n371));
  INV_X1    g185(.A(new_n342), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n334), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n221), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n320), .B(KEYINPUT8), .Z(new_n375));
  NAND3_X1  g189(.A1(new_n344), .A2(new_n334), .A3(new_n279), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT7), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n364), .A2(KEYINPUT92), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n364), .A2(KEYINPUT92), .ZN(new_n381));
  NOR4_X1   g195(.A1(new_n362), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n361), .B(KEYINPUT91), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n383), .A2(new_n356), .B1(KEYINPUT7), .B2(new_n365), .ZN(new_n384));
  OR3_X1    g198(.A1(new_n378), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n319), .B1(new_n368), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n366), .B1(new_n351), .B2(new_n353), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n378), .A2(new_n382), .A3(new_n384), .ZN(new_n388));
  INV_X1    g202(.A(new_n319), .ZN(new_n389));
  NOR4_X1   g203(.A1(new_n387), .A2(new_n388), .A3(G902), .A4(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n318), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n315), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G475), .ZN(new_n393));
  XNOR2_X1  g207(.A(G113), .B(G122), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(new_n212), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G214), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n397), .A2(G237), .A3(G953), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT93), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G237), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n189), .A3(G214), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT93), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n196), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT94), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n398), .A2(G143), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT94), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n400), .A2(new_n403), .A3(new_n407), .A4(new_n196), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT17), .A3(G131), .ZN(new_n410));
  XNOR2_X1  g224(.A(G125), .B(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT16), .ZN(new_n412));
  OR3_X1    g226(.A1(new_n359), .A2(KEYINPUT16), .A3(G140), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n194), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(G146), .A3(new_n413), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT97), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n409), .A2(G131), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n405), .A2(new_n239), .A3(new_n406), .A4(new_n408), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n410), .A2(KEYINPUT97), .A3(new_n418), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n411), .B(G146), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT95), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n405), .A2(new_n430), .A3(new_n406), .A4(new_n408), .ZN(new_n431));
  NAND2_X1  g245(.A1(KEYINPUT18), .A2(G131), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n432), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n429), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n396), .B1(new_n428), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n429), .ZN(new_n437));
  INV_X1    g251(.A(new_n434), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n431), .A2(new_n432), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n427), .A2(new_n395), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n393), .B1(new_n442), .B2(new_n299), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT96), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n411), .B(KEYINPUT19), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n194), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n416), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n422), .B2(new_n424), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n445), .B1(new_n435), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n449), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n440), .A2(new_n451), .A3(KEYINPUT96), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n396), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(G475), .B1(new_n453), .B2(new_n441), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n299), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n455), .B1(new_n454), .B2(new_n299), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n444), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G478), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(KEYINPUT15), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT13), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n196), .A3(G128), .ZN(new_n463));
  XNOR2_X1  g277(.A(G128), .B(G143), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(G134), .B(new_n463), .C1(new_n465), .C2(new_n462), .ZN(new_n466));
  INV_X1    g280(.A(G122), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n467), .A2(KEYINPUT98), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(KEYINPUT98), .ZN(new_n469));
  OAI21_X1  g283(.A(G116), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n325), .A2(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT99), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT99), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n474), .A3(new_n471), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n473), .A2(G107), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(G107), .B1(new_n473), .B2(new_n475), .ZN(new_n477));
  OAI221_X1 g291(.A(new_n466), .B1(new_n253), .B2(new_n465), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n253), .B(new_n464), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n470), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n471), .B(KEYINPUT14), .ZN(new_n482));
  OAI21_X1  g296(.A(G107), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n480), .A2(KEYINPUT100), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT100), .B1(new_n480), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n478), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G217), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n313), .A2(new_n487), .A3(G953), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n478), .B(new_n488), .C1(new_n484), .C2(new_n485), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT101), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI211_X1 g308(.A(KEYINPUT101), .B(G902), .C1(new_n490), .C2(new_n491), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n461), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI22_X1  g310(.A1(new_n492), .A2(new_n493), .B1(KEYINPUT15), .B2(new_n460), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n189), .A2(G952), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(G234), .B2(G237), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT21), .B(G898), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(G234), .A2(G237), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(G902), .A3(G953), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n500), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n459), .A2(new_n498), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n392), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT23), .B1(new_n259), .B2(G119), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT75), .B1(new_n259), .B2(G119), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G119), .B(G128), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT24), .B(G110), .Z(new_n513));
  OAI22_X1  g327(.A1(new_n511), .A2(G110), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n411), .A2(new_n194), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n416), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT76), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(G110), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n512), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n417), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT76), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n514), .A2(new_n521), .A3(new_n416), .A4(new_n515), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT22), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(G137), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n517), .A2(new_n520), .A3(new_n522), .A4(new_n526), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n299), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n528), .A2(KEYINPUT25), .A3(new_n299), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n487), .B1(G234), .B2(new_n299), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n530), .A2(new_n535), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n250), .A2(KEYINPUT66), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n253), .A2(new_n542), .A3(new_n249), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n241), .A2(G137), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G131), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n546), .A2(new_n252), .A3(new_n207), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n252), .A2(new_n256), .B1(new_n261), .B2(new_n263), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT30), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n257), .A2(new_n264), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n546), .A2(new_n252), .A3(new_n207), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n338), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n331), .A3(new_n552), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n556));
  NAND3_X1  g370(.A1(new_n401), .A2(new_n189), .A3(G210), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT26), .B(G101), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n554), .A2(new_n555), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT31), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n547), .A2(new_n548), .A3(new_n338), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT30), .B1(new_n547), .B2(new_n548), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n551), .A2(new_n550), .A3(new_n552), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n563), .B1(new_n566), .B2(new_n338), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n560), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n331), .B1(new_n551), .B2(new_n552), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT28), .B1(new_n563), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT28), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n555), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n560), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n562), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G472), .A2(G902), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n577), .A2(KEYINPUT69), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT69), .B1(new_n577), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n540), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n582));
  AOI211_X1 g396(.A(new_n563), .B(new_n560), .C1(new_n566), .C2(new_n338), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n575), .B1(new_n571), .B2(new_n573), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT71), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n338), .B1(new_n547), .B2(new_n548), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n572), .B1(new_n587), .B2(new_n555), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT72), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n573), .B(KEYINPUT73), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n590), .A2(KEYINPUT29), .A3(new_n560), .A4(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT71), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n593), .B(new_n582), .C1(new_n583), .C2(new_n584), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n586), .A2(new_n299), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n577), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n581), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT74), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT74), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n581), .A2(new_n596), .A3(new_n600), .A4(new_n597), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n539), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n508), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  INV_X1    g418(.A(G472), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n577), .B2(new_n299), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n606), .B(KEYINPUT102), .Z(new_n607));
  OR2_X1    g421(.A1(new_n579), .A2(new_n580), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n609), .A2(new_n315), .A3(new_n539), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n350), .A2(KEYINPUT6), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n348), .A2(new_n349), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n320), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n369), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n614), .B2(KEYINPUT6), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n385), .B(new_n299), .C1(new_n615), .C2(new_n366), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n389), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n368), .A2(new_n319), .A3(new_n385), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n317), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n506), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n490), .A2(new_n491), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT33), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n490), .A2(new_n624), .A3(new_n491), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(G478), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n492), .A2(new_n460), .ZN(new_n627));
  NAND2_X1  g441(.A1(G478), .A2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n459), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n621), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n610), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  NAND2_X1  g449(.A1(new_n453), .A2(new_n441), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n393), .A3(new_n299), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT20), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n457), .A2(KEYINPUT103), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n456), .B1(new_n458), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n444), .A3(new_n498), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n621), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n610), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  INV_X1    g461(.A(new_n609), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n648), .A2(new_n392), .A3(new_n507), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n527), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT104), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n523), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n535), .A2(G902), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n534), .A2(new_n535), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT37), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G110), .ZN(G12));
  NAND2_X1  g472(.A1(new_n599), .A2(new_n601), .ZN(new_n659));
  INV_X1    g473(.A(new_n500), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n504), .A2(G900), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n643), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n659), .A2(new_n664), .A3(new_n392), .A4(new_n655), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  NAND2_X1  g480(.A1(new_n617), .A2(new_n618), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT38), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n581), .A2(new_n597), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n567), .A2(new_n575), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n587), .A2(new_n555), .A3(new_n575), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n299), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n668), .A2(new_n654), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n662), .B(KEYINPUT39), .Z(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n311), .A2(new_n314), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT40), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n459), .A2(new_n498), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n317), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n675), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n682), .B(KEYINPUT105), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n196), .ZN(G45));
  AOI21_X1  g498(.A(new_n443), .B1(new_n638), .B2(new_n456), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n685), .A2(new_n629), .A3(new_n663), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n659), .A2(new_n392), .A3(new_n655), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  NAND3_X1  g502(.A1(new_n297), .A2(new_n299), .A3(new_n304), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G469), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n690), .A2(new_n314), .A3(new_n305), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n602), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n632), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT41), .B(G113), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G15));
  NAND3_X1  g509(.A1(new_n602), .A2(new_n644), .A3(new_n691), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n602), .A2(new_n644), .A3(KEYINPUT106), .A4(new_n691), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n690), .A2(new_n314), .A3(new_n305), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(new_n391), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n294), .A2(new_n295), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n287), .A2(KEYINPUT12), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n706), .B(KEYINPUT84), .C1(new_n290), .C2(new_n291), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n707), .A3(new_n271), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n303), .B1(new_n708), .B2(new_n192), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n298), .B1(new_n709), .B2(new_n299), .ZN(new_n710));
  INV_X1    g524(.A(new_n271), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n294), .B2(new_n295), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n191), .B1(new_n712), .B2(new_n707), .ZN(new_n713));
  NOR4_X1   g527(.A1(new_n713), .A2(G469), .A3(G902), .A4(new_n303), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(KEYINPUT107), .A3(new_n314), .A4(new_n619), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n704), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n654), .B1(new_n599), .B2(new_n601), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n507), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  NOR3_X1   g534(.A1(new_n703), .A2(new_n391), .A3(new_n680), .ZN(new_n721));
  INV_X1    g535(.A(new_n578), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n562), .A2(new_n569), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n571), .A2(new_n589), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n588), .A2(KEYINPUT72), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n591), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n575), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n722), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n539), .A2(new_n606), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n721), .A2(new_n620), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n728), .A2(new_n606), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(new_n655), .ZN(new_n734));
  NOR4_X1   g548(.A1(new_n728), .A2(new_n606), .A3(new_n654), .A4(KEYINPUT108), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n686), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT107), .B1(new_n691), .B2(new_n619), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n703), .A2(new_n391), .A3(new_n702), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n717), .A2(KEYINPUT109), .A3(new_n737), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT110), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n359), .ZN(G27));
  NAND2_X1  g560(.A1(new_n577), .A2(new_n578), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT32), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT112), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n539), .B1(new_n749), .B2(new_n596), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n667), .A2(new_n317), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n314), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n308), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n308), .A2(new_n753), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n307), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n306), .B1(new_n756), .B2(G469), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n305), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n752), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n750), .A2(new_n760), .A3(new_n686), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n760), .A2(new_n763), .A3(new_n602), .A4(new_n686), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n239), .ZN(G33));
  NAND3_X1  g580(.A1(new_n760), .A2(new_n602), .A3(new_n664), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  NAND2_X1  g582(.A1(new_n630), .A2(new_n685), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT114), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n629), .B(KEYINPUT113), .Z(new_n773));
  OAI21_X1  g587(.A(new_n770), .B1(new_n773), .B2(new_n459), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n609), .A3(new_n655), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n609), .A4(new_n655), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n751), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT115), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n756), .A2(KEYINPUT45), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n309), .A2(KEYINPUT45), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(G469), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n306), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n714), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n785), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n314), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n676), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n778), .A2(new_n792), .A3(new_n751), .A4(new_n779), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n781), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  AND3_X1   g609(.A1(new_n789), .A2(KEYINPUT47), .A3(new_n314), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT47), .B1(new_n789), .B2(new_n314), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n686), .B(new_n751), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n659), .A3(new_n538), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT116), .Z(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  XOR2_X1   g615(.A(new_n715), .B(KEYINPUT49), .Z(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n317), .A3(new_n668), .ZN(new_n803));
  INV_X1    g617(.A(new_n769), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n674), .A2(new_n539), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n314), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n796), .A2(new_n797), .ZN(new_n807));
  INV_X1    g621(.A(new_n715), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n314), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n660), .B1(new_n772), .B2(new_n774), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(new_n729), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n751), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(KEYINPUT121), .A3(new_n751), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n809), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n752), .A2(new_n660), .A3(new_n808), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n685), .A3(new_n629), .A4(new_n805), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n775), .B(new_n817), .C1(new_n735), .C2(new_n734), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT122), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n668), .A2(new_n318), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n810), .A2(new_n691), .A3(new_n729), .A4(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT50), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n816), .A2(new_n818), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n827), .A2(new_n828), .A3(new_n499), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n775), .A2(new_n750), .A3(new_n817), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT48), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n811), .A2(new_n717), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n817), .A2(new_n459), .A3(new_n630), .A4(new_n805), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n829), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n665), .A2(new_n687), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n742), .B2(new_n743), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n681), .A2(new_n667), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n759), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n655), .B1(new_n669), .B2(new_n673), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n840), .A3(new_n314), .A4(new_n662), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT117), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n718), .B(new_n392), .C1(new_n664), .C2(new_n686), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT109), .B1(new_n717), .B2(new_n737), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n741), .B(new_n736), .C1(new_n704), .C2(new_n716), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n843), .B(new_n841), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n835), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n719), .A2(new_n730), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n692), .A2(new_n632), .B1(new_n602), .B2(new_n508), .ZN(new_n851));
  INV_X1    g665(.A(new_n498), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n631), .B1(new_n459), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n853), .A2(new_n619), .A3(new_n620), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n649), .A2(new_n655), .B1(new_n610), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n850), .A2(new_n700), .A3(new_n851), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n718), .A2(new_n311), .A3(new_n852), .A4(new_n662), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n642), .A2(new_n444), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n857), .A2(new_n858), .B1(new_n736), .B2(new_n759), .ZN(new_n859));
  INV_X1    g673(.A(new_n752), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n762), .A2(new_n764), .A3(new_n767), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n856), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n846), .A2(new_n847), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n744), .A2(KEYINPUT117), .A3(new_n843), .A4(new_n841), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT52), .ZN(new_n867));
  AND4_X1   g681(.A1(KEYINPUT53), .A2(new_n849), .A3(new_n864), .A4(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(KEYINPUT118), .B(KEYINPUT52), .Z(new_n869));
  NAND3_X1  g683(.A1(new_n865), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n837), .A2(KEYINPUT52), .A3(new_n841), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT53), .B1(new_n872), .B2(new_n864), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT54), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(KEYINPUT53), .A3(new_n864), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT52), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(new_n865), .B2(new_n866), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n698), .A2(new_n699), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n854), .A2(new_n610), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n656), .A2(new_n719), .A3(new_n730), .A4(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n863), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n861), .A4(new_n851), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n877), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n875), .B(new_n876), .C1(new_n885), .C2(KEYINPUT53), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n874), .A2(KEYINPUT119), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n849), .A2(new_n864), .A3(new_n867), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n891), .A3(new_n875), .A4(new_n876), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT120), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n895), .A3(new_n892), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n834), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(G952), .A2(G953), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n806), .B1(new_n897), .B2(new_n898), .ZN(G75));
  AOI21_X1  g713(.A(new_n299), .B1(new_n890), .B2(new_n876), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G210), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n354), .A2(new_n367), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n387), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n901), .B2(new_n902), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n189), .A2(G952), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT123), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(G51));
  NAND2_X1  g725(.A1(new_n785), .A2(KEYINPUT57), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n785), .A2(KEYINPUT57), .ZN(new_n913));
  INV_X1    g727(.A(new_n886), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n875), .B1(new_n890), .B2(new_n876), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n912), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n709), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n900), .A2(G469), .A3(new_n783), .A4(new_n782), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n910), .B1(new_n917), .B2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n900), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n920), .A2(new_n636), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n636), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n910), .B1(new_n921), .B2(new_n922), .ZN(G60));
  NAND2_X1  g737(.A1(new_n623), .A2(new_n625), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n628), .B(KEYINPUT59), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n924), .B(new_n925), .C1(new_n914), .C2(new_n915), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n909), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n894), .A2(new_n896), .A3(new_n925), .ZN(new_n928));
  INV_X1    g742(.A(new_n924), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n890), .B2(new_n876), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n910), .B1(new_n933), .B2(new_n652), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n528), .A2(new_n529), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n936), .B2(new_n933), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g752(.A(G953), .B1(new_n502), .B2(new_n363), .ZN(new_n939));
  INV_X1    g753(.A(new_n856), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n615), .B1(G898), .B2(new_n189), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT124), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  OR2_X1    g758(.A1(new_n853), .A2(KEYINPUT125), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n678), .B1(new_n853), .B2(KEYINPUT125), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n945), .A2(new_n946), .A3(new_n602), .A4(new_n751), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(KEYINPUT126), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(KEYINPUT126), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n800), .A2(new_n794), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n683), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n837), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n189), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n566), .B(new_n446), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(G900), .A2(G953), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n790), .A2(new_n676), .A3(new_n838), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n863), .B1(new_n750), .B2(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n794), .A2(KEYINPUT127), .A3(new_n837), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT127), .B1(new_n794), .B2(new_n837), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n800), .B(new_n960), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n955), .B(new_n958), .C1(new_n963), .C2(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n966), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n957), .A2(new_n968), .A3(new_n964), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(G72));
  NOR3_X1   g784(.A1(new_n950), .A2(new_n953), .A3(new_n856), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n670), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n963), .B2(new_n856), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n910), .B1(new_n976), .B2(new_n583), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n670), .A2(new_n583), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n973), .B(new_n978), .C1(new_n868), .C2(new_n873), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n975), .A2(new_n977), .A3(new_n979), .ZN(G57));
endmodule


