//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n213));
  XNOR2_X1  g0013(.A(new_n212), .B(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n203), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n222), .B1(new_n201), .B2(new_n223), .C1(new_n202), .C2(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n221), .B(new_n225), .C1(G107), .C2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT66), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(G77), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n226), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(new_n210), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n214), .B(new_n219), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n224), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND3_X1  g0049(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n203), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT12), .B1(new_n252), .B2(KEYINPUT73), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(KEYINPUT73), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n250), .A2(new_n217), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n207), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G68), .A3(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n262));
  INV_X1    g0062(.A(G77), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n208), .A2(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(new_n217), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n267), .A2(KEYINPUT11), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(KEYINPUT11), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n255), .B(new_n260), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  OAI211_X1 g0072(.A(G232), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n276), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G97), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(G226), .A3(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n275), .A2(new_n277), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  OR2_X1    g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n284), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n286), .B1(new_n289), .B2(new_n220), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT13), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT13), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n283), .A2(new_n294), .A3(new_n291), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT75), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT74), .B(KEYINPUT14), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n296), .A2(new_n297), .A3(G169), .A4(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n294), .B1(new_n283), .B2(new_n291), .ZN(new_n300));
  AOI211_X1 g0100(.A(KEYINPUT13), .B(new_n290), .C1(new_n281), .C2(new_n282), .ZN(new_n301));
  OAI211_X1 g0101(.A(G169), .B(new_n298), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT75), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(G169), .B1(new_n300), .B2(new_n301), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT14), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n295), .A2(KEYINPUT72), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT72), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n283), .A2(new_n308), .A3(new_n294), .A4(new_n291), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n307), .A2(new_n293), .A3(G179), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n270), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n286), .B1(new_n289), .B2(new_n229), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n276), .A2(G232), .A3(new_n279), .ZN(new_n314));
  INV_X1    g0114(.A(G107), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n276), .A2(G1698), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n314), .B1(new_n315), .B2(new_n276), .C1(new_n316), .C2(new_n220), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n313), .B1(new_n317), .B2(new_n282), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n258), .A2(G77), .A3(new_n259), .ZN(new_n322));
  XOR2_X1   g0122(.A(new_n322), .B(KEYINPUT68), .Z(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(G20), .ZN(new_n327));
  XOR2_X1   g0127(.A(KEYINPUT8), .B(G58), .Z(new_n328));
  AOI22_X1  g0128(.A1(new_n325), .A2(new_n327), .B1(new_n328), .B2(new_n261), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n208), .B2(new_n230), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n266), .B1(new_n230), .B2(new_n251), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n318), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n321), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n323), .B(new_n331), .C1(new_n318), .C2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT69), .ZN(new_n338));
  INV_X1    g0138(.A(G190), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n337), .A2(new_n338), .B1(new_n339), .B2(new_n319), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n323), .A2(new_n331), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n319), .A2(G200), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT69), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n335), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n328), .A2(new_n259), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n345), .A2(new_n257), .B1(new_n250), .B2(new_n328), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT7), .B1(new_n276), .B2(G20), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n271), .A2(new_n272), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(new_n208), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n350), .A3(G68), .ZN(new_n351));
  XNOR2_X1  g0151(.A(G58), .B(G68), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(G20), .B1(G159), .B2(new_n261), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT16), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n266), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(KEYINPUT16), .A3(new_n353), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n346), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n286), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n223), .A2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G223), .B2(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G87), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n361), .A2(new_n348), .B1(new_n326), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n359), .B1(new_n363), .B2(new_n282), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n288), .A2(G232), .A3(new_n284), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT76), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n336), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n364), .A2(new_n367), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(G190), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n358), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n356), .A2(new_n357), .ZN(new_n374));
  INV_X1    g0174(.A(new_n346), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n364), .A2(new_n367), .A3(G179), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n320), .B1(new_n364), .B2(new_n367), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT18), .B1(new_n358), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n358), .A2(new_n370), .A3(KEYINPUT17), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n373), .A2(new_n381), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n344), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n286), .B1(new_n289), .B2(new_n223), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n276), .A2(G222), .A3(new_n279), .ZN(new_n388));
  INV_X1    g0188(.A(G223), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n388), .B1(new_n230), .B2(new_n276), .C1(new_n316), .C2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n390), .B2(new_n282), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(G179), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n328), .A2(new_n327), .B1(G150), .B2(new_n261), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(KEYINPUT67), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n394), .A2(KEYINPUT67), .B1(G20), .B2(new_n204), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n355), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n259), .A2(G50), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n257), .A2(new_n398), .B1(G50), .B2(new_n250), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n391), .A2(G169), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n393), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT70), .B1(new_n392), .B2(new_n339), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT70), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n391), .A2(new_n404), .A3(G190), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n399), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n395), .A2(new_n396), .ZN(new_n408));
  OAI211_X1 g0208(.A(KEYINPUT9), .B(new_n407), .C1(new_n408), .C2(new_n355), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT9), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n397), .B2(new_n399), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n392), .A2(G200), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT10), .B1(new_n406), .B2(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n411), .A2(new_n412), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n403), .A2(new_n405), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT10), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .A4(new_n409), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n402), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n270), .B1(new_n296), .B2(G200), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n307), .A2(new_n293), .A3(G190), .A4(new_n309), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AND4_X1   g0222(.A1(new_n312), .A2(new_n386), .A3(new_n419), .A4(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT5), .B(G41), .ZN(new_n424));
  INV_X1    g0224(.A(G45), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(G1), .ZN(new_n426));
  INV_X1    g0226(.A(new_n217), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n424), .A2(new_n426), .B1(new_n427), .B2(new_n287), .ZN(new_n428));
  NAND2_X1  g0228(.A1(KEYINPUT5), .A2(G41), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(KEYINPUT5), .A2(G41), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n285), .B1(new_n427), .B2(new_n287), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n428), .A2(G270), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(G264), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n436));
  INV_X1    g0236(.A(new_n272), .ZN(new_n437));
  NAND2_X1  g0237(.A1(KEYINPUT3), .A2(G33), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(G303), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(G257), .B(new_n279), .C1(new_n271), .C2(new_n272), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n436), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n282), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT77), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n326), .B2(G1), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n207), .A2(KEYINPUT77), .A3(G33), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n258), .A2(new_n447), .A3(G116), .ZN(new_n448));
  INV_X1    g0248(.A(G116), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n251), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n256), .A2(new_n217), .B1(G20), .B2(new_n449), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  INV_X1    g0252(.A(G97), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n208), .C1(G33), .C2(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n451), .A2(KEYINPUT20), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT20), .B1(new_n451), .B2(new_n454), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n448), .B(new_n450), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n443), .A2(new_n457), .A3(KEYINPUT21), .A4(G169), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n320), .B1(new_n435), .B2(new_n442), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n461), .A2(KEYINPUT79), .A3(KEYINPUT21), .A4(new_n457), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n457), .B1(new_n443), .B2(G200), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n339), .B2(new_n443), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n457), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT21), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n435), .A2(G179), .A3(new_n442), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n466), .A2(new_n467), .B1(new_n468), .B2(new_n457), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n463), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT80), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n327), .A2(G116), .ZN(new_n474));
  OR3_X1    g0274(.A1(new_n208), .A2(KEYINPUT23), .A3(G107), .ZN(new_n475));
  OAI211_X1 g0275(.A(KEYINPUT80), .B(KEYINPUT23), .C1(new_n208), .C2(G107), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n473), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n208), .B(G87), .C1(new_n271), .C2(new_n272), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT22), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT22), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n276), .A2(new_n481), .A3(new_n208), .A4(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT24), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n355), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n477), .B1(new_n480), .B2(new_n482), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT24), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n207), .A2(new_n315), .A3(G13), .A4(G20), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT25), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n258), .A2(new_n447), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n489), .B(new_n492), .C1(new_n493), .C2(new_n315), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n445), .A2(new_n446), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n257), .A2(new_n495), .A3(new_n315), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n490), .B(KEYINPUT25), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT81), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n486), .A2(new_n488), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  OAI211_X1 g0300(.A(G250), .B(new_n279), .C1(new_n271), .C2(new_n272), .ZN(new_n501));
  OAI211_X1 g0301(.A(G257), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G294), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n282), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n424), .A2(new_n288), .A3(G274), .A4(new_n426), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n428), .A2(G264), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n320), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n504), .A2(new_n282), .B1(new_n428), .B2(G264), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n333), .A3(new_n506), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n499), .A2(new_n500), .A3(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n509), .A2(new_n511), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n498), .A2(new_n494), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n266), .B1(new_n487), .B2(KEYINPUT24), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n484), .A2(new_n485), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT82), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  AND2_X1   g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G97), .A2(G107), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n315), .A2(KEYINPUT6), .A3(G97), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n347), .A2(new_n350), .A3(G107), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n266), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n251), .A2(new_n453), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n493), .B2(new_n453), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n432), .A2(new_n288), .ZN(new_n534));
  INV_X1    g0334(.A(G257), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n506), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(G244), .B(new_n279), .C1(new_n271), .C2(new_n272), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n276), .A2(KEYINPUT4), .A3(G244), .A4(new_n279), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n452), .A4(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n536), .B1(new_n542), .B2(new_n282), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n530), .B(new_n533), .C1(new_n543), .C2(new_n336), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n282), .ZN(new_n545));
  INV_X1    g0345(.A(new_n536), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(new_n339), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n355), .B1(new_n527), .B2(new_n528), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n543), .A2(G169), .B1(new_n549), .B2(new_n532), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n545), .A2(new_n333), .A3(new_n546), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n544), .A2(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n508), .A2(G200), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n510), .A2(G190), .A3(new_n506), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n518), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n208), .B1(new_n278), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n523), .A2(new_n362), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n208), .B(G68), .C1(new_n271), .C2(new_n272), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n557), .B1(new_n264), .B2(new_n453), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n266), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n324), .A2(new_n251), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n258), .A2(new_n447), .A3(G87), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(G238), .B(new_n279), .C1(new_n271), .C2(new_n272), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G116), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n282), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n426), .A2(G274), .ZN(new_n574));
  OAI21_X1  g0374(.A(G250), .B1(new_n425), .B2(G1), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n282), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G200), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n576), .B1(new_n572), .B2(new_n282), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n568), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n258), .A2(new_n447), .A3(new_n325), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n564), .A2(new_n565), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n563), .A2(new_n266), .B1(new_n251), .B2(new_n324), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT78), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n583), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n580), .A2(new_n320), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n333), .B(new_n576), .C1(new_n572), .C2(new_n282), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n582), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n552), .A2(new_n556), .A3(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n423), .A2(new_n470), .A3(new_n520), .A4(new_n594), .ZN(new_n595));
  XOR2_X1   g0395(.A(new_n595), .B(KEYINPUT83), .Z(G372));
  NAND2_X1  g0396(.A1(new_n414), .A2(new_n418), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n373), .A2(new_n384), .ZN(new_n598));
  INV_X1    g0398(.A(new_n335), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n422), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n598), .B1(new_n312), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n381), .A2(new_n383), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n402), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n578), .A2(G169), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n580), .A2(G179), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n607), .A2(new_n608), .B1(new_n586), .B2(new_n583), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n320), .B2(new_n580), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n585), .A3(new_n588), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n547), .A2(new_n320), .B1(new_n530), .B2(new_n533), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n543), .A2(new_n333), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .A4(new_n582), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n609), .B1(new_n614), .B2(KEYINPUT26), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n586), .B(new_n566), .C1(new_n580), .C2(new_n336), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n616), .A2(new_n617), .B1(G190), .B2(new_n580), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n568), .A2(new_n579), .A3(KEYINPUT84), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n609), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n530), .A2(new_n533), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n621), .B(new_n613), .C1(G169), .C2(new_n543), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n486), .A2(new_n488), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(new_n515), .A3(new_n554), .A4(new_n553), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n543), .A2(G190), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n549), .A2(new_n532), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n628), .B(new_n629), .C1(new_n336), .C2(new_n543), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n620), .A2(new_n627), .A3(new_n622), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n514), .A2(new_n518), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n632), .A2(new_n463), .A3(new_n469), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n615), .B(new_n625), .C1(new_n631), .C2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n423), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n606), .A2(new_n635), .ZN(G369));
  NAND2_X1  g0436(.A1(new_n463), .A2(new_n469), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n457), .A2(new_n643), .ZN(new_n644));
  MUX2_X1   g0444(.A(new_n637), .B(new_n470), .S(new_n644), .Z(new_n645));
  XNOR2_X1  g0445(.A(KEYINPUT85), .B(G330), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n556), .B1(new_n518), .B2(new_n643), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n520), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n643), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n632), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n637), .A2(new_n651), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n520), .A3(new_n649), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n514), .A2(new_n518), .A3(new_n651), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(G399));
  INV_X1    g0459(.A(new_n211), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(G41), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n559), .A2(G116), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G1), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n215), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT29), .B1(new_n634), .B2(new_n651), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n627), .A2(new_n622), .A3(new_n630), .ZN(new_n668));
  INV_X1    g0468(.A(new_n609), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n580), .A2(new_n336), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n617), .B1(new_n670), .B2(new_n567), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n581), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n616), .A2(new_n617), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n500), .B1(new_n499), .B2(new_n512), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n514), .A2(new_n518), .A3(KEYINPUT82), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(new_n463), .A4(new_n469), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n609), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n624), .B1(new_n593), .B2(new_n622), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT88), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n620), .A2(new_n623), .A3(KEYINPUT26), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n614), .A2(KEYINPUT88), .A3(new_n624), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n643), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n667), .B1(KEYINPUT29), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n578), .A2(KEYINPUT86), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT86), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n580), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n547), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n443), .A2(new_n508), .A3(new_n333), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT87), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n443), .A2(new_n508), .A3(new_n333), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n545), .A2(new_n546), .B1(new_n578), .B2(KEYINPUT86), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT87), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .A4(new_n691), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n510), .A2(new_n580), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n468), .A3(new_n543), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n699), .A2(new_n468), .A3(KEYINPUT30), .A4(new_n543), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n694), .A2(new_n698), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n643), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n594), .A2(new_n520), .A3(new_n470), .A4(new_n651), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n706), .B1(new_n707), .B2(KEYINPUT31), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n702), .B(new_n703), .C1(new_n693), .C2(new_n692), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n646), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n688), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n666), .B1(new_n713), .B2(G1), .ZN(G364));
  NOR2_X1   g0514(.A1(new_n645), .A2(new_n646), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n208), .A2(G13), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n207), .B1(new_n716), .B2(G45), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n715), .B(new_n648), .C1(new_n662), .C2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n717), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n661), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n211), .A2(new_n276), .ZN(new_n721));
  INV_X1    g0521(.A(G355), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n721), .A2(new_n722), .B1(G116), .B2(new_n211), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n660), .A2(new_n276), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n425), .B2(new_n216), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n245), .A2(new_n425), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n208), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT89), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n217), .B1(G20), .B2(new_n320), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n720), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n208), .A2(new_n339), .A3(new_n336), .A4(G179), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n362), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n208), .A2(new_n333), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G190), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n740), .A2(new_n339), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n742), .A2(new_n203), .B1(new_n744), .B2(new_n201), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n208), .B1(new_n746), .B2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n738), .B(new_n745), .C1(G97), .C2(new_n748), .ZN(new_n749));
  NOR4_X1   g0549(.A1(new_n208), .A2(new_n336), .A3(G179), .A4(G190), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n276), .B1(new_n751), .B2(new_n315), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n746), .A2(G20), .A3(new_n339), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(KEYINPUT32), .A3(G159), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT32), .ZN(new_n756));
  INV_X1    g0556(.A(G159), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n756), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n752), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n739), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT90), .ZN(new_n761));
  AOI21_X1  g0561(.A(G200), .B1(new_n760), .B2(KEYINPUT90), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n761), .A2(G190), .A3(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n749), .B(new_n759), .C1(new_n202), .C2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n761), .A2(new_n339), .A3(new_n762), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT91), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT91), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n230), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n743), .A2(G326), .ZN(new_n773));
  INV_X1    g0573(.A(G303), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n774), .B2(new_n737), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G283), .B2(new_n750), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n742), .B1(new_n777), .B2(KEYINPUT92), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(KEYINPUT92), .B2(new_n777), .ZN(new_n779));
  INV_X1    g0579(.A(new_n763), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G322), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n747), .A2(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n276), .B(new_n783), .C1(G329), .C2(new_n754), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n776), .A2(new_n779), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n764), .A2(new_n770), .B1(new_n772), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n735), .B1(new_n786), .B2(new_n732), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n731), .B(KEYINPUT93), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n645), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT94), .Z(new_n791));
  NOR2_X1   g0591(.A1(new_n718), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  NAND2_X1  g0593(.A1(new_n634), .A2(new_n651), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n335), .A2(new_n643), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n340), .A2(new_n343), .B1(new_n341), .B2(new_n651), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n335), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n797), .A2(new_n634), .A3(new_n651), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(new_n711), .ZN(new_n802));
  INV_X1    g0602(.A(new_n720), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n805), .A2(KEYINPUT96), .B1(new_n711), .B2(new_n801), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(KEYINPUT96), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n732), .A2(new_n729), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n720), .B1(G77), .B2(new_n809), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n348), .B1(new_n753), .B2(new_n771), .C1(new_n453), .C2(new_n747), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n736), .A2(G107), .B1(new_n750), .B2(G87), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n744), .B2(new_n774), .C1(new_n813), .C2(new_n742), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n811), .B(new_n814), .C1(G294), .C2(new_n780), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n449), .B2(new_n769), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n741), .A2(G150), .B1(new_n743), .B2(G137), .ZN(new_n817));
  INV_X1    g0617(.A(G143), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n817), .B1(new_n818), .B2(new_n763), .C1(new_n769), .C2(new_n757), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT95), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(KEYINPUT34), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n276), .B1(new_n753), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G58), .B2(new_n748), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n736), .A2(G50), .B1(new_n750), .B2(G68), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n820), .A2(KEYINPUT34), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n816), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n810), .B1(new_n828), .B2(new_n732), .ZN(new_n829));
  INV_X1    g0629(.A(new_n729), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n830), .B2(new_n797), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n807), .A2(new_n831), .ZN(G384));
  OR2_X1    g0632(.A1(new_n526), .A2(KEYINPUT35), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n526), .A2(KEYINPUT35), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n833), .A2(new_n834), .A3(G116), .A4(new_n218), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT36), .Z(new_n836));
  AOI21_X1  g0636(.A(new_n230), .B1(G58), .B2(G68), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n216), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n201), .A2(G68), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n207), .B(G13), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT103), .B1(new_n687), .B2(new_n423), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n679), .A2(new_n685), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n843), .A2(KEYINPUT29), .A3(new_n651), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT29), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n794), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g0646(.A1(KEYINPUT103), .A2(new_n423), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n606), .B1(new_n842), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT104), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n376), .A2(new_n380), .ZN(new_n850));
  INV_X1    g0650(.A(new_n641), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n376), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT37), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n850), .A2(new_n852), .A3(new_n853), .A4(new_n371), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n354), .A2(KEYINPUT99), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n351), .A2(new_n353), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT99), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(KEYINPUT16), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n266), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n375), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n851), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n380), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n861), .A2(new_n862), .A3(new_n371), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n854), .B1(new_n863), .B2(new_n853), .ZN(new_n864));
  INV_X1    g0664(.A(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n385), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT100), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n864), .A2(new_n866), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n864), .A2(KEYINPUT100), .A3(new_n866), .A4(KEYINPUT38), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n869), .A2(new_n872), .A3(KEYINPUT39), .A4(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n875));
  INV_X1    g0675(.A(new_n852), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n385), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n385), .A2(KEYINPUT102), .A3(new_n876), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n850), .A2(new_n852), .A3(new_n371), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n854), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n875), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n874), .B1(new_n886), .B2(KEYINPUT39), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n312), .A2(KEYINPUT97), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n299), .A2(new_n303), .A3(new_n306), .A4(new_n310), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT97), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n890), .A3(new_n270), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n643), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n795), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n800), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n889), .A2(new_n890), .A3(new_n270), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n890), .B1(new_n889), .B2(new_n270), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n270), .A2(new_n643), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n422), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n899), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n889), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT98), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n900), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n888), .A2(new_n891), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT98), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n908), .A3(new_n903), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n896), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n869), .A2(new_n873), .A3(new_n872), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n602), .A2(new_n641), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n894), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n849), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n707), .A2(KEYINPUT31), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT106), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT106), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n704), .A2(new_n920), .A3(KEYINPUT31), .A4(new_n643), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n917), .A2(new_n705), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(new_n798), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n907), .A2(new_n908), .A3(new_n903), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n908), .B1(new_n907), .B2(new_n903), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(new_n911), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n919), .A2(new_n921), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n797), .B1(new_n928), .B2(new_n708), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n905), .B2(new_n909), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT40), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n886), .A2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n926), .A2(new_n927), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n386), .A2(new_n419), .A3(new_n312), .A4(new_n422), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(new_n922), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n933), .B(new_n423), .C1(new_n708), .C2(new_n928), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n646), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n916), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n207), .B2(new_n716), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n916), .A2(new_n938), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n841), .B1(new_n940), .B2(new_n941), .ZN(G367));
  OAI211_X1 g0742(.A(new_n622), .B(new_n630), .C1(new_n629), .C2(new_n651), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n623), .A2(new_n643), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n656), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT42), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n943), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT107), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n519), .B2(new_n513), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n643), .B1(new_n949), .B2(new_n622), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT43), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n568), .A2(new_n651), .ZN(new_n952));
  MUX2_X1   g0752(.A(new_n674), .B(new_n669), .S(new_n952), .Z(new_n953));
  OAI22_X1  g0753(.A1(new_n946), .A2(new_n950), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n951), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n954), .B(new_n955), .Z(new_n956));
  INV_X1    g0756(.A(new_n948), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n653), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n956), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n956), .B2(new_n959), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n658), .A2(new_n947), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT45), .Z(new_n965));
  NOR2_X1   g0765(.A1(new_n658), .A2(new_n947), .ZN(new_n966));
  XNOR2_X1  g0766(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(new_n653), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n656), .B1(new_n652), .B2(new_n655), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n648), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n712), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n661), .B(KEYINPUT41), .Z(new_n974));
  OAI21_X1  g0774(.A(new_n717), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n953), .A2(new_n788), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n725), .A2(new_n241), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n733), .B1(new_n211), .B2(new_n324), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n720), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n744), .A2(new_n818), .B1(new_n202), .B2(new_n737), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n742), .A2(new_n757), .B1(new_n230), .B2(new_n751), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n348), .B1(new_n754), .B2(G137), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n203), .B2(new_n747), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(G150), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(new_n985), .B2(new_n763), .C1(new_n769), .C2(new_n201), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n736), .A2(G116), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT46), .Z(new_n988));
  INV_X1    g0788(.A(G317), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n348), .B1(new_n753), .B2(new_n989), .C1(new_n315), .C2(new_n747), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n742), .A2(new_n782), .B1(new_n453), .B2(new_n751), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n769), .B2(new_n813), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n763), .A2(new_n774), .B1(new_n771), .B2(new_n744), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT110), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n986), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n979), .B1(new_n997), .B2(new_n732), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n963), .A2(new_n975), .B1(new_n976), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(G387));
  NOR2_X1   g0800(.A1(new_n652), .A2(new_n789), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n238), .A2(G45), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT111), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n328), .A2(new_n201), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT50), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n663), .B(new_n425), .C1(new_n203), .C2(new_n263), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1003), .B(new_n724), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(G107), .B2(new_n211), .C1(new_n663), .C2(new_n721), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n733), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n720), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n276), .B1(new_n751), .B2(new_n453), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n741), .A2(new_n328), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n324), .B2(new_n747), .C1(new_n744), .C2(new_n757), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(G50), .C2(new_n780), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n737), .A2(new_n230), .B1(new_n985), .B2(new_n753), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT112), .Z(new_n1016));
  OAI211_X1 g0816(.A(new_n1014), .B(new_n1016), .C1(new_n203), .C2(new_n769), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n276), .B1(new_n754), .B2(G326), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n737), .A2(new_n782), .B1(new_n813), .B2(new_n747), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n741), .A2(G311), .B1(new_n743), .B2(G322), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n989), .B2(new_n763), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n768), .B2(G303), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1019), .B1(new_n1022), .B2(KEYINPUT48), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(KEYINPUT48), .B2(new_n1022), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT49), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1018), .B1(new_n449), .B2(new_n751), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1017), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1001), .B(new_n1010), .C1(new_n732), .C2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n972), .B2(new_n719), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n713), .A2(new_n972), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n661), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n713), .A2(new_n972), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(G393));
  INV_X1    g0834(.A(new_n1031), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n662), .B1(new_n970), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n970), .B2(new_n1035), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n734), .B1(G97), .B2(new_n660), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n724), .A2(new_n248), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n803), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n763), .A2(new_n757), .B1(new_n985), .B2(new_n744), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT51), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n736), .A2(G68), .B1(new_n754), .B2(G143), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n348), .B1(new_n750), .B2(G87), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n741), .A2(G50), .B1(G77), .B2(new_n748), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1044), .B(new_n1048), .C1(new_n768), .C2(new_n328), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n276), .B1(new_n754), .B2(G322), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n315), .B2(new_n751), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n741), .A2(G303), .B1(G116), .B2(new_n748), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n813), .B2(new_n737), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1051), .B(new_n1053), .C1(new_n768), .C2(G294), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n763), .A2(new_n771), .B1(new_n989), .B2(new_n744), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT52), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1042), .A2(new_n1049), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n732), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1040), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n957), .B2(new_n731), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n970), .B2(new_n719), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1037), .A2(new_n1061), .ZN(G390));
  INV_X1    g0862(.A(G330), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n917), .A2(new_n705), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n919), .A2(new_n921), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n797), .B(new_n1066), .C1(new_n924), .C2(new_n925), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n887), .B1(new_n910), .B2(new_n892), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n796), .A2(new_n335), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n686), .A2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n924), .A2(new_n925), .B1(new_n1070), .B2(new_n795), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n886), .A2(new_n892), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1067), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n896), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n924), .B2(new_n925), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n893), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1077), .A2(new_n887), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n646), .B(new_n797), .C1(new_n708), .C2(new_n710), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n924), .B2(new_n925), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1074), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g0882(.A1(new_n922), .A2(new_n1063), .A3(new_n935), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n606), .B(new_n1084), .C1(new_n842), .C2(new_n847), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n905), .A2(new_n909), .A3(new_n1079), .ZN(new_n1086));
  OAI211_X1 g0886(.A(G330), .B(new_n797), .C1(new_n928), .C2(new_n708), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n905), .B2(new_n909), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1075), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1070), .A2(new_n795), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n905), .A2(new_n1087), .A3(new_n909), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1081), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(KEYINPUT114), .B(new_n1085), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT114), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n423), .A2(new_n844), .A3(new_n846), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT103), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n423), .A2(new_n844), .A3(new_n846), .A4(KEYINPUT103), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n605), .B(new_n1083), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1094), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1082), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1081), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n905), .A2(new_n909), .A3(new_n1079), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n896), .B1(new_n1067), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1100), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(KEYINPUT114), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1068), .A2(new_n1073), .A3(new_n1081), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1078), .B2(new_n1067), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1095), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1102), .A2(new_n661), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n887), .A2(new_n729), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n720), .B1(new_n328), .B2(new_n809), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n769), .A2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n741), .A2(G137), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n348), .B(new_n1117), .C1(G125), .C2(new_n754), .ZN(new_n1118));
  INV_X1    g0918(.A(G128), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n744), .A2(new_n1119), .B1(new_n747), .B2(new_n757), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(G50), .B2(new_n750), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n780), .A2(G132), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n736), .A2(G150), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT53), .Z(new_n1124));
  NAND4_X1  g0924(.A1(new_n1118), .A2(new_n1121), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n769), .A2(new_n453), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n276), .B(new_n738), .C1(G294), .C2(new_n754), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n741), .A2(G107), .B1(new_n743), .B2(G283), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n780), .A2(G116), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n748), .A2(G77), .B1(new_n750), .B2(G68), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1116), .A2(new_n1125), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1114), .B1(new_n1132), .B2(new_n732), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1082), .A2(new_n719), .B1(new_n1113), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1112), .A2(new_n1134), .ZN(G378));
  NAND2_X1  g0935(.A1(new_n926), .A2(new_n927), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n930), .A2(new_n932), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1136), .A2(KEYINPUT117), .A3(new_n1137), .A4(G330), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n400), .A2(new_n641), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT55), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n419), .B(new_n1140), .ZN(new_n1141));
  XOR2_X1   g0941(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n1142));
  XOR2_X1   g0942(.A(new_n1141), .B(new_n1142), .Z(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT117), .B1(new_n933), .B2(G330), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1136), .A2(G330), .A3(new_n1137), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT117), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1148), .A2(new_n1149), .A3(new_n1143), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n914), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n1154), .A3(new_n915), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1109), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1151), .B(new_n1155), .C1(new_n1085), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n662), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1102), .A2(new_n1100), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1160), .A2(KEYINPUT57), .A3(new_n1155), .A4(new_n1151), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT118), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1147), .A2(new_n914), .A3(new_n1150), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n915), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1166), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n1160), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1159), .A2(new_n1163), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1151), .A2(new_n719), .A3(new_n1155), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n803), .B1(new_n201), .B2(new_n808), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1115), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n741), .A2(G132), .B1(new_n736), .B2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n743), .A2(G125), .B1(G150), .B2(new_n748), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n763), .C2(new_n1119), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n768), .B2(G137), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT59), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n750), .A2(G159), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n754), .C2(G124), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n742), .A2(new_n453), .B1(new_n202), .B2(new_n751), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G41), .B(new_n276), .C1(new_n754), .C2(G283), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n230), .B2(new_n737), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(G107), .C2(new_n780), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n743), .A2(G116), .B1(G68), .B2(new_n748), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT115), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(new_n324), .C2(new_n769), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT58), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n201), .B1(new_n271), .B2(G41), .ZN(new_n1192));
  AND4_X1   g0992(.A1(new_n1181), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1170), .B1(new_n1058), .B2(new_n1193), .C1(new_n1143), .C2(new_n830), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1169), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1168), .A2(new_n1195), .ZN(G375));
  NAND3_X1  g0996(.A1(new_n1089), .A2(new_n1085), .A3(new_n1092), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1107), .A2(new_n1110), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(new_n974), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT119), .Z(new_n1200));
  NAND2_X1  g1000(.A1(new_n1095), .A2(new_n719), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n924), .A2(new_n925), .A3(new_n830), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n768), .A2(G150), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n276), .B1(new_n1119), .B2(new_n753), .C1(new_n751), .C2(new_n202), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n741), .A2(new_n1171), .B1(G159), .B2(new_n736), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n201), .B2(new_n747), .C1(new_n822), .C2(new_n744), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G137), .C2(new_n780), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n348), .B1(new_n753), .B2(new_n774), .C1(new_n324), .C2(new_n747), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n736), .A2(G97), .B1(new_n750), .B2(G77), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n744), .B2(new_n782), .C1(new_n449), .C2(new_n742), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G283), .C2(new_n780), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n768), .A2(G107), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1203), .A2(new_n1207), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n720), .B1(G68), .B2(new_n809), .C1(new_n1213), .C2(new_n1058), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1201), .B1(new_n1202), .B2(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1200), .A2(new_n1215), .ZN(G381));
  INV_X1    g1016(.A(G390), .ZN(new_n1217));
  INV_X1    g1017(.A(G384), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OR4_X1    g1019(.A1(G396), .A2(G387), .A3(new_n1219), .A4(G393), .ZN(new_n1220));
  INV_X1    g1020(.A(G378), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1168), .A2(new_n1221), .A3(new_n1195), .ZN(new_n1222));
  OR3_X1    g1022(.A1(new_n1220), .A2(G381), .A3(new_n1222), .ZN(G407));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(G343), .C2(new_n1222), .ZN(G409));
  NAND2_X1  g1024(.A1(G387), .A2(new_n1217), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n999), .A2(G390), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(G393), .B(new_n792), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT125), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1225), .A2(new_n1226), .A3(KEYINPUT125), .A4(new_n1228), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(G387), .A2(new_n1217), .A3(KEYINPUT124), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT124), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n999), .B2(G390), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1235), .A3(new_n1226), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1231), .A2(new_n1232), .B1(new_n1227), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT61), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G375), .A2(G378), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n642), .A2(G213), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1157), .A2(new_n974), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1169), .A2(new_n1112), .A3(new_n1134), .A4(new_n1194), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1240), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(G2897), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1197), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n661), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1198), .B2(KEYINPUT60), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1251), .A2(new_n1218), .A3(new_n1215), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT120), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1218), .B1(new_n1251), .B2(new_n1215), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT120), .B(new_n1218), .C1(new_n1251), .C2(new_n1215), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1247), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT122), .ZN(new_n1258));
  INV_X1    g1058(.A(G2897), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1240), .B1(KEYINPUT121), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(KEYINPUT121), .B2(new_n1259), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1255), .A2(new_n1258), .A3(new_n1256), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1254), .A2(new_n1253), .ZN(new_n1263));
  OR3_X1    g1063(.A1(new_n1251), .A2(new_n1218), .A3(new_n1215), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1256), .A4(new_n1261), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT122), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1257), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1245), .B1(new_n1267), .B2(KEYINPUT123), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1262), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1257), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1269), .A2(KEYINPUT123), .A3(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1238), .B1(new_n1268), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1221), .B1(new_n1168), .B2(new_n1195), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1243), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1273), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1275), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1239), .A2(new_n1279), .A3(new_n1244), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1237), .B1(new_n1272), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT123), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1267), .A2(KEYINPUT123), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1245), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  NOR4_X1   g1089(.A1(new_n1274), .A2(new_n1275), .A3(new_n1289), .A4(new_n1243), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1237), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1280), .A2(new_n1289), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1288), .A2(new_n1291), .A3(new_n1238), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1283), .A2(new_n1293), .ZN(G405));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1222), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1295), .B1(new_n1296), .B2(new_n1274), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1239), .A2(KEYINPUT127), .A3(new_n1222), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1279), .A3(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1239), .A2(KEYINPUT127), .A3(new_n1222), .A4(new_n1275), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1236), .A2(new_n1227), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1299), .A2(new_n1300), .A3(new_n1237), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(G402));
endmodule


