//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT65), .B(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G58), .A2(G232), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G68), .Z(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G169), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G232), .A3(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(G226), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G97), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n248), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n257), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(G238), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT13), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT13), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n255), .A2(new_n264), .A3(new_n261), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n246), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT14), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(new_n265), .ZN(new_n268));
  INV_X1    g0068(.A(G179), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n265), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n264), .B1(new_n255), .B2(new_n261), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n267), .B(G169), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT75), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n266), .A2(KEYINPUT75), .A3(new_n267), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT74), .B(KEYINPUT12), .Z(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n279), .A2(new_n207), .A3(G1), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G68), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT65), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n278), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  OR3_X1    g0087(.A1(new_n281), .A2(KEYINPUT12), .A3(G68), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n206), .A2(G20), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT70), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n282), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n216), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n280), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n287), .A2(new_n288), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT11), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G50), .ZN(new_n298));
  XOR2_X1   g0098(.A(new_n298), .B(KEYINPUT73), .Z(new_n299));
  INV_X1    g0099(.A(G77), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n207), .A2(G33), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n286), .A2(new_n207), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n293), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n295), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n303), .A2(new_n296), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n277), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n268), .A2(G200), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n263), .A2(G190), .A3(new_n265), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n247), .A2(G222), .A3(new_n249), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n247), .A2(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G223), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n313), .B1(new_n300), .B2(new_n247), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n254), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT67), .B(G226), .Z(new_n318));
  AOI21_X1  g0118(.A(new_n258), .B1(new_n260), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n246), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n294), .B(KEYINPUT69), .ZN(new_n322));
  OR3_X1    g0122(.A1(new_n290), .A2(KEYINPUT71), .A3(new_n202), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT71), .B1(new_n290), .B2(new_n202), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n297), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT8), .B(G58), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT68), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G58), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n326), .B1(new_n332), .B2(new_n301), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(new_n293), .B1(new_n202), .B2(new_n280), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n325), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n317), .A2(new_n269), .A3(new_n319), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n321), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n335), .B(KEYINPUT9), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n320), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(G200), .B2(new_n320), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT10), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(KEYINPUT10), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n290), .A2(new_n300), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n294), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G77), .B2(new_n281), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT15), .B(G87), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n301), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n207), .A2(new_n251), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n327), .A2(new_n352), .B1(new_n207), .B2(new_n300), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(KEYINPUT72), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(KEYINPUT72), .B2(new_n353), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n349), .B1(new_n293), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n247), .A2(G232), .A3(new_n249), .ZN(new_n357));
  INV_X1    g0157(.A(G107), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n357), .B1(new_n358), .B2(new_n247), .C1(new_n314), .C2(new_n220), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n254), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n258), .B1(G244), .B2(new_n260), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n356), .B1(new_n340), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n362), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n356), .B1(new_n246), .B2(new_n362), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n269), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n312), .A2(new_n346), .A3(new_n367), .A4(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n247), .A2(G226), .A3(G1698), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G33), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n373), .A2(new_n375), .A3(G223), .A4(new_n249), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n254), .ZN(new_n379));
  INV_X1    g0179(.A(new_n216), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G41), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n256), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n260), .A2(G232), .B1(new_n382), .B2(new_n259), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n379), .A2(G190), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n365), .B1(new_n379), .B2(new_n383), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n332), .A2(new_n290), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n322), .A2(new_n387), .B1(new_n280), .B2(new_n332), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n373), .A2(new_n375), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n390), .B2(new_n207), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n247), .B2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT76), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n286), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n213), .B1(new_n219), .B2(new_n330), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(G20), .B1(G159), .B2(new_n297), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT16), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n392), .B(G20), .C1(new_n373), .C2(new_n375), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n391), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(new_n399), .A3(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n293), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n386), .B(new_n388), .C1(new_n400), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n389), .B1(new_n391), .B2(new_n401), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT76), .B1(new_n394), .B2(KEYINPUT7), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n219), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n201), .B1(new_n286), .B2(G58), .ZN(new_n412));
  INV_X1    g0212(.A(G159), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n412), .A2(new_n207), .B1(new_n413), .B2(new_n352), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n408), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n403), .A2(new_n293), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n417), .A2(KEYINPUT17), .A3(new_n388), .A4(new_n386), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n407), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT78), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n379), .A2(new_n383), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n269), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n246), .B1(new_n379), .B2(new_n383), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT77), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(G169), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT77), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n426), .B(new_n427), .C1(new_n269), .C2(new_n422), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n417), .A2(new_n388), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(KEYINPUT18), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n425), .A2(new_n428), .ZN(new_n433));
  INV_X1    g0233(.A(new_n388), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n415), .B2(new_n416), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n432), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n407), .A2(KEYINPUT78), .A3(new_n418), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n421), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n371), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G45), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(G1), .ZN(new_n442));
  INV_X1    g0242(.A(G41), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n442), .B(KEYINPUT83), .C1(KEYINPUT5), .C2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n206), .B(G45), .C1(new_n443), .C2(KEYINPUT5), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT83), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(KEYINPUT5), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n444), .A2(new_n447), .A3(new_n382), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n254), .ZN(new_n450));
  INV_X1    g0250(.A(new_n448), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n445), .ZN(new_n452));
  INV_X1    g0252(.A(G257), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n247), .A2(G244), .A3(new_n249), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT82), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT4), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT4), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(KEYINPUT82), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n390), .A2(new_n249), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n460), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n454), .B1(new_n462), .B2(new_n254), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n246), .ZN(new_n464));
  AOI211_X1 g0264(.A(new_n269), .B(new_n454), .C1(new_n462), .C2(new_n254), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT84), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n358), .B1(new_n409), .B2(new_n410), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT6), .ZN(new_n471));
  AND2_X1   g0271(.A1(G97), .A2(G107), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n358), .A2(KEYINPUT6), .A3(G97), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n207), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n297), .A2(KEYINPUT79), .A3(G77), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT79), .B1(new_n297), .B2(G77), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n470), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT79), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n352), .B2(new_n300), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n297), .A2(KEYINPUT79), .A3(G77), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g0284(.A(G97), .B(G107), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n471), .A2(new_n252), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n485), .A2(new_n471), .B1(new_n358), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(KEYINPUT80), .B(new_n484), .C1(new_n487), .C2(new_n207), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n293), .B1(new_n469), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT81), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT81), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(new_n293), .C1(new_n469), .C2(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n281), .A2(G97), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n251), .A2(G1), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n280), .A2(new_n293), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(new_n497), .B2(G97), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n468), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n498), .ZN(new_n500));
  AOI211_X1 g0300(.A(KEYINPUT84), .B(new_n500), .C1(new_n491), .C2(new_n493), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n467), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n491), .B2(new_n493), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n463), .A2(G190), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n503), .B(new_n504), .C1(new_n365), .C2(new_n463), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n390), .A2(G303), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n373), .A2(new_n375), .A3(G264), .A4(G1698), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n373), .A2(new_n375), .A3(G257), .A4(new_n249), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT90), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n450), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n507), .A2(KEYINPUT90), .A3(new_n508), .A4(new_n509), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n497), .A2(G116), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n281), .A2(G116), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G116), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G20), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n293), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n207), .C1(G33), .C2(new_n252), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT20), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n293), .A3(new_n519), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n515), .B(new_n517), .C1(new_n523), .C2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n450), .B(G270), .C1(new_n451), .C2(new_n445), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n449), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n514), .A2(G179), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT91), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n514), .A2(new_n530), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n524), .B(new_n525), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n516), .B1(new_n497), .B2(G116), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n246), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(KEYINPUT21), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT21), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n527), .A2(G169), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n529), .B1(new_n512), .B2(new_n513), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n541), .A2(KEYINPUT91), .A3(G179), .A4(new_n527), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n533), .A2(new_n538), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n527), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n541), .B2(new_n365), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(G190), .B2(new_n541), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT87), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n549), .A2(new_n550), .A3(new_n207), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n549), .B2(new_n207), .ZN(new_n552));
  NOR3_X1   g0352(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n373), .A2(new_n375), .A3(new_n207), .A4(G68), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n301), .A2(new_n252), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(KEYINPUT19), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n293), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n350), .A2(new_n280), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n497), .A2(G87), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n442), .A2(G250), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n442), .A2(new_n256), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n450), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n251), .A2(new_n518), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G238), .A2(G1698), .ZN(new_n566));
  INV_X1    g0366(.A(G244), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(G1698), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n568), .B2(new_n247), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT85), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n254), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n220), .A2(new_n249), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n390), .A2(new_n574), .B1(new_n251), .B2(new_n518), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(KEYINPUT85), .ZN(new_n576));
  OAI211_X1 g0376(.A(G190), .B(new_n564), .C1(new_n571), .C2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n561), .B1(new_n577), .B2(KEYINPUT89), .ZN(new_n578));
  INV_X1    g0378(.A(new_n564), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n450), .B1(new_n575), .B2(KEYINPUT85), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n569), .A2(new_n570), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT89), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(G190), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n578), .B(new_n584), .C1(new_n365), .C2(new_n582), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n269), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n582), .A2(KEYINPUT86), .A3(new_n269), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n564), .B1(new_n571), .B2(new_n576), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n246), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n294), .B1(G1), .B2(new_n251), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n350), .B(KEYINPUT88), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n558), .B(new_n559), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n588), .A2(new_n589), .A3(new_n591), .A4(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n585), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n373), .A2(new_n375), .A3(G257), .A4(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n373), .A2(new_n375), .A3(G250), .A4(new_n249), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G294), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n254), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n450), .B(G264), .C1(new_n451), .C2(new_n445), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT93), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT93), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(G179), .A3(new_n449), .A4(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n601), .A2(new_n449), .A3(new_n602), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G169), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n373), .A2(new_n375), .A3(new_n207), .A4(G87), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT92), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT22), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT23), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n207), .B2(G107), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n358), .A2(KEYINPUT23), .A3(G20), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n565), .A2(new_n207), .ZN(new_n619));
  XNOR2_X1  g0419(.A(KEYINPUT92), .B(KEYINPUT22), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n619), .C1(new_n610), .C2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT24), .B1(new_n614), .B2(new_n621), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n610), .A2(new_n620), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT24), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n618), .A2(new_n619), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .A4(new_n613), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n293), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT25), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n281), .B2(G107), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n280), .A2(KEYINPUT25), .A3(new_n358), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n630), .A2(new_n631), .B1(new_n497), .B2(G107), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n607), .A2(new_n609), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n604), .A2(new_n449), .A3(new_n606), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n365), .ZN(new_n635));
  INV_X1    g0435(.A(new_n608), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n340), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n628), .A2(new_n632), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n633), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n548), .A2(new_n596), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n440), .A2(new_n506), .A3(new_n642), .ZN(G372));
  NOR2_X1   g0443(.A1(new_n423), .A2(new_n424), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT18), .B1(new_n435), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n435), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n432), .ZN(new_n647));
  INV_X1    g0447(.A(new_n370), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n307), .B1(new_n310), .B2(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n407), .A2(KEYINPUT78), .A3(new_n418), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT78), .B1(new_n407), .B2(new_n418), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n645), .B(new_n647), .C1(new_n649), .C2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n344), .A2(new_n345), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n338), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n533), .A2(new_n538), .A3(new_n543), .ZN(new_n657));
  INV_X1    g0457(.A(new_n542), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n657), .A2(new_n633), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT94), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n582), .B2(new_n365), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n590), .A2(KEYINPUT94), .A3(G200), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n578), .A2(new_n661), .A3(new_n662), .A4(new_n584), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n586), .A2(new_n591), .A3(new_n594), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n634), .A2(new_n365), .B1(new_n340), .B2(new_n636), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n663), .B(new_n664), .C1(new_n665), .C2(new_n639), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n502), .A3(new_n505), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n596), .B(new_n467), .C1(new_n499), .C2(new_n501), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n503), .A2(new_n466), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n663), .A2(new_n664), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n668), .A2(new_n670), .A3(new_n675), .A4(new_n664), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n440), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n656), .A2(new_n677), .ZN(G369));
  NAND3_X1  g0478(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G213), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(G343), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n639), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n641), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT95), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n633), .A2(new_n684), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n684), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n548), .B1(new_n545), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n544), .A2(new_n527), .A3(new_n684), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT96), .Z(new_n699));
  OAI211_X1 g0499(.A(new_n544), .B(new_n692), .C1(new_n689), .C2(new_n690), .ZN(new_n700));
  INV_X1    g0500(.A(new_n633), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n684), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n210), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n553), .A2(new_n518), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(G1), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n215), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n707), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n668), .A2(new_n664), .ZN(new_n714));
  NOR4_X1   g0514(.A1(new_n672), .A2(new_n503), .A3(new_n466), .A4(new_n674), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n669), .B2(new_n674), .ZN(new_n716));
  OAI211_X1 g0516(.A(KEYINPUT29), .B(new_n692), .C1(new_n714), .C2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n676), .A2(new_n692), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(KEYINPUT29), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n642), .A2(new_n502), .A3(new_n505), .A4(new_n692), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n463), .A2(new_n604), .A3(new_n606), .A4(new_n582), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n541), .A2(G179), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n723), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n604), .A2(new_n582), .A3(new_n606), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT30), .A4(new_n463), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n541), .A2(new_n582), .A3(G179), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n462), .A2(new_n254), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n728), .B(new_n634), .C1(new_n729), .C2(new_n454), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n724), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT31), .B1(new_n731), .B2(new_n684), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n720), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G330), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n719), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n713), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n279), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n206), .B1(new_n740), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n706), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT101), .Z(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n695), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n216), .B1(G20), .B2(new_n246), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n215), .A2(new_n441), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n705), .A2(new_n247), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(new_n244), .C2(new_n441), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n705), .A2(new_n390), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n757), .A2(G355), .B1(new_n518), .B2(new_n705), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n753), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n340), .A2(G179), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n207), .ZN(new_n761));
  INV_X1    g0561(.A(G294), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n207), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(G303), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n761), .A2(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(new_n340), .A3(new_n365), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n247), .B1(new_n768), .B2(G329), .ZN(new_n769));
  INV_X1    g0569(.A(G283), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n763), .A2(new_n340), .A3(G200), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(G20), .A2(G179), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT97), .Z(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n340), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n766), .B(new_n772), .C1(G326), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n775), .A2(G190), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT33), .B(G317), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT98), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n774), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(G200), .B1(new_n774), .B2(new_n783), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n784), .A2(new_n340), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G322), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n784), .A2(G190), .A3(new_n785), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n781), .B1(new_n782), .B2(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n330), .A2(new_n788), .B1(new_n786), .B2(new_n300), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT99), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n767), .A2(new_n413), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  INV_X1    g0593(.A(new_n778), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(new_n252), .B2(new_n761), .C1(new_n282), .C2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n795), .B1(G50), .B2(new_n776), .ZN(new_n796));
  INV_X1    g0596(.A(G87), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n247), .B1(new_n771), .B2(new_n358), .C1(new_n797), .C2(new_n764), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT100), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n791), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n789), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n759), .B1(new_n801), .B2(new_n751), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n744), .B1(new_n750), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n695), .B(new_n696), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n744), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT102), .ZN(G396));
  NAND2_X1  g0606(.A1(new_n648), .A2(new_n692), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n363), .A2(new_n366), .B1(new_n356), .B2(new_n692), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n370), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n718), .B(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(new_n736), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n743), .B1(new_n812), .B2(new_n736), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n751), .A2(new_n745), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n744), .B1(new_n300), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n788), .A2(new_n762), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n797), .A2(new_n771), .B1(new_n764), .B2(new_n358), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n390), .B1(new_n767), .B2(new_n782), .C1(new_n761), .C2(new_n252), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(new_n778), .C2(G283), .ZN(new_n821));
  INV_X1    g0621(.A(new_n776), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n765), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n786), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n818), .B(new_n823), .C1(G116), .C2(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G137), .A2(new_n776), .B1(new_n778), .B2(G150), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n827), .B2(new_n788), .C1(new_n413), .C2(new_n786), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT34), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n247), .B1(new_n767), .B2(new_n831), .C1(new_n202), .C2(new_n764), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n761), .A2(new_n330), .B1(new_n771), .B2(new_n282), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n828), .C2(new_n829), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n825), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n751), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n817), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT103), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n746), .B2(new_n811), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n838), .B2(new_n837), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT104), .Z(new_n842));
  NOR2_X1   g0642(.A1(new_n815), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G384));
  INV_X1    g0644(.A(new_n487), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n845), .A2(KEYINPUT35), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(KEYINPUT35), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n846), .A2(new_n847), .A3(G116), .A4(new_n217), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT36), .ZN(new_n849));
  OAI21_X1  g0649(.A(G77), .B1(new_n219), .B2(new_n330), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n711), .A2(new_n850), .B1(G50), .B2(new_n282), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(G1), .A3(new_n279), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT105), .Z(new_n853));
  NAND2_X1  g0653(.A1(new_n277), .A2(new_n310), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n684), .B1(new_n304), .B2(new_n305), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n855), .B(KEYINPUT106), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n310), .B(new_n858), .C1(new_n277), .C2(new_n306), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n676), .A2(new_n692), .A3(new_n811), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n807), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n435), .A2(new_n682), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n429), .A2(new_n430), .ZN(new_n867));
  XNOR2_X1  g0667(.A(KEYINPUT109), .B(KEYINPUT37), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n866), .A2(new_n867), .A3(new_n405), .A4(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n282), .B1(new_n394), .B2(new_n395), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n408), .B1(new_n414), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n403), .A3(new_n293), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n388), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT107), .ZN(new_n875));
  INV_X1    g0675(.A(new_n644), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT107), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n873), .A2(new_n877), .A3(new_n388), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n405), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT108), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT108), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n879), .A2(new_n882), .A3(new_n405), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n875), .A2(new_n878), .ZN(new_n884));
  INV_X1    g0684(.A(new_n682), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n870), .B1(new_n887), .B2(KEYINPUT37), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n652), .B2(new_n437), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n864), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n886), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n439), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n880), .A2(KEYINPUT108), .B1(new_n885), .B2(new_n884), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(new_n883), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n892), .B(KEYINPUT38), .C1(new_n895), .C2(new_n870), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n863), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n647), .A2(new_n645), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n682), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n307), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n684), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n890), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n904));
  INV_X1    g0704(.A(new_n868), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n405), .B1(new_n435), .B2(new_n682), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n646), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT110), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT110), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n909), .B(new_n905), .C1(new_n906), .C2(new_n646), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n908), .A2(new_n869), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT111), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n407), .A2(new_n912), .A3(new_n418), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n647), .A3(new_n645), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n407), .B2(new_n418), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n865), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n864), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n896), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n903), .B(new_n904), .C1(new_n920), .C2(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n901), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n440), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n656), .B1(new_n719), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n810), .B1(new_n857), .B2(new_n859), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n735), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n897), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n735), .A2(new_n926), .A3(KEYINPUT40), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n919), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n440), .A2(new_n735), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(G330), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n925), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n206), .B2(new_n740), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n925), .A2(new_n938), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n849), .B(new_n853), .C1(new_n940), .C2(new_n941), .ZN(G367));
  OR2_X1    g0742(.A1(new_n503), .A2(new_n692), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n506), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT113), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT113), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n506), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n671), .A2(new_n684), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT42), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n544), .A2(new_n692), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n950), .A2(new_n951), .A3(new_n691), .A4(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n945), .A2(new_n947), .B1(new_n671), .B2(new_n684), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT42), .B1(new_n955), .B2(new_n700), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT43), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n561), .A2(new_n684), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n664), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT112), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n673), .B2(new_n960), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n502), .B1(new_n955), .B2(new_n701), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n692), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n958), .A2(new_n959), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(new_n959), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n963), .A2(new_n959), .ZN(new_n968));
  INV_X1    g0768(.A(new_n965), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n967), .B(new_n968), .C1(new_n969), .C2(new_n957), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n699), .A2(new_n955), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n706), .B(KEYINPUT41), .Z(new_n975));
  INV_X1    g0775(.A(KEYINPUT44), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n950), .B2(new_n703), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n955), .A2(new_n702), .A3(KEYINPUT44), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n950), .A2(KEYINPUT45), .A3(new_n703), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n955), .B2(new_n702), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n699), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n691), .A2(new_n953), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n700), .A2(new_n697), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n697), .B1(new_n986), .B2(new_n700), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n738), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n979), .A2(new_n699), .A3(new_n983), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n985), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n975), .B1(new_n993), .B2(new_n738), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n973), .B(new_n974), .C1(new_n994), .C2(new_n742), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n237), .A2(new_n705), .A3(new_n247), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n752), .B1(new_n210), .B2(new_n350), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n743), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(G137), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n247), .B1(new_n767), .B2(new_n999), .C1(new_n300), .C2(new_n771), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n761), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(G68), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n330), .B2(new_n764), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1000), .B(new_n1003), .C1(G159), .C2(new_n778), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n202), .B2(new_n786), .C1(new_n827), .C2(new_n822), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n788), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1005), .B1(G150), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT46), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n764), .A2(new_n1008), .A3(new_n518), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT114), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n794), .B2(new_n762), .C1(new_n782), .C2(new_n822), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n771), .A2(new_n252), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n247), .B(new_n1012), .C1(G317), .C2(new_n768), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1008), .B1(new_n764), .B2(new_n518), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n358), .C2(new_n761), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n770), .A2(new_n786), .B1(new_n788), .B2(new_n765), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1011), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1007), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT47), .Z(new_n1019));
  AOI21_X1  g0819(.A(new_n998), .B1(new_n1019), .B2(new_n751), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n963), .A2(new_n749), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n995), .A2(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n1006), .A2(G317), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G311), .A2(new_n778), .B1(new_n776), .B2(G322), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n765), .C2(new_n786), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n764), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1001), .A2(G283), .B1(new_n1030), .B2(G294), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT49), .Z(new_n1033));
  AOI21_X1  g0833(.A(new_n247), .B1(new_n768), .B2(G326), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n518), .B2(new_n771), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n788), .A2(new_n202), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n593), .A2(new_n761), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n764), .A2(new_n300), .ZN(new_n1039));
  INV_X1    g0839(.A(G150), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n247), .B1(new_n767), .B2(new_n1040), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1038), .A2(new_n1012), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n413), .B2(new_n822), .C1(new_n332), .C2(new_n794), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1037), .B(new_n1043), .C1(G68), .C2(new_n824), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n751), .B1(new_n1036), .B2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n757), .A2(new_n708), .B1(new_n358), .B2(new_n705), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n327), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n202), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n709), .B(new_n441), .C1(new_n282), .C2(new_n300), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n755), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT115), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n233), .B2(new_n441), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1046), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n744), .B1(new_n1056), .B2(new_n752), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1045), .B(new_n1057), .C1(new_n691), .C2(new_n748), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT116), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n742), .B2(new_n989), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n990), .A2(new_n706), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n989), .A2(new_n738), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(G393));
  INV_X1    g0863(.A(new_n992), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT117), .ZN(new_n1065));
  OAI21_X1  g0865(.A(KEYINPUT117), .B1(new_n1064), .B2(new_n984), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n742), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n247), .B1(new_n767), .B2(new_n827), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n761), .A2(new_n300), .B1(new_n764), .B2(new_n219), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n771), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1068), .B(new_n1069), .C1(G87), .C2(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n202), .B2(new_n794), .C1(new_n327), .C2(new_n786), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1006), .A2(G159), .B1(G150), .B2(new_n776), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1006), .A2(G311), .B1(G317), .B2(new_n776), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT52), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n390), .B1(new_n767), .B2(new_n787), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n761), .A2(new_n518), .B1(new_n764), .B2(new_n770), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G107), .C2(new_n1070), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n765), .B2(new_n794), .C1(new_n762), .C2(new_n786), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1072), .A2(new_n1074), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n751), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n755), .A2(new_n241), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n753), .B1(G97), .B2(new_n705), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n744), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n747), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1082), .B(new_n1085), .C1(new_n950), .C2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n991), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n993), .A2(new_n706), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1067), .B(new_n1087), .C1(new_n1088), .C2(new_n1089), .ZN(G390));
  INV_X1    g0890(.A(new_n904), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT39), .B1(new_n918), .B2(new_n896), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1091), .A2(new_n1092), .B1(new_n863), .B2(new_n903), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n692), .B(new_n809), .C1(new_n714), .C2(new_n716), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT118), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n807), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n1094), .B2(new_n807), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n861), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n919), .B1(new_n902), .B2(new_n684), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1093), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n696), .B1(new_n720), .B2(new_n734), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n811), .A3(new_n860), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1093), .B(new_n1102), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n440), .A2(new_n1101), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n656), .B(new_n1107), .C1(new_n719), .C2(new_n923), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1094), .A2(new_n807), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT118), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1094), .A2(new_n1095), .A3(new_n807), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n860), .B1(new_n1101), .B2(new_n811), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1103), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n862), .A2(new_n807), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1103), .B2(new_n1113), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1108), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1106), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1104), .A2(new_n1105), .A3(new_n1118), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n706), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1104), .A2(new_n742), .A3(new_n1105), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT120), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n745), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n390), .B1(new_n768), .B2(G125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n202), .B2(new_n771), .C1(new_n413), .C2(new_n761), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT53), .B1(new_n1030), .B2(G150), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1030), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n794), .A2(new_n999), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1127), .B(new_n1130), .C1(G128), .C2(new_n776), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1131), .B1(new_n831), .B2(new_n788), .C1(new_n786), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT119), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n390), .B1(new_n767), .B2(new_n762), .C1(new_n797), .C2(new_n764), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n761), .A2(new_n300), .B1(new_n771), .B2(new_n282), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n794), .B2(new_n358), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G283), .B2(new_n776), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n252), .B2(new_n786), .C1(new_n518), .C2(new_n788), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n751), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n744), .B1(new_n332), .B2(new_n816), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1125), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1123), .A2(new_n1124), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1124), .B1(new_n1123), .B2(new_n1146), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1122), .B1(new_n1147), .B2(new_n1148), .ZN(G378));
  INV_X1    g0949(.A(new_n1108), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1121), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n927), .B1(new_n896), .B2(new_n890), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n933), .B(G330), .C1(new_n1153), .C2(KEYINPUT40), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n335), .A2(new_n885), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n346), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n346), .A2(new_n1155), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OR3_X1    g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1154), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n931), .A2(G330), .A3(new_n933), .A4(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n922), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n921), .A4(new_n901), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1152), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1151), .A2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1121), .A2(new_n1150), .B1(new_n1168), .B2(new_n1167), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n706), .C1(KEYINPUT57), .C2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n741), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1002), .B1(new_n330), .B2(new_n771), .C1(new_n770), .C2(new_n767), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n390), .A2(new_n443), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1039), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT121), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n776), .A2(G116), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1177), .B2(new_n1176), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1174), .B(new_n1179), .C1(G97), .C2(new_n778), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n358), .B2(new_n788), .C1(new_n593), .C2(new_n786), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT58), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1175), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1132), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1030), .A2(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n1040), .B2(new_n761), .C1(new_n794), .C2(new_n831), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G125), .B2(new_n776), .ZN(new_n1190));
  INV_X1    g0990(.A(G128), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1190), .B1(new_n1191), .B2(new_n788), .C1(new_n999), .C2(new_n786), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1070), .A2(G159), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n768), .C2(G124), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n751), .B1(new_n1186), .B2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT122), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n744), .B1(new_n202), .B2(new_n816), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT123), .Z(new_n1202));
  OAI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(new_n746), .C2(new_n1162), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT124), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1173), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1172), .A2(new_n1205), .ZN(G375));
  OAI21_X1  g1006(.A(new_n861), .B1(new_n736), .B2(new_n810), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1207), .A2(new_n1102), .B1(new_n807), .B2(new_n862), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1108), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n975), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1119), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1209), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n861), .A2(new_n745), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n771), .A2(new_n300), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n390), .B1(new_n767), .B2(new_n765), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G97), .C2(new_n1030), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n593), .B2(new_n761), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n518), .A2(new_n794), .B1(new_n822), .B2(new_n762), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n824), .B2(G107), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT125), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1218), .B(new_n1221), .C1(G283), .C2(new_n1006), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n788), .A2(new_n999), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n761), .A2(new_n202), .B1(new_n764), .B2(new_n413), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n247), .B1(new_n767), .B2(new_n1191), .C1(new_n330), .C2(new_n771), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n776), .C2(G132), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n794), .B2(new_n1132), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1223), .B(new_n1227), .C1(G150), .C2(new_n824), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n751), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n744), .B1(new_n282), .B2(new_n816), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1213), .A2(new_n742), .B1(new_n1214), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1212), .A2(new_n1232), .ZN(G381));
  NOR4_X1   g1033(.A1(G381), .A2(G393), .A3(G384), .A4(G396), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1089), .B1(new_n1235), .B2(new_n990), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1067), .A2(new_n1087), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1123), .A2(new_n1146), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n707), .B1(new_n1106), .B2(new_n1119), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1241), .B2(new_n1121), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OR4_X1    g1043(.A1(G387), .A2(new_n1239), .A3(G375), .A4(new_n1243), .ZN(G407));
  NAND2_X1  g1044(.A1(new_n683), .A2(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G407), .B(G213), .C1(G375), .C2(new_n1247), .ZN(G409));
  INV_X1    g1048(.A(KEYINPUT63), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1172), .A2(G378), .A3(new_n1205), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1171), .A2(new_n1211), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1205), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1242), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1245), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n1108), .A4(new_n1117), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT127), .ZN(new_n1257));
  XOR2_X1   g1057(.A(KEYINPUT126), .B(KEYINPUT60), .Z(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1210), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1118), .A2(new_n707), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G384), .B1(new_n1262), .B2(new_n1232), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT127), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1256), .B(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1232), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(new_n843), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1263), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1249), .B1(new_n1255), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1246), .A2(G2897), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1263), .B2(new_n1268), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1262), .A2(G384), .A3(new_n1232), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1267), .A2(new_n843), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1276), .A3(new_n1272), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT61), .B1(new_n1255), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(new_n1238), .ZN(new_n1280));
  XOR2_X1   g1080(.A(G393), .B(G396), .Z(new_n1281));
  NAND3_X1  g1081(.A1(G390), .A2(new_n995), .A3(new_n1022), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1281), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1246), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(KEYINPUT63), .A3(new_n1269), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1271), .A2(new_n1279), .A3(new_n1285), .A4(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1286), .A2(new_n1289), .A3(new_n1269), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT61), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1286), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1289), .B1(new_n1286), .B2(new_n1269), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1290), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1288), .B1(new_n1295), .B2(new_n1285), .ZN(G405));
  OR2_X1    g1096(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1172), .A2(G378), .A3(new_n1205), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1243), .B1(new_n1172), .B2(new_n1205), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1270), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1269), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1297), .B(new_n1303), .ZN(G402));
endmodule


