//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n607, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n452), .B(new_n453), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  NAND2_X1  g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT68), .Z(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n468), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(G137), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G137), .A4(new_n466), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n475), .A2(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n472), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n472), .A2(new_n466), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NOR2_X1   g065(.A1(new_n466), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n485), .B2(G126), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n470), .B2(new_n471), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n496), .B(new_n499), .C1(new_n471), .C2(new_n470), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT70), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .A3(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n509), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n511), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(new_n506), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n518), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  AOI22_X1  g097(.A1(new_n507), .A2(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n516), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n510), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n524), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n506), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(G90), .A2(new_n523), .B1(new_n510), .B2(G52), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n534), .A2(new_n535), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n506), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n510), .A2(G43), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n523), .A2(G81), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n517), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n523), .A2(KEYINPUT73), .A3(G91), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n516), .A2(G65), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n554), .A2(new_n555), .B1(G651), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n513), .A2(G53), .A3(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n510), .A2(new_n563), .A3(G53), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n562), .B1(new_n561), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  XNOR2_X1  g143(.A(new_n531), .B(KEYINPUT74), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G286));
  NAND2_X1  g145(.A1(new_n523), .A2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n510), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(G86), .A2(new_n523), .B1(new_n510), .B2(G48), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  INV_X1    g151(.A(new_n515), .ZN(new_n577));
  NOR2_X1   g152(.A1(KEYINPUT5), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G61), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n576), .B1(new_n581), .B2(G651), .ZN(new_n582));
  AOI211_X1 g157(.A(KEYINPUT75), .B(new_n506), .C1(new_n579), .C2(new_n580), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n575), .B1(new_n582), .B2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(G85), .A2(new_n523), .B1(new_n510), .B2(G47), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT76), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n506), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(new_n523), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  AOI22_X1  g166(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n506), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n593), .B2(new_n592), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n510), .A2(G54), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(G171), .ZN(G284));
  XOR2_X1   g175(.A(G284), .B(KEYINPUT78), .Z(G321));
  INV_X1    g176(.A(G299), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n598), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n598), .B2(G286), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G297));
  XNOR2_X1  g180(.A(new_n604), .B(KEYINPUT79), .ZN(G280));
  AND3_X1   g181(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n485), .A2(G123), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT81), .Z(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(KEYINPUT82), .ZN(new_n617));
  INV_X1    g192(.A(G111), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n616), .A2(KEYINPUT82), .B1(new_n618), .B2(G2105), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n483), .A2(G135), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT83), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n478), .A2(new_n467), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  NOR2_X1   g202(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n623), .B(new_n629), .C1(new_n627), .C2(new_n624), .ZN(G156));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT85), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n665), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT20), .Z(new_n669));
  AOI211_X1 g244(.A(new_n667), .B(new_n669), .C1(new_n662), .C2(new_n666), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  XOR2_X1   g246(.A(G1981), .B(G1986), .Z(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n671), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G229));
  MUX2_X1   g253(.A(G6), .B(G305), .S(G16), .Z(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT32), .B(G1981), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G166), .B2(new_n682), .ZN(new_n684));
  INV_X1    g259(.A(G1971), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(G23), .ZN(new_n687));
  INV_X1    g262(.A(G288), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n682), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT33), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  AND3_X1   g266(.A1(new_n681), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n682), .A2(G24), .ZN(new_n695));
  INV_X1    g270(.A(G290), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n682), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1986), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n483), .A2(G131), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n485), .A2(G119), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n466), .A2(G107), .ZN(new_n701));
  OAI21_X1  g276(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G25), .B(new_n703), .S(G29), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n698), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n694), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(KEYINPUT87), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n694), .A2(new_n711), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n692), .A2(new_n693), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT36), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n713), .A2(new_n718), .A3(new_n715), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G29), .A2(G35), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G162), .B2(G29), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G2090), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G1961), .ZN(new_n727));
  NOR2_X1   g302(.A1(G171), .A2(new_n682), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G5), .B2(new_n682), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT93), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n733), .B(new_n734), .Z(new_n735));
  AOI22_X1  g310(.A1(new_n485), .A2(G129), .B1(G105), .B2(new_n467), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n483), .A2(G141), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n731), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n731), .B2(G32), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  NAND2_X1  g318(.A1(G160), .A2(G29), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT24), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n731), .B1(new_n745), .B2(G34), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(KEYINPUT91), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(G34), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n746), .B2(KEYINPUT91), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n744), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n742), .B1(new_n743), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n731), .A2(G27), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n731), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2078), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n546), .A2(G16), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G16), .B2(G19), .ZN(new_n756));
  INV_X1    g331(.A(G1341), .ZN(new_n757));
  OAI22_X1  g332(.A1(new_n756), .A2(new_n757), .B1(new_n750), .B2(new_n743), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n754), .B(new_n758), .C1(new_n740), .C2(new_n741), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n682), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n682), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n756), .A2(new_n757), .B1(G1966), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n751), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n483), .A2(G140), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n485), .A2(G128), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n466), .A2(G116), .ZN(new_n766));
  OAI21_X1  g341(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G29), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n731), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT88), .Z(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G2067), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G33), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT89), .Z(new_n776));
  NAND3_X1  g351(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT25), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n478), .A2(G127), .ZN(new_n779));
  NAND2_X1  g354(.A1(G115), .A2(G2104), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n466), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n778), .B(new_n781), .C1(G139), .C2(new_n483), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n776), .B1(new_n783), .B2(new_n731), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT90), .B(G2072), .Z(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT31), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G11), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(G11), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(G28), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n731), .B1(new_n791), .B2(G28), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n789), .B(new_n790), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n621), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G29), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n786), .A2(new_n787), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n773), .A2(G2067), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n729), .B2(new_n727), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n763), .A2(new_n774), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n682), .A2(G4), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n607), .B2(new_n682), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(G1348), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n682), .A2(G20), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT96), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT23), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G299), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G1956), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n802), .A2(G1348), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n761), .A2(G1966), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT94), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n803), .A2(new_n809), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n720), .A2(new_n730), .A3(new_n800), .A4(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  NOR2_X1   g390(.A1(new_n597), .A2(new_n608), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n523), .A2(G93), .ZN(new_n819));
  INV_X1    g394(.A(new_n510), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT98), .B(G55), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n819), .B1(new_n820), .B2(new_n821), .C1(new_n506), .C2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n545), .B(new_n823), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n818), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n826));
  AOI21_X1  g401(.A(G860), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n823), .A2(G860), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT37), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(G145));
  XNOR2_X1  g406(.A(new_n703), .B(new_n626), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n485), .A2(G130), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT101), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n483), .A2(G142), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n466), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n832), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n498), .A2(new_n840), .A3(new_n500), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n498), .B2(new_n500), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n494), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n768), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n735), .A2(new_n738), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n782), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n782), .B(new_n847), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n839), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n851), .A3(new_n839), .ZN(new_n854));
  XNOR2_X1  g429(.A(G160), .B(G162), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n621), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n839), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n850), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n856), .B1(new_n850), .B2(new_n859), .ZN(new_n861));
  AOI21_X1  g436(.A(G37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g439(.A1(new_n607), .A2(G299), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n602), .A2(new_n597), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n824), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n610), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT105), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT41), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n866), .A2(KEYINPUT106), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n602), .A2(new_n597), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n875), .A2(new_n865), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n874), .B1(new_n878), .B2(KEYINPUT41), .ZN(new_n879));
  INV_X1    g454(.A(new_n871), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n869), .A2(new_n882), .A3(new_n871), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n873), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT42), .ZN(new_n885));
  XNOR2_X1  g460(.A(G290), .B(G288), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(G303), .B(G305), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n889), .B1(new_n886), .B2(new_n887), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n884), .A2(KEYINPUT42), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n885), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n885), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(G868), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n823), .A2(new_n598), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(G295));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n899), .ZN(G331));
  NAND2_X1  g476(.A1(G301), .A2(new_n531), .ZN(new_n902));
  NAND2_X1  g477(.A1(G171), .A2(new_n569), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n824), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n870), .A2(new_n903), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT108), .B1(new_n867), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n867), .A2(KEYINPUT108), .A3(new_n910), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n875), .A2(KEYINPUT41), .A3(new_n865), .A4(new_n877), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n908), .B(new_n909), .C1(new_n911), .C2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n911), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(new_n907), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n869), .A2(new_n907), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT109), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n915), .B(new_n893), .C1(new_n917), .C2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n905), .A2(new_n906), .B1(new_n865), .B2(new_n866), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n879), .B2(new_n908), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n894), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT110), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n920), .A2(new_n924), .A3(new_n927), .A4(new_n921), .ZN(new_n928));
  INV_X1    g503(.A(new_n924), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n894), .A2(new_n923), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n921), .B1(new_n929), .B2(new_n930), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n920), .A2(KEYINPUT43), .A3(new_n924), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(G397));
  INV_X1    g514(.A(KEYINPUT126), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n768), .A2(G2067), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n478), .A2(G2105), .ZN(new_n943));
  INV_X1    g518(.A(G126), .ZN(new_n944));
  OAI22_X1  g519(.A1(new_n943), .A2(new_n944), .B1(new_n491), .B2(new_n492), .ZN(new_n945));
  INV_X1    g520(.A(new_n500), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n499), .B1(new_n478), .B2(new_n496), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT99), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n498), .A2(new_n840), .A3(new_n500), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n942), .B1(new_n950), .B2(G1384), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n475), .A2(G40), .A3(new_n481), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G2067), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n768), .B(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT112), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(new_n845), .A3(G1996), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n843), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n475), .A2(G40), .A3(new_n481), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT111), .B1(new_n964), .B2(G1996), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n966));
  INV_X1    g541(.A(G1996), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n953), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(new_n738), .A3(new_n735), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n960), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n703), .A2(new_n706), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n941), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n703), .B(new_n706), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n953), .A2(new_n974), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n960), .A2(new_n975), .A3(new_n970), .ZN(new_n976));
  INV_X1    g551(.A(G1986), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n953), .A2(new_n696), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT48), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n973), .A2(new_n953), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n969), .B(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n953), .B1(new_n956), .B2(new_n845), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT125), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(KEYINPUT125), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n986), .A2(KEYINPUT47), .A3(new_n987), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n980), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n950), .A2(G1384), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(new_n963), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n688), .A2(G1976), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n963), .A2(new_n843), .A3(new_n961), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(G8), .A3(new_n997), .A4(new_n999), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT114), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1005), .B(new_n575), .C1(new_n582), .C2(new_n583), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n581), .A2(G651), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n510), .A2(G48), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT115), .B(G86), .Z(new_n1009));
  NAND2_X1  g584(.A1(new_n523), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G1981), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT116), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1006), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1001), .A2(new_n1015), .A3(G8), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(KEYINPUT116), .A3(new_n1013), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1001), .A2(G8), .A3(new_n997), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1016), .A2(new_n1018), .B1(KEYINPUT52), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1004), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G303), .A2(G8), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n952), .B1(new_n994), .B2(KEYINPUT45), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n502), .A2(new_n961), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n942), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1971), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n950), .B2(G1384), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n494), .B2(new_n501), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT50), .ZN(new_n1032));
  AOI211_X1 g607(.A(G2090), .B(new_n952), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(G8), .B(new_n1024), .C1(new_n1028), .C2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT113), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n843), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(new_n963), .A3(new_n1027), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n685), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT50), .B1(new_n843), .B2(new_n961), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1032), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n963), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1038), .B1(G2090), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(G8), .A4(new_n1024), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1035), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n952), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n725), .C1(new_n994), .C2(new_n1029), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n993), .B1(new_n1038), .B2(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1048), .A2(new_n1024), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n952), .B1(KEYINPUT45), .B2(new_n1031), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1966), .B1(new_n951), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n963), .A2(new_n743), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1053));
  OAI21_X1  g628(.A(G8), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1054), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1021), .B1(new_n1045), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n963), .B1(new_n1026), .B2(new_n942), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n962), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n952), .A2(G2084), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n993), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1004), .A2(new_n1020), .A3(new_n569), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1024), .B1(new_n1042), .B2(G8), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT63), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n995), .B(KEYINPUT117), .ZN(new_n1067));
  AOI211_X1 g642(.A(G1976), .B(G288), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1006), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1057), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n531), .A2(G8), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT122), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1054), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT121), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1060), .A2(new_n1062), .A3(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1079), .A3(G8), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1074), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1077), .A2(new_n1079), .A3(new_n1074), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1084));
  OAI211_X1 g659(.A(KEYINPUT62), .B(new_n1076), .C1(new_n1082), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G2078), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n951), .A2(new_n1050), .A3(KEYINPUT123), .A4(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1087), .A2(KEYINPUT53), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n951), .A2(new_n1050), .A3(new_n1086), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1088), .A2(new_n1091), .B1(new_n727), .B2(new_n1041), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1036), .A2(new_n1086), .A3(new_n1027), .A4(new_n963), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT124), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(KEYINPUT124), .A3(new_n1094), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G301), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1004), .B(new_n1020), .C1(new_n1048), .C2(new_n1024), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1035), .B2(new_n1044), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1085), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(KEYINPUT51), .A3(new_n1083), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT62), .B1(new_n1104), .B2(new_n1076), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1072), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n559), .B(KEYINPUT57), .C1(new_n565), .C2(new_n566), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n558), .A2(G651), .ZN(new_n1109));
  INV_X1    g684(.A(new_n555), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT73), .B1(new_n523), .B2(G91), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n561), .A2(new_n564), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1108), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1107), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1029), .B1(new_n843), .B2(new_n961), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n963), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n808), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1036), .A2(new_n963), .A3(new_n1027), .A4(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1116), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1119), .A2(new_n1121), .A3(new_n1116), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n994), .A2(new_n954), .A3(new_n963), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n952), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT60), .B(new_n1127), .C1(new_n1128), .C2(G1348), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1125), .A2(new_n1126), .B1(new_n1130), .B2(new_n597), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1036), .A2(new_n967), .A3(new_n1027), .A4(new_n963), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1001), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n546), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT59), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1138), .A3(new_n546), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1127), .B1(new_n1128), .B2(G1348), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(new_n607), .A3(new_n1129), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1116), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1107), .A2(new_n1115), .A3(KEYINPUT119), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT61), .B(new_n1124), .C1(new_n1145), .C2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1131), .A2(new_n1140), .A3(new_n1144), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1141), .A2(new_n607), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n1124), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT120), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1086), .A2(KEYINPUT53), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n843), .A2(new_n961), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(new_n942), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1041), .A2(new_n727), .B1(new_n1025), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1093), .A2(KEYINPUT124), .A3(new_n1094), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1160), .B(G301), .C1(new_n1161), .C2(new_n1095), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1156), .B1(new_n1099), .B2(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1165), .A2(new_n1103), .B1(new_n1054), .B2(new_n1075), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1160), .B1(new_n1161), .B2(new_n1095), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1156), .B1(new_n1167), .B2(G171), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1092), .A2(new_n1098), .A3(G301), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1164), .A2(new_n1166), .A3(new_n1170), .A4(new_n1101), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1155), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1140), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1119), .A2(new_n1121), .A3(new_n1116), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1126), .B1(new_n1174), .B2(new_n1122), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1130), .A2(new_n597), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(KEYINPUT120), .B(new_n1154), .C1(new_n1173), .C2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1106), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(G290), .B(new_n977), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n976), .B1(new_n964), .B2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n940), .B(new_n992), .C1(new_n1179), .C2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1035), .A2(new_n1044), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1066), .B(new_n1070), .C1(new_n1183), .C2(new_n1021), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1100), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1045), .A2(new_n1099), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1186), .B1(KEYINPUT62), .B2(new_n1166), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1105), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1184), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AND4_X1   g764(.A1(new_n1170), .A2(new_n1101), .A3(new_n1076), .A4(new_n1104), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1154), .B1(new_n1173), .B2(new_n1177), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT120), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1190), .A2(new_n1193), .A3(new_n1178), .A4(new_n1164), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1181), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n980), .A2(new_n990), .A3(new_n991), .ZN(new_n1196));
  OAI21_X1  g771(.A(KEYINPUT126), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1182), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g773(.A1(G401), .A2(new_n464), .A3(G227), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n677), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g775(.A(new_n1201), .B(KEYINPUT127), .ZN(new_n1202));
  NAND3_X1  g776(.A1(new_n932), .A2(new_n863), .A3(new_n1202), .ZN(G225));
  INV_X1    g777(.A(G225), .ZN(G308));
endmodule


