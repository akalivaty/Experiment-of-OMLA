//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(new_n204), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n213), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n216), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G200), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  OR3_X1    g0055(.A1(new_n254), .A2(KEYINPUT66), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT66), .B1(new_n254), .B2(new_n255), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n258), .A2(G223), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n254), .A2(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G222), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n249), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  OAI211_X1 g0066(.A(G1), .B(G13), .C1(new_n250), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G274), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n249), .A2(new_n270), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(G226), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n248), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT9), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n209), .B1(new_n213), .B2(new_n250), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n210), .B1(new_n201), .B2(new_n203), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n250), .A2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n279), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n277), .B1(new_n278), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  INV_X1    g0087(.A(G1), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G13), .A3(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n291), .A2(new_n288), .A3(G13), .A4(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(new_n277), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n288), .A2(G20), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G50), .A3(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n287), .B(new_n297), .C1(G50), .C2(new_n293), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n275), .B1(new_n276), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n265), .A2(new_n274), .ZN(new_n303));
  OR3_X1    g0103(.A1(new_n298), .A2(new_n276), .A3(new_n299), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n301), .B1(new_n302), .B2(new_n303), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT10), .B1(new_n275), .B2(KEYINPUT73), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT77), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n251), .A2(new_n253), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n250), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n210), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT7), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n311), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n312), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n315), .A2(KEYINPUT78), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT78), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n313), .A2(new_n318), .A3(new_n314), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G68), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT79), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n315), .A2(KEYINPUT78), .A3(new_n316), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT79), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(G68), .A4(new_n319), .ZN(new_n324));
  INV_X1    g0124(.A(G58), .ZN(new_n325));
  INV_X1    g0125(.A(G68), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(G20), .B1(new_n327), .B2(new_n203), .ZN(new_n328));
  INV_X1    g0128(.A(G159), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(KEYINPUT80), .B1(new_n329), .B2(new_n284), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n328), .A2(KEYINPUT80), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n321), .A2(KEYINPUT16), .A3(new_n324), .A4(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n314), .B1(new_n263), .B2(G20), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(G68), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT16), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n277), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n333), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n279), .B1(new_n288), .B2(G20), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n295), .A2(new_n343), .B1(new_n294), .B2(new_n279), .ZN(new_n344));
  INV_X1    g0144(.A(G274), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n249), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n270), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n273), .A2(G232), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n250), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n263), .B2(new_n310), .ZN(new_n351));
  INV_X1    g0151(.A(G226), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G223), .B2(G1698), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n351), .A2(new_n354), .B1(new_n250), .B2(new_n218), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n349), .B1(new_n249), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n248), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(G190), .B2(new_n356), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n342), .A2(new_n344), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT17), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n344), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n333), .B2(new_n341), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(KEYINPUT17), .A3(new_n358), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n342), .A2(new_n344), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT81), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(KEYINPUT81), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n355), .A2(new_n249), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n347), .A3(new_n348), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G169), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n356), .A2(G179), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n368), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n365), .B1(KEYINPUT18), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT81), .B1(new_n342), .B2(new_n344), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n367), .B(new_n362), .C1(new_n333), .C2(new_n341), .ZN(new_n378));
  INV_X1    g0178(.A(new_n374), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n347), .A2(KEYINPUT74), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT74), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n272), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT13), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G226), .A2(G1698), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n233), .B2(G1698), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n390), .A2(new_n263), .B1(G33), .B2(G97), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(new_n267), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n273), .A2(G238), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n387), .A2(new_n388), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n385), .B1(new_n346), .B2(new_n270), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n268), .A2(KEYINPUT74), .A3(new_n271), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n393), .B1(new_n391), .B2(new_n267), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT13), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n394), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n387), .A2(new_n393), .A3(new_n392), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(KEYINPUT75), .A3(KEYINPUT13), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(G169), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT14), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT76), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(KEYINPUT76), .A3(KEYINPUT14), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT14), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n401), .A2(new_n403), .A3(new_n410), .A4(G169), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n394), .A2(G179), .A3(new_n400), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n281), .A2(new_n262), .B1(new_n210), .B2(G68), .ZN(new_n416));
  INV_X1    g0216(.A(G50), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n284), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n277), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT11), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n294), .A2(new_n326), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT12), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n295), .A2(G68), .A3(new_n296), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n302), .B1(new_n402), .B2(KEYINPUT13), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n426), .B2(new_n394), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n401), .A2(G200), .A3(new_n403), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G169), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n303), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G179), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n265), .A2(new_n433), .A3(new_n274), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n300), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n435), .B(KEYINPUT69), .ZN(new_n436));
  INV_X1    g0236(.A(G238), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n256), .B2(new_n257), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT70), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n260), .A2(G232), .B1(G107), .B2(new_n254), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n441), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT70), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n249), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n272), .B1(G244), .B2(new_n273), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G200), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n295), .A2(G77), .A3(new_n296), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT71), .ZN(new_n450));
  INV_X1    g0250(.A(new_n279), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT15), .B(G87), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n452), .B1(new_n281), .B2(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n454), .A2(new_n277), .B1(new_n262), .B2(new_n294), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n448), .B(new_n457), .C1(new_n302), .C2(new_n447), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n447), .A2(new_n431), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n445), .A2(new_n433), .A3(new_n446), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n436), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NOR4_X1   g0262(.A1(new_n309), .A2(new_n383), .A3(new_n430), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT6), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n464), .A2(new_n220), .A3(G107), .ZN(new_n465));
  XNOR2_X1  g0265(.A(G97), .B(G107), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  OAI22_X1  g0267(.A1(new_n467), .A2(new_n210), .B1(new_n262), .B2(new_n284), .ZN(new_n468));
  INV_X1    g0268(.A(G107), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n334), .B2(new_n336), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n277), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n294), .A2(new_n220), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n311), .A2(new_n312), .ZN(new_n474));
  INV_X1    g0274(.A(G244), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1698), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT4), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT4), .A2(G244), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n263), .A2(new_n255), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n249), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n269), .A2(G1), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n267), .A3(G274), .A4(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G257), .A3(new_n267), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n490), .A2(KEYINPUT83), .A3(G257), .A4(new_n267), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n483), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n288), .A2(G33), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n293), .A2(new_n340), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n293), .A2(new_n340), .A3(KEYINPUT82), .A4(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(G97), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n483), .A2(new_n495), .A3(G190), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n473), .A2(new_n497), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n496), .A2(new_n431), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n471), .A2(new_n503), .A3(new_n472), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n507), .C1(G179), .C2(new_n496), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n437), .A2(new_n255), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n475), .A2(G1698), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n311), .B2(new_n312), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G116), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT84), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT84), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n515), .C1(new_n351), .C2(new_n513), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n519), .A3(new_n249), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n249), .A2(new_n219), .A3(new_n485), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n346), .B2(new_n485), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT85), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT85), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n520), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n433), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n474), .A2(new_n210), .A3(G68), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT19), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n281), .B2(new_n220), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n210), .A2(new_n532), .B1(new_n533), .B2(new_n218), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT86), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n277), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n294), .A2(new_n453), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n501), .A2(new_n502), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n453), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n520), .A2(new_n525), .A3(new_n522), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n525), .B1(new_n520), .B2(new_n522), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n527), .B(new_n539), .C1(new_n542), .C2(G169), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n524), .A2(G190), .A3(new_n526), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n501), .A2(G87), .A3(new_n502), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n536), .A2(new_n537), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n544), .B(new_n547), .C1(new_n542), .C2(new_n248), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n510), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n221), .A2(new_n255), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G264), .B2(new_n255), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n312), .B2(new_n311), .ZN(new_n553));
  INV_X1    g0353(.A(G303), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n263), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n249), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n490), .A2(G270), .A3(new_n267), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n486), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G116), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n294), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n293), .A2(new_n340), .A3(G116), .A4(new_n498), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n481), .B(new_n210), .C1(G33), .C2(new_n220), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(G20), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n277), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT20), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n562), .B(new_n563), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n560), .A2(new_n570), .A3(G169), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n560), .A2(new_n433), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n570), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n560), .A2(new_n570), .A3(KEYINPUT21), .A4(G169), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n560), .A2(G200), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n351), .A2(new_n552), .B1(new_n554), .B2(new_n263), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n558), .B1(new_n579), .B2(new_n249), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  INV_X1    g0381(.A(new_n570), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT87), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n578), .A2(new_n581), .A3(KEYINPUT87), .A4(new_n582), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n577), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n255), .A2(G250), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT89), .B1(new_n351), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g0389(.A1(KEYINPUT90), .A2(G294), .ZN(new_n590));
  NAND2_X1  g0390(.A1(KEYINPUT90), .A2(G294), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n250), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n221), .A2(new_n255), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(new_n474), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT89), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n474), .A2(new_n595), .A3(G250), .A4(new_n255), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n589), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n249), .B1(new_n485), .B2(new_n484), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n249), .B1(G264), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT91), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(G179), .A4(new_n486), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT24), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n474), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT23), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n210), .B2(G107), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n469), .A2(KEYINPUT23), .A3(G20), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n606), .A2(new_n607), .B1(new_n280), .B2(G116), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n254), .A2(G20), .A3(new_n218), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(KEYINPUT22), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n602), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n609), .A2(KEYINPUT22), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n612), .A2(KEYINPUT24), .A3(new_n603), .A4(new_n608), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n613), .A3(new_n277), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n501), .A2(G107), .A3(new_n502), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n290), .A2(new_n469), .A3(new_n292), .ZN(new_n616));
  XOR2_X1   g0416(.A(new_n616), .B(KEYINPUT25), .Z(new_n617));
  INV_X1    g0417(.A(KEYINPUT88), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n615), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n614), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n599), .A2(G179), .A3(new_n486), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT91), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n431), .B1(new_n599), .B2(new_n486), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n601), .B(new_n621), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n599), .A2(G190), .A3(new_n486), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n597), .A2(new_n249), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n598), .A2(G264), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n628), .A2(new_n486), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n627), .B1(new_n630), .B2(new_n248), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(new_n621), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n463), .A2(new_n550), .A3(new_n587), .A4(new_n633), .ZN(G372));
  INV_X1    g0434(.A(new_n577), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(new_n635), .B2(new_n625), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n248), .B1(new_n520), .B2(new_n522), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n546), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT92), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT92), .B1(new_n546), .B2(new_n637), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n544), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n523), .A2(new_n431), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n527), .A2(new_n539), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n636), .A2(new_n645), .A3(new_n510), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  INV_X1    g0447(.A(new_n508), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n644), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n543), .A2(new_n548), .A3(new_n648), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(KEYINPUT26), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n646), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n463), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n436), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n363), .A2(new_n379), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n381), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT18), .B1(new_n363), .B2(new_n379), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n461), .A2(KEYINPUT93), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT93), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n459), .A2(new_n662), .A3(new_n456), .A4(new_n460), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n429), .A3(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n425), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n660), .B1(new_n665), .B2(new_n365), .ZN(new_n666));
  INV_X1    g0466(.A(new_n309), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n655), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n654), .A2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n288), .A2(new_n210), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n570), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n587), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n635), .B2(new_n676), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n675), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n626), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n621), .A2(new_n675), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n625), .B1(new_n632), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT94), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n635), .A2(new_n675), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n633), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(new_n681), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  NAND3_X1  g0492(.A1(new_n533), .A2(new_n218), .A3(new_n561), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n214), .A2(new_n266), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(G1), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n207), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n524), .A2(new_n526), .ZN(new_n700));
  INV_X1    g0500(.A(new_n496), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n599), .A3(new_n574), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n699), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n628), .A2(new_n629), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n580), .A2(new_n483), .A3(new_n495), .A4(G179), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n542), .A2(new_n706), .A3(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n599), .A2(new_n486), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n580), .A2(G179), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n708), .A2(new_n496), .A3(new_n523), .A4(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n703), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n675), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n619), .A2(new_n620), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n708), .A2(G200), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n614), .A3(new_n627), .A4(new_n718), .ZN(new_n719));
  AND4_X1   g0519(.A1(new_n587), .A2(new_n625), .A3(new_n719), .A4(new_n680), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT95), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(new_n550), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n587), .A2(new_n625), .A3(new_n719), .A4(new_n680), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT95), .B1(new_n723), .B2(new_n549), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n716), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G330), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT96), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n715), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n711), .B2(new_n675), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n721), .B1(new_n720), .B2(new_n550), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n723), .A2(new_n549), .A3(KEYINPUT95), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT96), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(G330), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT98), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n509), .B(new_n737), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n738), .A2(new_n636), .A3(new_n645), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n642), .A2(new_n648), .A3(new_n644), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT26), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n543), .A2(new_n548), .A3(new_n647), .A4(new_n648), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n644), .A3(new_n742), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT29), .B(new_n680), .C1(new_n739), .C2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n653), .A2(new_n680), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n736), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n698), .B1(new_n749), .B2(G1), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT99), .Z(G364));
  AND2_X1   g0551(.A1(new_n210), .A2(G13), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n288), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n695), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n679), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G330), .B2(new_n678), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n756), .B(KEYINPUT100), .Z(new_n759));
  NAND2_X1  g0559(.A1(new_n263), .A2(new_n214), .ZN(new_n760));
  INV_X1    g0560(.A(G355), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(G116), .B2(new_n214), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n243), .A2(G45), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n351), .A2(new_n214), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n269), .B2(new_n208), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n209), .B1(G20), .B2(new_n431), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n759), .B1(new_n766), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n210), .A2(new_n433), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n302), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT102), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n590), .A2(new_n591), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n302), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n210), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n778), .A2(G326), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT103), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(KEYINPUT103), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n210), .A2(new_n248), .A3(G179), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n786), .A2(new_n302), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT101), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT101), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G283), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G190), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n793), .A2(G20), .A3(new_n433), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n795), .A2(G311), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G322), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n774), .A2(G190), .A3(new_n248), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n798), .B(new_n254), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n775), .A2(G190), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n786), .A2(G190), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n554), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n784), .A2(new_n785), .A3(new_n792), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(new_n218), .ZN(new_n809));
  INV_X1    g0609(.A(new_n776), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n797), .A2(G159), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n810), .A2(new_n417), .B1(KEYINPUT32), .B2(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n809), .B(new_n812), .C1(G68), .C2(new_n802), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n791), .A2(G107), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n263), .B1(new_n800), .B2(new_n325), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G77), .B2(new_n795), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n781), .A2(new_n220), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(KEYINPUT32), .B2(new_n811), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n808), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n773), .B1(new_n820), .B2(new_n770), .ZN(new_n821));
  INV_X1    g0621(.A(new_n769), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n678), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n758), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NAND4_X1  g0625(.A1(new_n661), .A2(new_n456), .A3(new_n663), .A4(new_n675), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n458), .B(new_n461), .C1(new_n457), .C2(new_n680), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n745), .B(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n756), .B1(new_n829), .B2(new_n736), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n736), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n770), .A2(new_n767), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT104), .Z(new_n833));
  OAI21_X1  g0633(.A(new_n759), .B1(new_n833), .B2(G77), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n803), .A2(KEYINPUT105), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n803), .A2(KEYINPUT105), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(G283), .ZN(new_n839));
  INV_X1    g0639(.A(G294), .ZN(new_n840));
  INV_X1    g0640(.A(G311), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n800), .A2(new_n840), .B1(new_n841), .B2(new_n796), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n263), .B(new_n842), .C1(G116), .C2(new_n795), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n805), .A2(new_n469), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n817), .B(new_n844), .C1(G303), .C2(new_n776), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n791), .A2(G87), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n839), .A2(new_n843), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n800), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G143), .B1(new_n795), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n803), .B2(new_n282), .C1(new_n850), .C2(new_n810), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n791), .A2(G68), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n805), .A2(new_n417), .B1(new_n781), .B2(new_n325), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n351), .B(new_n856), .C1(G132), .C2(new_n797), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n847), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n834), .B1(new_n859), .B2(new_n770), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n828), .B2(new_n768), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n831), .A2(new_n861), .ZN(G384));
  INV_X1    g0662(.A(KEYINPUT107), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n333), .A2(new_n277), .ZN(new_n864));
  INV_X1    g0664(.A(new_n332), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n322), .A2(G68), .A3(new_n319), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n866), .B2(KEYINPUT79), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT16), .B1(new_n867), .B2(new_n324), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n344), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n673), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n376), .B2(new_n382), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n359), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n377), .A2(new_n378), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n875), .B1(new_n876), .B2(new_n374), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n368), .A2(new_n369), .A3(new_n870), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n869), .A2(new_n374), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n871), .A2(new_n879), .A3(new_n359), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n877), .A2(new_n878), .B1(new_n880), .B2(KEYINPUT37), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n872), .A2(new_n873), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n871), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n363), .A2(KEYINPUT17), .A3(new_n358), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT17), .B1(new_n363), .B2(new_n358), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n380), .B2(new_n381), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n375), .A2(KEYINPUT18), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n883), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n375), .A2(new_n878), .A3(new_n874), .A4(new_n359), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n863), .B1(new_n882), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n873), .B1(new_n872), .B2(new_n881), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(KEYINPUT107), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n429), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n424), .B(new_n675), .C1(new_n415), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n424), .A2(new_n675), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n413), .B1(new_n407), .B2(new_n408), .ZN(new_n902));
  INV_X1    g0702(.A(new_n424), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n429), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n733), .A2(new_n905), .A3(new_n828), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT40), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n377), .A2(new_n378), .A3(new_n673), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n659), .B2(new_n365), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n380), .A2(new_n908), .A3(new_n875), .ZN(new_n910));
  INV_X1    g0710(.A(new_n359), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n656), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n874), .B1(new_n878), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n909), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n873), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n896), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n733), .A2(new_n905), .A3(KEYINPUT40), .A4(new_n828), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n907), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n463), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(new_n725), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n919), .A2(new_n921), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n922), .A2(new_n923), .A3(new_n726), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n653), .A2(new_n680), .A3(new_n828), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n461), .A2(new_n675), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n905), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n895), .A2(KEYINPUT107), .A3(new_n896), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT107), .B1(new_n895), .B2(new_n896), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n878), .A2(new_n912), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n890), .B1(new_n935), .B2(new_n874), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n936), .B2(new_n909), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n882), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n415), .A2(new_n424), .A3(new_n680), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n660), .A2(new_n870), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n933), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n463), .B(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n668), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n945), .B(new_n947), .Z(new_n948));
  OAI22_X1  g0748(.A1(new_n924), .A2(new_n948), .B1(new_n288), .B2(new_n752), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n924), .ZN(new_n950));
  INV_X1    g0750(.A(new_n467), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(KEYINPUT35), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n952), .A2(G116), .A3(new_n211), .A4(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT36), .Z(new_n955));
  NOR3_X1   g0755(.A1(new_n207), .A2(new_n262), .A3(new_n327), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT106), .B1(new_n201), .B2(G68), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n201), .A2(KEYINPUT106), .A3(G68), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n288), .B(G13), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n950), .A2(new_n955), .A3(new_n960), .ZN(G367));
  OAI221_X1 g0761(.A(new_n771), .B1(new_n214), .B2(new_n453), .C1(new_n239), .C2(new_n764), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n759), .A2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n838), .A2(G159), .B1(G143), .B2(new_n778), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n791), .A2(G77), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n800), .A2(new_n282), .B1(new_n850), .B2(new_n796), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n254), .B(new_n966), .C1(new_n202), .C2(new_n795), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n781), .A2(new_n326), .ZN(new_n968));
  INV_X1    g0768(.A(new_n805), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(G58), .B2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n964), .A2(new_n965), .A3(new_n967), .A4(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n790), .A2(new_n220), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n474), .B(new_n972), .C1(G317), .C2(new_n797), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT112), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n969), .A2(KEYINPUT46), .A3(G116), .ZN(new_n976));
  INV_X1    g0776(.A(G283), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n800), .A2(new_n554), .B1(new_n794), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT46), .B1(new_n969), .B2(G116), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(G107), .C2(new_n782), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n838), .A2(new_n779), .B1(G311), .B2(new_n778), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n975), .A2(new_n976), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n973), .A2(new_n974), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n971), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n963), .B1(new_n985), .B2(new_n770), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n546), .A2(new_n675), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n645), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n644), .A2(new_n987), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n769), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n507), .A2(new_n675), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n738), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n648), .A2(new_n675), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n691), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n997), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n690), .A2(new_n681), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n691), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n687), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n687), .B1(new_n1008), .B2(new_n1004), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n679), .A2(KEYINPUT110), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n690), .B1(new_n684), .B2(new_n689), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1013), .B(new_n1014), .Z(new_n1015));
  NAND2_X1  g0815(.A1(new_n749), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT111), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n688), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n1009), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT111), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1020), .A2(new_n1021), .A3(new_n749), .A4(new_n1015), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n749), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n695), .B(KEYINPUT41), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n754), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT42), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n1001), .B2(new_n690), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n997), .A2(KEYINPUT42), .A3(new_n633), .A4(new_n689), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n508), .B1(new_n995), .B2(new_n625), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1029), .A2(new_n1030), .B1(new_n680), .B2(new_n1031), .ZN(new_n1032));
  OR3_X1    g0832(.A1(new_n1032), .A2(KEYINPUT108), .A3(new_n991), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n991), .B1(new_n1032), .B2(KEYINPUT108), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT43), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  AND3_X1   g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT43), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n688), .A2(new_n1001), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n993), .B1(new_n1027), .B2(new_n1041), .ZN(G387));
  NAND2_X1  g0842(.A1(new_n1015), .A2(new_n754), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n760), .A2(new_n694), .B1(G107), .B2(new_n214), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n236), .A2(new_n269), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n279), .A2(G50), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT50), .ZN(new_n1047));
  AOI211_X1 g0847(.A(G45), .B(new_n693), .C1(G68), .C2(G77), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n764), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1044), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT113), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n771), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n759), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n474), .B1(G326), .B2(new_n797), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n779), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n805), .A2(new_n1056), .B1(new_n781), .B2(new_n977), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n848), .A2(G317), .B1(new_n795), .B2(G303), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n799), .B2(new_n777), .C1(new_n837), .C2(new_n841), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT49), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1055), .B1(new_n561), .B2(new_n790), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n781), .A2(new_n453), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n805), .A2(new_n262), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n451), .C2(new_n802), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n800), .A2(new_n417), .B1(new_n794), .B2(new_n326), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G150), .B2(new_n797), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n351), .B1(G159), .B2(new_n776), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1064), .A2(new_n1065), .B1(new_n972), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1054), .B1(new_n1073), .B2(new_n770), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n684), .B2(new_n822), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1016), .A2(new_n755), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n749), .A2(new_n1015), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1043), .B(new_n1075), .C1(new_n1076), .C2(new_n1077), .ZN(G393));
  NOR2_X1   g0878(.A1(new_n781), .A2(new_n262), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n795), .A2(new_n451), .B1(new_n797), .B2(G143), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n474), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(G68), .C2(new_n969), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1082), .B(new_n846), .C1(new_n201), .C2(new_n837), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G150), .A2(new_n776), .B1(new_n848), .B2(G159), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT51), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G317), .A2(new_n776), .B1(new_n848), .B2(G311), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n254), .B1(new_n796), .B2(new_n799), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n805), .A2(new_n977), .B1(new_n781), .B2(new_n561), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G294), .C2(new_n795), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n814), .B(new_n1090), .C1(new_n554), .C2(new_n837), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1083), .A2(new_n1085), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n770), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n771), .B1(new_n220), .B2(new_n214), .C1(new_n246), .C2(new_n764), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n759), .A3(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT114), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1001), .B2(new_n769), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1020), .B2(new_n754), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT115), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n695), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1023), .A2(KEYINPUT116), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT116), .B1(new_n1023), .B2(new_n1100), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(G390));
  AND4_X1   g0904(.A1(G330), .A2(new_n733), .A3(new_n905), .A4(new_n828), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n938), .A2(new_n941), .B1(new_n939), .B2(new_n929), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n828), .B(new_n680), .C1(new_n739), .C2(new_n743), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n927), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n905), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n916), .A3(new_n939), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1105), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n929), .A2(new_n939), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n1114));
  AOI21_X1  g0914(.A(KEYINPUT39), .B1(new_n915), .B2(new_n896), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n727), .A2(new_n735), .A3(new_n828), .A4(new_n905), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1110), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n753), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n767), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n759), .B1(new_n833), .B2(new_n451), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT117), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n838), .A2(G107), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n800), .A2(new_n561), .B1(new_n794), .B2(new_n220), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n263), .B(new_n1125), .C1(G294), .C2(new_n797), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1079), .B(new_n809), .C1(G283), .C2(new_n776), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1124), .A2(new_n855), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n805), .A2(new_n282), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT119), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT118), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  INV_X1    g0933(.A(G125), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n794), .A2(new_n1133), .B1(new_n796), .B2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n254), .B(new_n1135), .C1(G132), .C2(new_n848), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G159), .A2(new_n782), .B1(new_n776), .B2(G128), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n850), .B2(new_n837), .C1(new_n201), .C2(new_n790), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1128), .B1(new_n1132), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1123), .B1(new_n1140), .B2(new_n770), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1120), .B1(new_n1121), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n733), .A2(G330), .A3(new_n828), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n905), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1108), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1117), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n727), .A2(new_n735), .A3(new_n828), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1105), .B1(new_n1147), .B2(new_n1144), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n928), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n725), .A2(new_n726), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n463), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1152), .B(new_n668), .C1(new_n920), .C2(new_n747), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1119), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1112), .A2(new_n1118), .A3(new_n1150), .A4(new_n1154), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n755), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1142), .A2(new_n1158), .ZN(G378));
  AOI21_X1  g0959(.A(new_n943), .B1(new_n898), .B2(new_n930), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n882), .A2(new_n937), .ZN(new_n1161));
  OAI21_X1  g0961(.A(G330), .B1(new_n1161), .B2(new_n917), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n942), .B(new_n1160), .C1(new_n907), .C2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n906), .B1(new_n931), .B2(new_n932), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT40), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1162), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n945), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT121), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n667), .A2(new_n1168), .A3(new_n435), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n435), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT121), .B1(new_n309), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n300), .A2(new_n870), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT55), .Z(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1174), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1169), .A2(new_n1177), .A3(new_n1171), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1176), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1163), .A2(new_n1167), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1181), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1157), .A2(new_n1154), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT57), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1181), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1157), .B2(new_n1154), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1163), .A2(new_n1167), .A3(new_n1181), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1189), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n755), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1186), .A2(new_n1194), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n755), .B(new_n754), .C1(new_n201), .C2(new_n832), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n770), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n791), .A2(G58), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n220), .A2(new_n803), .B1(new_n810), .B2(new_n561), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1199), .A2(new_n968), .A3(new_n1067), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n794), .A2(new_n453), .B1(new_n796), .B2(new_n977), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n351), .A2(new_n266), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G107), .C2(new_n848), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1198), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT58), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1202), .B(new_n417), .C1(G33), .C2(G41), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G132), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n803), .A2(new_n1210), .B1(new_n805), .B2(new_n1133), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n848), .A2(G128), .B1(new_n795), .B2(G137), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n282), .B2(new_n781), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(G125), .C2(new_n776), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT120), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n797), .C2(G124), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n790), .B2(new_n329), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1215), .B2(KEYINPUT59), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1206), .B(new_n1209), .C1(new_n1216), .C2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1196), .B1(new_n1197), .B2(new_n1220), .C1(new_n1181), .C2(new_n768), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1184), .B2(new_n754), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1195), .A2(new_n1223), .ZN(G375));
  OAI211_X1 g1024(.A(new_n1153), .B(new_n1146), .C1(new_n1149), .C2(new_n1148), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1155), .A2(new_n1026), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1144), .A2(new_n767), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n759), .B1(new_n833), .B2(G68), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n810), .A2(new_n1210), .B1(new_n850), .B2(new_n800), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1133), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(new_n838), .B2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT124), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n969), .A2(G159), .B1(new_n782), .B2(G50), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n795), .A2(G150), .B1(new_n797), .B2(G128), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1233), .A2(new_n474), .A3(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(new_n1198), .A3(new_n1235), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n810), .A2(new_n840), .B1(new_n794), .B2(new_n469), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n838), .B2(G116), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT123), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n254), .B1(new_n796), .B2(new_n554), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G283), .B2(new_n848), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1066), .B1(G97), .B2(new_n969), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n965), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1236), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1228), .B1(new_n1244), .B2(new_n770), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT125), .Z(new_n1246));
  AOI22_X1  g1046(.A1(new_n1150), .A2(new_n754), .B1(new_n1227), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1226), .A2(new_n1247), .ZN(G381));
  INV_X1    g1048(.A(new_n1040), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1039), .B(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n748), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n753), .B1(new_n1251), .B2(new_n1025), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1250), .A2(new_n1252), .B1(new_n992), .B2(new_n986), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1099), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1103), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(new_n1101), .ZN(new_n1256));
  INV_X1    g1056(.A(G381), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1253), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OR3_X1    g1059(.A1(G375), .A2(G378), .A3(new_n1259), .ZN(G407));
  INV_X1    g1060(.A(G378), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n674), .A2(G213), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G407), .B(G213), .C1(G375), .C2(new_n1264), .ZN(G409));
  INV_X1    g1065(.A(KEYINPUT61), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G378), .B(new_n1223), .C1(new_n1186), .C2(new_n1194), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1189), .A2(new_n1026), .A3(new_n1185), .A4(new_n1192), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1189), .A2(new_n754), .A3(new_n1192), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1221), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1261), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1263), .B1(new_n1267), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1274), .A2(KEYINPUT60), .A3(new_n1153), .A4(new_n1146), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1225), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1275), .A2(new_n1277), .A3(new_n755), .A4(new_n1155), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1278), .A2(G384), .A3(new_n1247), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1278), .B2(new_n1247), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1273), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1247), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1278), .A2(G384), .A3(new_n1247), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(KEYINPUT126), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1263), .A2(G2897), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1281), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(G2897), .A3(new_n1263), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1266), .B1(new_n1272), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1281), .A2(new_n1286), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1272), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(G393), .B(new_n824), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(new_n1256), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1253), .A2(G390), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1299), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  AOI211_X1 g1104(.A(KEYINPUT127), .B(new_n1298), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1294), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1293), .A2(new_n1297), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT62), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1272), .A2(new_n1309), .A3(new_n1294), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1272), .B2(new_n1294), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1310), .A2(new_n1292), .A3(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1308), .B1(new_n1312), .B2(new_n1306), .ZN(G405));
  NOR2_X1   g1113(.A1(G387), .A2(new_n1256), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1253), .A2(G390), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1303), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1298), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1302), .A2(new_n1303), .A3(new_n1299), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G375), .A2(new_n1261), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(new_n1267), .A3(new_n1289), .ZN(new_n1321));
  AOI21_X1  g1121(.A(G378), .B1(new_n1195), .B2(new_n1223), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1267), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1294), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1319), .A2(new_n1321), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1319), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(G402));
endmodule


