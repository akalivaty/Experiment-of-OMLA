//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n207), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n208), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT27), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G183gat), .ZN(new_n221));
  INV_X1    g020(.A(G190gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT28), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT28), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n222), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n215), .A2(new_n217), .A3(new_n224), .A4(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n218), .A2(new_n222), .ZN(new_n230));
  NAND3_X1  g029(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT65), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT65), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n240));
  NAND2_X1  g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(G169gat), .B2(G176gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n229), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n240), .A2(KEYINPUT25), .A3(new_n243), .A4(new_n241), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n233), .B1(KEYINPUT66), .B2(KEYINPUT24), .ZN(new_n248));
  AND2_X1   g047(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n247), .B1(new_n250), .B2(new_n232), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n228), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT74), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT74), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n228), .B(new_n254), .C1(new_n246), .C2(new_n251), .ZN(new_n255));
  AND2_X1   g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT29), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(G211gat), .A2(G218gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT22), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT73), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G211gat), .B(G218gat), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n264), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n232), .B1(new_n249), .B2(new_n248), .ZN(new_n271));
  INV_X1    g070(.A(new_n247), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n230), .A2(new_n231), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(new_n235), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n244), .B1(new_n275), .B2(new_n238), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n273), .B1(new_n276), .B2(new_n229), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(new_n256), .A3(new_n228), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n270), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n255), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n254), .B1(new_n277), .B2(new_n228), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n256), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n252), .A2(new_n257), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n270), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n206), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n206), .A2(KEYINPUT37), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n253), .A2(new_n255), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n289), .A2(new_n256), .B1(new_n252), .B2(new_n257), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n279), .B1(new_n290), .B2(new_n270), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT37), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n202), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n279), .B(new_n205), .C1(new_n290), .C2(new_n270), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n206), .B1(new_n291), .B2(KEYINPUT37), .ZN(new_n295));
  INV_X1    g094(.A(new_n270), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n258), .A2(new_n296), .A3(new_n278), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT37), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n202), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n294), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n304));
  INV_X1    g103(.A(G113gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(G120gat), .ZN(new_n306));
  INV_X1    g105(.A(G134gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G127gat), .ZN(new_n308));
  INV_X1    g107(.A(G127gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G134gat), .ZN(new_n310));
  AND4_X1   g109(.A1(new_n303), .A2(new_n306), .A3(new_n308), .A4(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G113gat), .B(G120gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT68), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n305), .A2(G120gat), .ZN(new_n315));
  INV_X1    g114(.A(G120gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(G113gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n303), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n308), .A2(new_n310), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G141gat), .B(G148gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(G155gat), .B2(G162gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G148gat), .ZN(new_n330));
  INV_X1    g129(.A(G148gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G141gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G155gat), .B(G162gat), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT2), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n328), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n321), .B1(KEYINPUT3), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n328), .A2(new_n338), .A3(KEYINPUT75), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT75), .B1(new_n328), .B2(new_n338), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT3), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g144(.A(KEYINPUT76), .B(KEYINPUT3), .C1(new_n341), .C2(new_n342), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n311), .A2(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n328), .A3(new_n338), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n347), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n321), .B1(new_n341), .B2(new_n342), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n356), .B2(new_n349), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT5), .B1(new_n357), .B2(KEYINPUT77), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n328), .A2(new_n338), .A3(KEYINPUT75), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n348), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n321), .A2(new_n339), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n353), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n358), .A2(new_n366), .A3(KEYINPUT78), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n369), .B1(new_n364), .B2(new_n365), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n357), .A2(KEYINPUT77), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n355), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n369), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT0), .ZN(new_n377));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n375), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT78), .B1(new_n358), .B2(new_n366), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n370), .A2(new_n368), .A3(new_n371), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n354), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n354), .A2(new_n369), .ZN(new_n385));
  OAI211_X1 g184(.A(KEYINPUT6), .B(new_n380), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT80), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n379), .A3(new_n374), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n302), .A2(new_n381), .A3(new_n388), .A4(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n347), .A2(new_n351), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n352), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT39), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n380), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n356), .A2(new_n352), .A3(new_n349), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT39), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n399), .A2(KEYINPUT86), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(KEYINPUT86), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n400), .B(new_n401), .C1(new_n352), .C2(new_n394), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n397), .A2(new_n402), .A3(KEYINPUT40), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT40), .B1(new_n397), .B2(new_n402), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OR3_X1    g204(.A1(new_n291), .A2(KEYINPUT30), .A3(new_n206), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n286), .A2(KEYINPUT30), .A3(new_n294), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT85), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT85), .B1(new_n406), .B2(new_n407), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n405), .B(new_n390), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n263), .A2(new_n268), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n266), .A2(new_n262), .A3(new_n259), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT81), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(new_n263), .B2(new_n268), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT81), .B1(new_n417), .B2(new_n412), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n339), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT82), .B(new_n339), .C1(new_n416), .C2(new_n418), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n413), .B1(new_n339), .B2(KEYINPUT3), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n270), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G22gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n267), .A2(new_n413), .A3(new_n269), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n429), .A2(new_n415), .B1(new_n361), .B2(new_n360), .ZN(new_n430));
  INV_X1    g229(.A(new_n424), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n430), .A2(new_n431), .A3(new_n426), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n427), .A2(new_n428), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT31), .B(G50gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n436), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n432), .B1(new_n425), .B2(new_n426), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT83), .B1(new_n442), .B2(new_n428), .ZN(new_n443));
  INV_X1    g242(.A(new_n440), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT84), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n442), .A2(new_n428), .ZN(new_n446));
  AOI211_X1 g245(.A(G22gat), .B(new_n432), .C1(new_n425), .C2(new_n426), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n441), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n441), .B2(new_n445), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n393), .A2(new_n410), .A3(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n243), .A2(new_n241), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n230), .B(new_n231), .C1(new_n237), .C2(KEYINPUT65), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n233), .A2(new_n234), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT65), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n453), .B(new_n240), .C1(new_n454), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n229), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n458), .A2(new_n459), .B1(new_n271), .B2(new_n272), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n217), .A2(new_n224), .A3(new_n227), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n216), .B1(new_n208), .B2(new_n213), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n321), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G227gat), .ZN(new_n465));
  INV_X1    g264(.A(G233gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n228), .B(new_n348), .C1(new_n246), .C2(new_n251), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n464), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT70), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n472), .B(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n469), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n348), .B1(new_n277), .B2(new_n228), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n467), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT32), .ZN(new_n479));
  XNOR2_X1  g278(.A(G15gat), .B(G43gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT33), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT69), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n482), .B1(new_n478), .B2(KEYINPUT32), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n464), .A2(new_n469), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT33), .B1(new_n489), .B2(new_n467), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n487), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n482), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT32), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n496), .A2(KEYINPUT69), .A3(new_n490), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n475), .B(new_n486), .C1(new_n492), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT72), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n488), .A2(new_n491), .A3(new_n487), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT69), .B1(new_n496), .B2(new_n490), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n485), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(new_n475), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n502), .A2(KEYINPUT72), .A3(new_n475), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT36), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n486), .B1(new_n492), .B2(new_n497), .ZN(new_n507));
  INV_X1    g306(.A(new_n475), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n498), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n406), .A2(new_n407), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n392), .A2(KEYINPUT79), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n389), .A2(new_n390), .A3(new_n516), .A4(new_n391), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n381), .A2(new_n388), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n514), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n452), .B(new_n513), .C1(new_n521), .C2(new_n451), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT35), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n441), .A2(new_n445), .A3(new_n448), .ZN(new_n524));
  INV_X1    g323(.A(new_n448), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n437), .B1(new_n436), .B2(new_n440), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n443), .A2(KEYINPUT84), .A3(new_n444), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n524), .B(new_n528), .C1(new_n504), .C2(new_n505), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n523), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT35), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n392), .A2(new_n381), .A3(new_n388), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n509), .A2(new_n498), .ZN(new_n534));
  AND4_X1   g333(.A1(new_n451), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n522), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT101), .ZN(new_n537));
  NAND2_X1  g336(.A1(G230gat), .A2(G233gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G85gat), .A2(G92gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G99gat), .B(G106gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546));
  INV_X1    g345(.A(G85gat), .ZN(new_n547));
  INV_X1    g346(.A(G92gat), .ZN(new_n548));
  AOI22_X1  g347(.A1(KEYINPUT8), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n542), .A3(new_n543), .ZN(new_n551));
  INV_X1    g350(.A(new_n545), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G64gat), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n554), .A2(G57gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(G57gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  OR2_X1    g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n559), .A2(KEYINPUT92), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n561), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(new_n558), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n558), .B1(new_n555), .B2(new_n556), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n550), .B(new_n553), .C1(new_n564), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n568), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n560), .A2(new_n563), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n551), .A2(new_n552), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n545), .B1(new_n544), .B2(new_n549), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(KEYINPUT98), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n573), .A2(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n571), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT10), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(KEYINPUT99), .A3(new_n582), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n570), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT10), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n539), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n576), .A2(new_n580), .A3(new_n539), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n576), .A2(KEYINPUT100), .A3(new_n580), .A4(new_n539), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n537), .B1(new_n590), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT99), .B1(new_n581), .B2(new_n582), .ZN(new_n600));
  AOI211_X1 g399(.A(new_n584), .B(KEYINPUT10), .C1(new_n576), .C2(new_n580), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n589), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n538), .ZN(new_n603));
  INV_X1    g402(.A(new_n598), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(KEYINPUT101), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n597), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n538), .B(KEYINPUT102), .Z(new_n608));
  AOI21_X1  g407(.A(new_n608), .B1(new_n587), .B2(new_n589), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G43gat), .B(G50gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT87), .B(G29gat), .ZN(new_n615));
  INV_X1    g414(.A(G36gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(G29gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(new_n616), .A3(KEYINPUT14), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT14), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(G29gat), .B2(G36gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(KEYINPUT15), .B(new_n614), .C1(new_n617), .C2(new_n622), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n614), .A2(KEYINPUT15), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n614), .A2(KEYINPUT15), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n624), .B(new_n625), .C1(new_n616), .C2(new_n615), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n622), .B(KEYINPUT88), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT17), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT91), .ZN(new_n630));
  XNOR2_X1  g429(.A(G15gat), .B(G22gat), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n631), .A2(G1gat), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT16), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n633), .B2(G1gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(G8gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT89), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n634), .A2(KEYINPUT90), .ZN(new_n638));
  INV_X1    g437(.A(G8gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(KEYINPUT90), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n632), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n636), .A2(KEYINPUT89), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n630), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n628), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n628), .B(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT91), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n648), .A2(KEYINPUT18), .A3(new_n649), .A4(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n652), .A2(new_n649), .A3(new_n647), .A4(new_n645), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT18), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n646), .A2(new_n628), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n647), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n649), .B(KEYINPUT13), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n653), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G113gat), .B(G141gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G197gat), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT11), .B(G169gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT12), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n666), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n653), .A2(new_n656), .A3(new_n668), .A4(new_n660), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n613), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n646), .B1(KEYINPUT21), .B2(new_n578), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n673));
  NAND3_X1  g472(.A1(new_n572), .A2(new_n571), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G231gat), .A2(G233gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G127gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n672), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G155gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(G183gat), .B(G211gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n678), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(G232gat), .A2(G233gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT94), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n628), .B2(new_n577), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n651), .B2(new_n577), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n692), .A2(KEYINPUT95), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(KEYINPUT95), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(G190gat), .B(G218gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n696), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n693), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n688), .A2(new_n689), .ZN(new_n700));
  XOR2_X1   g499(.A(G134gat), .B(G162gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT96), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n697), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n703), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT97), .Z(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n697), .A2(new_n699), .A3(new_n704), .A4(new_n707), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n671), .A2(new_n686), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n536), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n519), .B1(new_n515), .B2(new_n517), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT103), .B(G1gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1324gat));
  NOR2_X1   g517(.A1(new_n408), .A2(new_n409), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n639), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT16), .B(G8gat), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n713), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT42), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(KEYINPUT42), .B2(new_n723), .ZN(G1325gat));
  NAND3_X1  g524(.A1(new_n509), .A2(KEYINPUT72), .A3(new_n498), .ZN(new_n726));
  INV_X1    g525(.A(new_n505), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n511), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n512), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT104), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n506), .A2(new_n731), .A3(new_n512), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G15gat), .B1(new_n713), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n510), .A2(G15gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n713), .B2(new_n736), .ZN(G1326gat));
  NOR2_X1   g536(.A1(new_n713), .A2(new_n451), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT43), .B(G22gat), .Z(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1327gat));
  NAND4_X1  g539(.A1(new_n711), .A2(new_n613), .A3(new_n670), .A4(new_n686), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n528), .A2(new_n524), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n510), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(new_n533), .A3(new_n532), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n714), .A2(new_n529), .A3(new_n514), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n523), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n741), .B1(new_n746), .B2(new_n522), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n714), .A3(new_n615), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT45), .ZN(new_n749));
  INV_X1    g548(.A(new_n711), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n536), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n685), .B(KEYINPUT105), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n671), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n742), .B1(new_n714), .B2(new_n514), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n757), .A2(new_n452), .A3(new_n732), .A4(new_n730), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n750), .B1(new_n746), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n753), .B(new_n756), .C1(new_n759), .C2(KEYINPUT44), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n715), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n749), .B1(new_n615), .B2(new_n761), .ZN(G1328gat));
  INV_X1    g561(.A(new_n719), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n616), .A3(new_n763), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT46), .Z(new_n765));
  OAI21_X1  g564(.A(G36gat), .B1(new_n760), .B2(new_n719), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1329gat));
  OAI21_X1  g566(.A(G43gat), .B1(new_n760), .B2(new_n734), .ZN(new_n768));
  INV_X1    g567(.A(G43gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n747), .A2(new_n769), .A3(new_n534), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g571(.A(G50gat), .B1(new_n760), .B2(new_n451), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(KEYINPUT106), .B(G50gat), .C1(new_n760), .C2(new_n451), .ZN(new_n776));
  INV_X1    g575(.A(G50gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n747), .A2(new_n777), .A3(new_n742), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n760), .B2(new_n451), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G50gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n760), .A2(new_n782), .A3(new_n451), .ZN(new_n785));
  OAI211_X1 g584(.A(KEYINPUT48), .B(new_n778), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n781), .A2(new_n786), .ZN(G1331gat));
  INV_X1    g586(.A(new_n670), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n750), .A2(new_n788), .A3(new_n685), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n613), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT108), .Z(new_n791));
  NAND2_X1  g590(.A1(new_n746), .A2(new_n758), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n714), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n792), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n719), .ZN(new_n797));
  NOR2_X1   g596(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n798));
  AND2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n797), .B2(new_n798), .ZN(G1333gat));
  INV_X1    g600(.A(G71gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n793), .A2(new_n802), .A3(new_n534), .ZN(new_n803));
  OAI21_X1  g602(.A(G71gat), .B1(new_n796), .B2(new_n734), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(G1334gat));
  NOR2_X1   g606(.A1(new_n796), .A2(new_n451), .ZN(new_n808));
  XOR2_X1   g607(.A(KEYINPUT109), .B(G78gat), .Z(new_n809));
  XNOR2_X1  g608(.A(new_n808), .B(new_n809), .ZN(G1335gat));
  AND4_X1   g609(.A1(new_n757), .A2(new_n452), .A3(new_n732), .A4(new_n730), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n521), .A2(new_n530), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n535), .B1(new_n812), .B2(KEYINPUT35), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n711), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n751), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n670), .A2(new_n685), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT110), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n612), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n815), .A2(new_n816), .A3(new_n753), .A4(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n753), .B(new_n819), .C1(new_n759), .C2(KEYINPUT44), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT111), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n820), .A2(new_n822), .A3(new_n714), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n759), .A2(new_n818), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n759), .A2(KEYINPUT51), .A3(new_n818), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n714), .A2(new_n547), .A3(new_n612), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT112), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n823), .A2(new_n547), .B1(new_n829), .B2(new_n831), .ZN(G1336gat));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833));
  OAI21_X1  g632(.A(G92gat), .B1(new_n821), .B2(new_n719), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n763), .A2(new_n548), .A3(new_n612), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n833), .B(new_n834), .C1(new_n829), .C2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n822), .A3(new_n763), .ZN(new_n837));
  INV_X1    g636(.A(new_n835), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n837), .A2(G92gat), .B1(new_n828), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n839), .B2(new_n833), .ZN(G1337gat));
  NAND3_X1  g639(.A1(new_n820), .A2(new_n822), .A3(new_n733), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n820), .A2(new_n822), .A3(KEYINPUT113), .A4(new_n733), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(G99gat), .A3(new_n844), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n613), .A2(G99gat), .A3(new_n510), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(G1338gat));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n849));
  OAI21_X1  g648(.A(G106gat), .B1(new_n821), .B2(new_n451), .ZN(new_n850));
  OR3_X1    g649(.A1(new_n451), .A2(new_n613), .A3(G106gat), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n849), .B(new_n850), .C1(new_n829), .C2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n826), .B2(new_n827), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n820), .A2(new_n822), .A3(new_n742), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(G106gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n855), .B2(new_n849), .ZN(G1339gat));
  INV_X1    g655(.A(new_n608), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n588), .B2(KEYINPUT10), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n600), .B2(new_n601), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT55), .B1(new_n590), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n602), .A2(new_n862), .A3(new_n857), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n607), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT101), .B1(new_n603), .B2(new_n604), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n537), .B(new_n598), .C1(new_n602), .C2(new_n538), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n861), .A2(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n863), .A2(new_n607), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n603), .A2(KEYINPUT54), .A3(new_n859), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT55), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT114), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n590), .A2(new_n860), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n864), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n868), .A2(KEYINPUT55), .A3(new_n869), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n606), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n877), .A3(new_n670), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n649), .B1(new_n648), .B2(new_n652), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n658), .A2(new_n659), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n665), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n612), .A2(new_n669), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n711), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n669), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n709), .B2(new_n710), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n871), .A3(new_n877), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n754), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n789), .A2(new_n612), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n715), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n788), .A2(G113gat), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n891), .A2(new_n719), .A3(new_n530), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n888), .A2(new_n890), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n715), .A2(new_n763), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n894), .A2(new_n743), .A3(new_n670), .A4(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(G113gat), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n896), .B2(G113gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n893), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n900), .B(new_n901), .ZN(G1340gat));
  INV_X1    g701(.A(new_n743), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(new_n888), .B2(new_n890), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n895), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(new_n316), .A3(new_n613), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n530), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n763), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n612), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n906), .B1(new_n909), .B2(new_n316), .ZN(G1341gat));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n309), .A3(new_n685), .ZN(new_n911));
  OAI21_X1  g710(.A(G127gat), .B1(new_n905), .B2(new_n754), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1342gat));
  NAND3_X1  g712(.A1(new_n711), .A2(new_n307), .A3(new_n719), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT56), .ZN(new_n916));
  OAI21_X1  g715(.A(G134gat), .B1(new_n905), .B2(new_n750), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(KEYINPUT56), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G1343gat));
  AOI21_X1  g718(.A(new_n451), .B1(new_n888), .B2(new_n890), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n714), .A2(new_n719), .ZN(new_n923));
  OR3_X1    g722(.A1(new_n733), .A2(KEYINPUT117), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT117), .B1(new_n733), .B2(new_n923), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n874), .A2(new_n875), .A3(new_n606), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n882), .B1(new_n788), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n750), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n685), .B1(new_n929), .B2(new_n886), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n742), .B1(new_n930), .B2(new_n889), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT57), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n922), .A2(new_n926), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G141gat), .B1(new_n933), .B2(new_n788), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n891), .A2(new_n742), .A3(new_n734), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n763), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n329), .A3(new_n670), .ZN(new_n937));
  XNOR2_X1  g736(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n934), .B2(new_n937), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(G1344gat));
  NAND3_X1  g740(.A1(new_n936), .A2(new_n331), .A3(new_n612), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n922), .A2(new_n932), .A3(new_n612), .A4(new_n926), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n331), .A2(KEYINPUT59), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n943), .A2(KEYINPUT119), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT119), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n920), .A2(new_n921), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n885), .A2(new_n606), .A3(new_n874), .A4(new_n875), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n685), .B1(new_n929), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n921), .B(new_n742), .C1(new_n951), .C2(new_n889), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n949), .A2(new_n612), .A3(new_n926), .A4(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n948), .B1(new_n953), .B2(G148gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n942), .B1(new_n947), .B2(new_n954), .ZN(G1345gat));
  NOR3_X1   g754(.A1(new_n933), .A2(new_n335), .A3(new_n754), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n935), .A2(new_n763), .A3(new_n686), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n957), .A2(KEYINPUT120), .ZN(new_n958));
  AOI21_X1  g757(.A(G155gat), .B1(new_n957), .B2(KEYINPUT120), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1346gat));
  OAI21_X1  g759(.A(G162gat), .B1(new_n933), .B2(new_n750), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n711), .A2(new_n336), .A3(new_n719), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n935), .B2(new_n962), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n714), .A2(new_n719), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n894), .A2(new_n743), .A3(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n904), .A2(KEYINPUT123), .A3(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n969), .A2(new_n209), .A3(new_n788), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n714), .B1(new_n888), .B2(new_n890), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n530), .A2(new_n763), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT121), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n974), .A2(KEYINPUT122), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(KEYINPUT122), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(new_n670), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n970), .B1(new_n209), .B2(new_n977), .ZN(G1348gat));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n612), .A3(new_n976), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n210), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n612), .A2(G176gat), .ZN(new_n981));
  OR3_X1    g780(.A1(new_n969), .A2(KEYINPUT124), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(KEYINPUT124), .B1(new_n969), .B2(new_n981), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(G1349gat));
  NAND4_X1  g783(.A1(new_n971), .A2(new_n225), .A3(new_n685), .A4(new_n973), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n967), .A2(new_n755), .A3(new_n968), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(new_n218), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT60), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  OAI221_X1 g790(.A(new_n985), .B1(new_n988), .B2(new_n989), .C1(new_n986), .C2(new_n218), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1350gat));
  NAND4_X1  g792(.A1(new_n975), .A2(new_n222), .A3(new_n711), .A4(new_n976), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n967), .A2(new_n711), .A3(new_n968), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n995), .A2(new_n996), .A3(G190gat), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n996), .B1(new_n995), .B2(G190gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(G1351gat));
  AND2_X1   g798(.A1(new_n949), .A2(new_n952), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n733), .A2(new_n714), .A3(new_n719), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n1000), .A2(new_n1001), .A3(new_n670), .A4(new_n1002), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n949), .A2(new_n952), .A3(new_n1002), .ZN(new_n1004));
  OAI21_X1  g803(.A(KEYINPUT127), .B1(new_n1004), .B2(new_n788), .ZN(new_n1005));
  XNOR2_X1  g804(.A(KEYINPUT126), .B(G197gat), .ZN(new_n1006));
  INV_X1    g805(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n733), .A2(new_n451), .A3(new_n719), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n971), .A2(new_n670), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1008), .A2(new_n1010), .ZN(G1352gat));
  OAI21_X1  g810(.A(G204gat), .B1(new_n1004), .B2(new_n613), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n971), .A2(new_n1009), .ZN(new_n1013));
  OR2_X1    g812(.A1(new_n613), .A2(G204gat), .ZN(new_n1014));
  OAI21_X1  g813(.A(KEYINPUT62), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OR3_X1    g814(.A1(new_n1013), .A2(KEYINPUT62), .A3(new_n1014), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(G1353gat));
  OR3_X1    g816(.A1(new_n1013), .A2(G211gat), .A3(new_n686), .ZN(new_n1018));
  NAND4_X1  g817(.A1(new_n949), .A2(new_n685), .A3(new_n952), .A4(new_n1002), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1019), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1020));
  INV_X1    g819(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g820(.A(KEYINPUT63), .B1(new_n1019), .B2(G211gat), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(G1354gat));
  OAI21_X1  g822(.A(G218gat), .B1(new_n1004), .B2(new_n750), .ZN(new_n1024));
  OR2_X1    g823(.A1(new_n750), .A2(G218gat), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1024), .B1(new_n1013), .B2(new_n1025), .ZN(G1355gat));
endmodule


