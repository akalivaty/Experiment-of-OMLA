

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803;

  OR2_X1 U363 ( .A1(n703), .A2(G902), .ZN(n503) );
  BUF_X1 U364 ( .A(G146), .Z(n341) );
  XNOR2_X2 U365 ( .A(n546), .B(n495), .ZN(n795) );
  AND2_X1 U366 ( .A1(n695), .A2(n694), .ZN(n461) );
  INV_X1 U367 ( .A(n341), .ZN(n530) );
  INV_X1 U368 ( .A(G953), .ZN(n796) );
  XNOR2_X1 U369 ( .A(n584), .B(KEYINPUT32), .ZN(n694) );
  BUF_X1 U370 ( .A(G128), .Z(n368) );
  AND2_X1 U371 ( .A1(n375), .A2(n374), .ZN(n342) );
  XNOR2_X2 U372 ( .A(n463), .B(n464), .ZN(n460) );
  NOR2_X2 U373 ( .A1(n684), .A2(n677), .ZN(n463) );
  INV_X2 U374 ( .A(n701), .ZN(n466) );
  AND2_X1 U375 ( .A1(n353), .A2(n351), .ZN(n343) );
  AND2_X2 U376 ( .A1(n473), .A2(n472), .ZN(n471) );
  NOR2_X2 U377 ( .A1(n589), .A2(n556), .ZN(n558) );
  XNOR2_X2 U378 ( .A(n565), .B(n564), .ZN(n355) );
  XNOR2_X2 U379 ( .A(n428), .B(n485), .ZN(n505) );
  XNOR2_X1 U380 ( .A(n505), .B(n348), .ZN(n781) );
  AND2_X1 U381 ( .A1(n370), .A2(n655), .ZN(n722) );
  NAND2_X1 U382 ( .A1(n482), .A2(n433), .ZN(n346) );
  OR2_X1 U383 ( .A1(n658), .A2(n413), .ZN(n668) );
  INV_X1 U384 ( .A(n401), .ZN(n400) );
  OR2_X1 U385 ( .A1(n637), .A2(n636), .ZN(n401) );
  INV_X1 U386 ( .A(n754), .ZN(n399) );
  INV_X1 U387 ( .A(n402), .ZN(n725) );
  INV_X1 U388 ( .A(n405), .ZN(n662) );
  XNOR2_X1 U389 ( .A(n622), .B(n621), .ZN(n482) );
  NAND2_X1 U390 ( .A1(n619), .A2(n618), .ZN(n402) );
  OR2_X1 U391 ( .A1(n411), .A2(n636), .ZN(n622) );
  OR2_X1 U392 ( .A1(n411), .A2(n566), .ZN(n352) );
  XNOR2_X1 U393 ( .A(n607), .B(n369), .ZN(n411) );
  NAND2_X1 U394 ( .A1(n636), .A2(n490), .ZN(n489) );
  AND2_X1 U395 ( .A1(n691), .A2(G953), .ZN(n780) );
  XNOR2_X1 U396 ( .A(G113), .B(KEYINPUT71), .ZN(n499) );
  NAND2_X1 U397 ( .A1(G902), .A2(G469), .ZN(n382) );
  BUF_X1 U398 ( .A(G104), .Z(n475) );
  INV_X1 U399 ( .A(KEYINPUT19), .ZN(n453) );
  INV_X1 U400 ( .A(G469), .ZN(n380) );
  INV_X1 U401 ( .A(G902), .ZN(n379) );
  AND2_X1 U402 ( .A1(n443), .A2(n441), .ZN(n440) );
  AND2_X1 U403 ( .A1(n450), .A2(n448), .ZN(n447) );
  AND2_X1 U404 ( .A1(n367), .A2(n604), .ZN(n473) );
  OR2_X1 U405 ( .A1(n714), .A2(n728), .ZN(n620) );
  NAND2_X1 U406 ( .A1(n350), .A2(KEYINPUT66), .ZN(n349) );
  BUF_X1 U407 ( .A(n598), .Z(n803) );
  AND2_X1 U408 ( .A1(n407), .A2(n410), .ZN(n674) );
  NOR2_X1 U409 ( .A1(n750), .A2(n613), .ZN(n590) );
  OR2_X1 U410 ( .A1(n613), .A2(n605), .ZN(n606) );
  NOR2_X1 U411 ( .A1(n480), .A2(n667), .ZN(n409) );
  NOR2_X1 U412 ( .A1(n457), .A2(KEYINPUT48), .ZN(n479) );
  XNOR2_X1 U413 ( .A(n396), .B(n648), .ZN(n480) );
  XNOR2_X1 U414 ( .A(n426), .B(G131), .ZN(G33) );
  NAND2_X1 U415 ( .A1(n358), .A2(n356), .ZN(n589) );
  AND2_X1 U416 ( .A1(n723), .A2(n652), .ZN(n653) );
  AND2_X1 U417 ( .A1(n361), .A2(n359), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n397), .B(n412), .ZN(n426) );
  XNOR2_X1 U419 ( .A(n418), .B(n417), .ZN(n416) );
  NAND2_X1 U420 ( .A1(n634), .A2(n725), .ZN(n397) );
  XNOR2_X1 U421 ( .A(n646), .B(n645), .ZN(n427) );
  NAND2_X1 U422 ( .A1(n388), .A2(n387), .ZN(n750) );
  NAND2_X1 U423 ( .A1(n357), .A2(n342), .ZN(n356) );
  XNOR2_X1 U424 ( .A(n651), .B(n650), .ZN(n723) );
  XNOR2_X1 U425 ( .A(n371), .B(n654), .ZN(n370) );
  AND2_X1 U426 ( .A1(n376), .A2(n452), .ZN(n357) );
  NOR2_X1 U427 ( .A1(n669), .A2(n405), .ZN(n418) );
  AND2_X1 U428 ( .A1(n390), .A2(n389), .ZN(n388) );
  XNOR2_X1 U429 ( .A(n346), .B(n633), .ZN(n634) );
  NAND2_X1 U430 ( .A1(n406), .A2(n423), .ZN(n376) );
  NAND2_X1 U431 ( .A1(n400), .A2(n399), .ZN(n639) );
  NOR2_X1 U432 ( .A1(n755), .A2(n401), .ZN(n756) );
  NAND2_X1 U433 ( .A1(n423), .A2(n488), .ZN(n656) );
  AND2_X1 U434 ( .A1(n630), .A2(n487), .ZN(n372) );
  NAND2_X1 U435 ( .A1(n414), .A2(n751), .ZN(n413) );
  INV_X1 U436 ( .A(n366), .ZN(n403) );
  XNOR2_X1 U437 ( .A(n425), .B(KEYINPUT28), .ZN(n424) );
  INV_X1 U438 ( .A(n429), .ZN(n488) );
  OR2_X1 U439 ( .A1(n657), .A2(n402), .ZN(n658) );
  AND2_X1 U440 ( .A1(n421), .A2(n431), .ZN(n452) );
  BUF_X1 U441 ( .A(n738), .Z(n366) );
  INV_X1 U442 ( .A(n659), .ZN(n414) );
  OR2_X1 U443 ( .A1(n405), .A2(KEYINPUT109), .ZN(n395) );
  AND2_X1 U444 ( .A1(n352), .A2(n741), .ZN(n351) );
  NOR2_X1 U445 ( .A1(n411), .A2(n659), .ZN(n425) );
  NAND2_X1 U446 ( .A1(n429), .A2(KEYINPUT19), .ZN(n375) );
  NAND2_X1 U447 ( .A1(n487), .A2(n486), .ZN(n423) );
  XNOR2_X1 U448 ( .A(n588), .B(n587), .ZN(n738) );
  INV_X1 U449 ( .A(n741), .ZN(n404) );
  NAND2_X1 U450 ( .A1(n364), .A2(n489), .ZN(n429) );
  OR2_X2 U451 ( .A1(n381), .A2(n377), .ZN(n643) );
  XNOR2_X1 U452 ( .A(n616), .B(n615), .ZN(n619) );
  NAND2_X1 U453 ( .A1(n460), .A2(n490), .ZN(n364) );
  NAND2_X1 U454 ( .A1(n383), .A2(n382), .ZN(n381) );
  AND2_X1 U455 ( .A1(n489), .A2(n453), .ZN(n422) );
  XNOR2_X1 U456 ( .A(n538), .B(n537), .ZN(n616) );
  XNOR2_X1 U457 ( .A(n459), .B(n579), .ZN(n458) );
  NOR2_X1 U458 ( .A1(G902), .A2(n698), .ZN(n538) );
  NOR2_X1 U459 ( .A1(n709), .A2(G902), .ZN(n459) );
  NAND2_X1 U460 ( .A1(n419), .A2(G469), .ZN(n383) );
  XNOR2_X1 U461 ( .A(n555), .B(KEYINPUT21), .ZN(n740) );
  AND2_X1 U462 ( .A1(n486), .A2(KEYINPUT19), .ZN(n420) );
  INV_X1 U463 ( .A(n798), .ZN(n345) );
  XNOR2_X1 U464 ( .A(n781), .B(n511), .ZN(n347) );
  XNOR2_X1 U465 ( .A(n793), .B(n530), .ZN(n570) );
  XNOR2_X1 U466 ( .A(n559), .B(n504), .ZN(n348) );
  XNOR2_X1 U467 ( .A(n529), .B(KEYINPUT10), .ZN(n793) );
  OR2_X1 U468 ( .A1(n677), .A2(n552), .ZN(n554) );
  INV_X1 U469 ( .A(n435), .ZN(n391) );
  NAND2_X1 U470 ( .A1(n380), .A2(n379), .ZN(n378) );
  XNOR2_X1 U471 ( .A(n512), .B(KEYINPUT15), .ZN(n677) );
  INV_X1 U472 ( .A(n635), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n499), .B(KEYINPUT3), .ZN(n428) );
  XNOR2_X1 U474 ( .A(n670), .B(KEYINPUT112), .ZN(n417) );
  XNOR2_X1 U475 ( .A(G131), .B(G122), .ZN(n531) );
  XNOR2_X1 U476 ( .A(KEYINPUT16), .B(G122), .ZN(n504) );
  INV_X1 U477 ( .A(KEYINPUT107), .ZN(n369) );
  XNOR2_X1 U478 ( .A(KEYINPUT4), .B(G146), .ZN(n494) );
  XNOR2_X1 U479 ( .A(KEYINPUT18), .B(G125), .ZN(n507) );
  XNOR2_X1 U480 ( .A(G116), .B(G122), .ZN(n542) );
  XNOR2_X1 U481 ( .A(G134), .B(G107), .ZN(n539) );
  BUF_X1 U482 ( .A(KEYINPUT39), .Z(n633) );
  XNOR2_X1 U483 ( .A(G902), .B(KEYINPUT89), .ZN(n512) );
  XOR2_X1 U484 ( .A(KEYINPUT33), .B(KEYINPUT110), .Z(n435) );
  XNOR2_X2 U485 ( .A(n344), .B(n792), .ZN(n365) );
  XNOR2_X1 U486 ( .A(n347), .B(n344), .ZN(n684) );
  XNOR2_X2 U487 ( .A(n795), .B(G101), .ZN(n344) );
  XNOR2_X1 U488 ( .A(n674), .B(n345), .ZN(n797) );
  INV_X1 U489 ( .A(n634), .ZN(n672) );
  NAND2_X2 U490 ( .A1(n343), .A2(n349), .ZN(n695) );
  INV_X1 U491 ( .A(n355), .ZN(n350) );
  NAND2_X1 U492 ( .A1(n355), .A2(n354), .ZN(n353) );
  AND2_X1 U493 ( .A1(n411), .A2(n566), .ZN(n354) );
  NAND2_X1 U494 ( .A1(n360), .A2(n434), .ZN(n359) );
  NAND2_X1 U495 ( .A1(n452), .A2(n375), .ZN(n360) );
  NAND2_X1 U496 ( .A1(n362), .A2(n434), .ZN(n361) );
  INV_X1 U497 ( .A(n376), .ZN(n362) );
  INV_X1 U498 ( .A(n363), .ZN(n406) );
  NAND2_X1 U499 ( .A1(n364), .A2(n422), .ZN(n363) );
  XNOR2_X2 U500 ( .A(n365), .B(n563), .ZN(n419) );
  XNOR2_X1 U501 ( .A(n365), .B(n481), .ZN(n703) );
  AND2_X1 U502 ( .A1(n386), .A2(n394), .ZN(n385) );
  NAND2_X1 U503 ( .A1(n477), .A2(n391), .ZN(n384) );
  NAND2_X1 U504 ( .A1(n599), .A2(KEYINPUT44), .ZN(n367) );
  NAND2_X1 U505 ( .A1(n680), .A2(n676), .ZN(n678) );
  NAND2_X1 U506 ( .A1(n675), .A2(n674), .ZN(n680) );
  NOR2_X1 U507 ( .A1(n409), .A2(n408), .ZN(n407) );
  NAND2_X1 U508 ( .A1(n416), .A2(n631), .ZN(n733) );
  INV_X1 U509 ( .A(n607), .ZN(n611) );
  NAND2_X1 U510 ( .A1(n665), .A2(n666), .ZN(n457) );
  NAND2_X1 U511 ( .A1(n482), .A2(n372), .ZN(n371) );
  NAND2_X1 U512 ( .A1(n395), .A2(n373), .ZN(n392) );
  INV_X1 U513 ( .A(n657), .ZN(n373) );
  INV_X1 U514 ( .A(n434), .ZN(n374) );
  XNOR2_X2 U515 ( .A(n643), .B(KEYINPUT1), .ZN(n405) );
  NOR2_X1 U516 ( .A1(n419), .A2(n378), .ZN(n377) );
  NOR2_X1 U517 ( .A1(n384), .A2(n657), .ZN(n386) );
  NAND2_X1 U518 ( .A1(n394), .A2(n477), .ZN(n393) );
  NAND2_X1 U519 ( .A1(n385), .A2(n395), .ZN(n387) );
  NAND2_X1 U520 ( .A1(n393), .A2(n435), .ZN(n389) );
  NAND2_X1 U521 ( .A1(n392), .A2(n435), .ZN(n390) );
  NAND2_X1 U522 ( .A1(n476), .A2(n405), .ZN(n394) );
  NAND2_X1 U523 ( .A1(n398), .A2(n426), .ZN(n396) );
  INV_X1 U524 ( .A(n427), .ZN(n398) );
  AND2_X1 U525 ( .A1(n662), .A2(n404), .ZN(n602) );
  NOR2_X1 U526 ( .A1(n662), .A2(n403), .ZN(n612) );
  AND2_X1 U527 ( .A1(n662), .A2(n403), .ZN(n739) );
  NOR2_X1 U528 ( .A1(n662), .A2(n404), .ZN(n582) );
  NAND2_X1 U529 ( .A1(n478), .A2(n673), .ZN(n408) );
  NAND2_X1 U530 ( .A1(n479), .A2(n480), .ZN(n410) );
  NOR2_X1 U531 ( .A1(n658), .A2(n659), .ZN(n415) );
  NAND2_X1 U532 ( .A1(n415), .A2(n656), .ZN(n661) );
  XNOR2_X1 U533 ( .A(n419), .B(n772), .ZN(n773) );
  NAND2_X1 U534 ( .A1(n487), .A2(n420), .ZN(n421) );
  AND2_X1 U535 ( .A1(n643), .A2(n424), .ZN(n649) );
  XNOR2_X1 U536 ( .A(n427), .B(n693), .ZN(G39) );
  XNOR2_X2 U537 ( .A(n484), .B(n483), .ZN(n559) );
  INV_X1 U538 ( .A(KEYINPUT84), .ZN(n490) );
  XNOR2_X1 U539 ( .A(G119), .B(G116), .ZN(n485) );
  XNOR2_X1 U540 ( .A(G125), .B(G140), .ZN(n528) );
  NOR2_X1 U541 ( .A1(n442), .A2(n780), .ZN(n441) );
  NOR2_X1 U542 ( .A1(n455), .A2(G210), .ZN(n442) );
  NAND2_X1 U543 ( .A1(n446), .A2(n690), .ZN(n439) );
  XOR2_X1 U544 ( .A(n475), .B(KEYINPUT100), .Z(n523) );
  XNOR2_X1 U545 ( .A(KEYINPUT91), .B(KEYINPUT17), .ZN(n506) );
  INV_X1 U546 ( .A(G234), .ZN(n552) );
  NOR2_X1 U547 ( .A1(n636), .A2(n490), .ZN(n486) );
  INV_X1 U548 ( .A(n502), .ZN(n481) );
  NAND2_X1 U549 ( .A1(n620), .A2(n652), .ZN(n472) );
  XNOR2_X1 U550 ( .A(n368), .B(G119), .ZN(n571) );
  INV_X1 U551 ( .A(G143), .ZN(n492) );
  INV_X1 U552 ( .A(n458), .ZN(n741) );
  NOR2_X1 U553 ( .A1(n449), .A2(n780), .ZN(n448) );
  NOR2_X1 U554 ( .A1(n456), .A2(G475), .ZN(n449) );
  NAND2_X1 U555 ( .A1(n446), .A2(n699), .ZN(n445) );
  INV_X1 U556 ( .A(KEYINPUT56), .ZN(n454) );
  XOR2_X1 U557 ( .A(n467), .B(KEYINPUT45), .Z(n430) );
  OR2_X1 U558 ( .A1(n623), .A2(n520), .ZN(n431) );
  XOR2_X1 U559 ( .A(n656), .B(KEYINPUT19), .Z(n432) );
  AND2_X1 U560 ( .A1(n630), .A2(n752), .ZN(n433) );
  XNOR2_X1 U561 ( .A(KEYINPUT88), .B(KEYINPUT0), .ZN(n434) );
  INV_X1 U562 ( .A(n690), .ZN(n455) );
  XNOR2_X1 U563 ( .A(n689), .B(n688), .ZN(n690) );
  INV_X1 U564 ( .A(n699), .ZN(n456) );
  XNOR2_X1 U565 ( .A(n698), .B(n697), .ZN(n699) );
  AND2_X1 U566 ( .A1(n456), .A2(G475), .ZN(n436) );
  AND2_X1 U567 ( .A1(n455), .A2(G210), .ZN(n437) );
  XNOR2_X1 U568 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n438) );
  NAND2_X1 U569 ( .A1(n440), .A2(n439), .ZN(n444) );
  NAND2_X1 U570 ( .A1(n466), .A2(n437), .ZN(n443) );
  XNOR2_X1 U571 ( .A(n444), .B(n454), .ZN(G51) );
  NAND2_X1 U572 ( .A1(n447), .A2(n445), .ZN(n451) );
  INV_X1 U573 ( .A(n466), .ZN(n446) );
  NAND2_X1 U574 ( .A1(n466), .A2(n436), .ZN(n450) );
  XNOR2_X1 U575 ( .A(n451), .B(n438), .ZN(G60) );
  NAND2_X1 U576 ( .A1(n457), .A2(KEYINPUT48), .ZN(n478) );
  BUF_X1 U577 ( .A(n589), .Z(n613) );
  AND2_X1 U578 ( .A1(n738), .A2(KEYINPUT109), .ZN(n476) );
  OR2_X1 U579 ( .A1(n738), .A2(KEYINPUT109), .ZN(n477) );
  NAND2_X1 U580 ( .A1(n695), .A2(n694), .ZN(n462) );
  XOR2_X1 U581 ( .A(n514), .B(KEYINPUT92), .Z(n464) );
  BUF_X1 U582 ( .A(n474), .Z(n465) );
  NAND2_X1 U583 ( .A1(n465), .A2(n471), .ZN(n467) );
  NAND2_X1 U584 ( .A1(n474), .A2(n471), .ZN(n470) );
  XNOR2_X1 U585 ( .A(n470), .B(KEYINPUT45), .ZN(n675) );
  NAND2_X1 U586 ( .A1(n462), .A2(n491), .ZN(n468) );
  NAND2_X1 U587 ( .A1(n469), .A2(n468), .ZN(n474) );
  NAND2_X1 U588 ( .A1(n461), .A2(n595), .ZN(n469) );
  XNOR2_X2 U589 ( .A(G110), .B(KEYINPUT90), .ZN(n483) );
  XNOR2_X2 U590 ( .A(G107), .B(G104), .ZN(n484) );
  INV_X1 U591 ( .A(n460), .ZN(n487) );
  AND2_X1 U592 ( .A1(n597), .A2(n596), .ZN(n491) );
  AND2_X1 U593 ( .A1(n643), .A2(n641), .ZN(n628) );
  INV_X1 U594 ( .A(KEYINPUT66), .ZN(n566) );
  XNOR2_X1 U595 ( .A(n776), .B(KEYINPUT126), .ZN(n777) );
  XNOR2_X1 U596 ( .A(n778), .B(n777), .ZN(n779) );
  XNOR2_X2 U597 ( .A(KEYINPUT79), .B(G128), .ZN(n493) );
  XNOR2_X2 U598 ( .A(n493), .B(n492), .ZN(n546) );
  XNOR2_X1 U599 ( .A(n494), .B(KEYINPUT69), .ZN(n495) );
  INV_X1 U600 ( .A(KEYINPUT70), .ZN(n496) );
  XNOR2_X1 U601 ( .A(n496), .B(G131), .ZN(n498) );
  XNOR2_X1 U602 ( .A(G137), .B(G134), .ZN(n497) );
  XNOR2_X1 U603 ( .A(n498), .B(n497), .ZN(n792) );
  NOR2_X1 U604 ( .A1(G953), .A2(G237), .ZN(n521) );
  NAND2_X1 U605 ( .A1(n521), .A2(G210), .ZN(n500) );
  XNOR2_X1 U606 ( .A(n500), .B(KEYINPUT5), .ZN(n501) );
  XNOR2_X1 U607 ( .A(n505), .B(n501), .ZN(n502) );
  INV_X1 U608 ( .A(G472), .ZN(n700) );
  XNOR2_X2 U609 ( .A(n503), .B(n700), .ZN(n607) );
  XNOR2_X1 U610 ( .A(n507), .B(n506), .ZN(n510) );
  NAND2_X1 U611 ( .A1(n796), .A2(G224), .ZN(n508) );
  XNOR2_X1 U612 ( .A(n508), .B(KEYINPUT77), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U614 ( .A(G237), .ZN(n513) );
  NAND2_X1 U615 ( .A1(n379), .A2(n513), .ZN(n515) );
  NAND2_X1 U616 ( .A1(n515), .A2(G210), .ZN(n514) );
  NAND2_X1 U617 ( .A1(n515), .A2(G214), .ZN(n751) );
  INV_X1 U618 ( .A(n751), .ZN(n636) );
  NAND2_X1 U619 ( .A1(G234), .A2(G237), .ZN(n516) );
  XNOR2_X1 U620 ( .A(n516), .B(KEYINPUT14), .ZN(n517) );
  XNOR2_X1 U621 ( .A(KEYINPUT74), .B(n517), .ZN(n519) );
  NAND2_X1 U622 ( .A1(n519), .A2(G952), .ZN(n518) );
  XNOR2_X1 U623 ( .A(n518), .B(KEYINPUT93), .ZN(n763) );
  AND2_X1 U624 ( .A1(n763), .A2(n796), .ZN(n623) );
  NAND2_X1 U625 ( .A1(G902), .A2(n519), .ZN(n624) );
  XOR2_X1 U626 ( .A(G898), .B(KEYINPUT94), .Z(n787) );
  NAND2_X1 U627 ( .A1(G953), .A2(n787), .ZN(n783) );
  NOR2_X1 U628 ( .A1(n624), .A2(n783), .ZN(n520) );
  NAND2_X1 U629 ( .A1(G214), .A2(n521), .ZN(n522) );
  XNOR2_X1 U630 ( .A(n523), .B(n522), .ZN(n527) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n525) );
  XNOR2_X1 U632 ( .A(G113), .B(KEYINPUT99), .ZN(n524) );
  XNOR2_X1 U633 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U634 ( .A(n527), .B(n526), .Z(n536) );
  INV_X1 U635 ( .A(n528), .ZN(n529) );
  XOR2_X1 U636 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n533) );
  XOR2_X1 U637 ( .A(n531), .B(G143), .Z(n532) );
  XNOR2_X1 U638 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U639 ( .A(n570), .B(n534), .ZN(n535) );
  XNOR2_X1 U640 ( .A(n536), .B(n535), .ZN(n698) );
  XNOR2_X1 U641 ( .A(KEYINPUT13), .B(G475), .ZN(n537) );
  XOR2_X1 U642 ( .A(KEYINPUT7), .B(KEYINPUT104), .Z(n540) );
  XNOR2_X1 U643 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U644 ( .A(n541), .B(KEYINPUT9), .Z(n543) );
  XNOR2_X1 U645 ( .A(n543), .B(n542), .ZN(n548) );
  AND2_X1 U646 ( .A1(G234), .A2(n796), .ZN(n544) );
  XNOR2_X1 U647 ( .A(KEYINPUT8), .B(n544), .ZN(n572) );
  NAND2_X1 U648 ( .A1(n572), .A2(G217), .ZN(n545) );
  XNOR2_X1 U649 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U650 ( .A(n548), .B(n547), .ZN(n776) );
  OR2_X1 U651 ( .A1(n776), .A2(G902), .ZN(n549) );
  XNOR2_X1 U652 ( .A(n549), .B(G478), .ZN(n617) );
  NOR2_X1 U653 ( .A1(n616), .A2(n617), .ZN(n551) );
  INV_X1 U654 ( .A(KEYINPUT106), .ZN(n550) );
  XNOR2_X1 U655 ( .A(n551), .B(n550), .ZN(n754) );
  XOR2_X1 U656 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n553) );
  XNOR2_X1 U657 ( .A(n554), .B(n553), .ZN(n577) );
  NAND2_X1 U658 ( .A1(n577), .A2(G221), .ZN(n555) );
  XNOR2_X1 U659 ( .A(n740), .B(KEYINPUT96), .ZN(n585) );
  OR2_X1 U660 ( .A1(n754), .A2(n585), .ZN(n556) );
  XOR2_X1 U661 ( .A(KEYINPUT73), .B(KEYINPUT22), .Z(n557) );
  XNOR2_X1 U662 ( .A(n558), .B(n557), .ZN(n580) );
  XOR2_X1 U663 ( .A(G140), .B(KEYINPUT76), .Z(n561) );
  NAND2_X1 U664 ( .A1(G227), .A2(n796), .ZN(n560) );
  XNOR2_X1 U665 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U666 ( .A(n559), .B(n562), .ZN(n563) );
  NAND2_X1 U667 ( .A1(n580), .A2(n662), .ZN(n565) );
  INV_X1 U668 ( .A(KEYINPUT108), .ZN(n564) );
  XNOR2_X1 U669 ( .A(G110), .B(G137), .ZN(n568) );
  XNOR2_X1 U670 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n567) );
  XNOR2_X1 U671 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U672 ( .A(n570), .B(n569), .ZN(n576) );
  XNOR2_X1 U673 ( .A(n571), .B(KEYINPUT72), .ZN(n574) );
  NAND2_X1 U674 ( .A1(n572), .A2(G221), .ZN(n573) );
  XNOR2_X1 U675 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U676 ( .A(n576), .B(n575), .ZN(n709) );
  NAND2_X1 U677 ( .A1(n577), .A2(G217), .ZN(n578) );
  XNOR2_X1 U678 ( .A(n578), .B(KEYINPUT25), .ZN(n579) );
  XNOR2_X1 U679 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n581) );
  XNOR2_X1 U680 ( .A(n607), .B(n581), .ZN(n657) );
  NAND2_X1 U681 ( .A1(n580), .A2(n657), .ZN(n601) );
  INV_X1 U682 ( .A(n601), .ZN(n583) );
  NAND2_X1 U683 ( .A1(n583), .A2(n582), .ZN(n584) );
  INV_X1 U684 ( .A(n585), .ZN(n586) );
  NAND2_X1 U685 ( .A1(n586), .A2(n458), .ZN(n588) );
  INV_X1 U686 ( .A(KEYINPUT68), .ZN(n587) );
  XNOR2_X1 U687 ( .A(n590), .B(KEYINPUT34), .ZN(n591) );
  AND2_X1 U688 ( .A1(n616), .A2(n617), .ZN(n655) );
  NAND2_X1 U689 ( .A1(n591), .A2(n655), .ZN(n593) );
  INV_X1 U690 ( .A(KEYINPUT35), .ZN(n592) );
  XNOR2_X2 U691 ( .A(n593), .B(n592), .ZN(n598) );
  NOR2_X1 U692 ( .A1(KEYINPUT44), .A2(KEYINPUT83), .ZN(n594) );
  NAND2_X1 U693 ( .A1(n803), .A2(n594), .ZN(n595) );
  NAND2_X1 U694 ( .A1(n598), .A2(KEYINPUT83), .ZN(n597) );
  INV_X1 U695 ( .A(KEYINPUT44), .ZN(n596) );
  INV_X1 U696 ( .A(n598), .ZN(n599) );
  INV_X1 U697 ( .A(KEYINPUT82), .ZN(n600) );
  XNOR2_X1 U698 ( .A(n601), .B(n600), .ZN(n603) );
  AND2_X1 U699 ( .A1(n603), .A2(n602), .ZN(n712) );
  INV_X1 U700 ( .A(n712), .ZN(n604) );
  NAND2_X1 U701 ( .A1(n643), .A2(n366), .ZN(n605) );
  XNOR2_X1 U702 ( .A(n606), .B(KEYINPUT97), .ZN(n608) );
  NAND2_X1 U703 ( .A1(n608), .A2(n607), .ZN(n610) );
  INV_X1 U704 ( .A(KEYINPUT98), .ZN(n609) );
  XNOR2_X1 U705 ( .A(n610), .B(n609), .ZN(n714) );
  NAND2_X1 U706 ( .A1(n612), .A2(n611), .ZN(n746) );
  OR2_X1 U707 ( .A1(n613), .A2(n746), .ZN(n614) );
  XNOR2_X1 U708 ( .A(n614), .B(KEYINPUT31), .ZN(n728) );
  INV_X1 U709 ( .A(KEYINPUT103), .ZN(n615) );
  INV_X1 U710 ( .A(n617), .ZN(n618) );
  NOR2_X1 U711 ( .A1(n619), .A2(n618), .ZN(n727) );
  NOR2_X1 U712 ( .A1(n727), .A2(n725), .ZN(n755) );
  INV_X1 U713 ( .A(n755), .ZN(n652) );
  XNOR2_X1 U714 ( .A(KEYINPUT113), .B(KEYINPUT30), .ZN(n621) );
  INV_X1 U715 ( .A(n623), .ZN(n627) );
  NOR2_X1 U716 ( .A1(G900), .A2(n624), .ZN(n625) );
  NAND2_X1 U717 ( .A1(n625), .A2(G953), .ZN(n626) );
  NAND2_X1 U718 ( .A1(n627), .A2(n626), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n738), .A2(n628), .ZN(n629) );
  XNOR2_X1 U720 ( .A(n629), .B(KEYINPUT75), .ZN(n630) );
  BUF_X1 U721 ( .A(n460), .Z(n631) );
  INV_X1 U722 ( .A(KEYINPUT38), .ZN(n632) );
  XNOR2_X1 U723 ( .A(n631), .B(n632), .ZN(n637) );
  INV_X1 U724 ( .A(n637), .ZN(n752) );
  XNOR2_X1 U725 ( .A(KEYINPUT115), .B(KEYINPUT40), .ZN(n635) );
  INV_X1 U726 ( .A(KEYINPUT41), .ZN(n638) );
  XNOR2_X1 U727 ( .A(n639), .B(n638), .ZN(n765) );
  INV_X1 U728 ( .A(n740), .ZN(n640) );
  AND2_X1 U729 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U730 ( .A1(n642), .A2(n741), .ZN(n659) );
  INV_X1 U731 ( .A(n649), .ZN(n644) );
  OR2_X1 U732 ( .A1(n765), .A2(n644), .ZN(n646) );
  INV_X1 U733 ( .A(KEYINPUT42), .ZN(n645) );
  XNOR2_X1 U734 ( .A(KEYINPUT81), .B(KEYINPUT46), .ZN(n647) );
  XNOR2_X1 U735 ( .A(n647), .B(KEYINPUT64), .ZN(n648) );
  NAND2_X1 U736 ( .A1(n649), .A2(n432), .ZN(n651) );
  INV_X1 U737 ( .A(KEYINPUT78), .ZN(n650) );
  XNOR2_X1 U738 ( .A(n653), .B(KEYINPUT47), .ZN(n666) );
  INV_X1 U739 ( .A(KEYINPUT114), .ZN(n654) );
  XNOR2_X1 U740 ( .A(KEYINPUT116), .B(KEYINPUT36), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n661), .B(n660), .ZN(n663) );
  OR2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n730) );
  INV_X1 U743 ( .A(n730), .ZN(n664) );
  NOR2_X1 U744 ( .A1(n722), .A2(n664), .ZN(n665) );
  INV_X1 U745 ( .A(KEYINPUT48), .ZN(n667) );
  XOR2_X1 U746 ( .A(KEYINPUT111), .B(n668), .Z(n669) );
  INV_X1 U747 ( .A(KEYINPUT43), .ZN(n670) );
  INV_X1 U748 ( .A(n727), .ZN(n671) );
  OR2_X1 U749 ( .A1(n672), .A2(n671), .ZN(n692) );
  AND2_X1 U750 ( .A1(n733), .A2(n692), .ZN(n673) );
  INV_X1 U751 ( .A(KEYINPUT2), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n679), .B(KEYINPUT65), .ZN(n683) );
  BUF_X1 U754 ( .A(n680), .Z(n735) );
  INV_X1 U755 ( .A(n735), .ZN(n681) );
  NAND2_X1 U756 ( .A1(n681), .A2(KEYINPUT2), .ZN(n682) );
  NAND2_X1 U757 ( .A1(n683), .A2(n682), .ZN(n701) );
  BUF_X1 U758 ( .A(n684), .Z(n689) );
  XNOR2_X1 U759 ( .A(KEYINPUT86), .B(KEYINPUT55), .ZN(n685) );
  XNOR2_X1 U760 ( .A(n685), .B(KEYINPUT87), .ZN(n687) );
  XOR2_X1 U761 ( .A(KEYINPUT124), .B(KEYINPUT54), .Z(n686) );
  XOR2_X1 U762 ( .A(n687), .B(n686), .Z(n688) );
  INV_X1 U763 ( .A(G952), .ZN(n691) );
  XNOR2_X1 U764 ( .A(n692), .B(G134), .ZN(G36) );
  XNOR2_X1 U765 ( .A(G137), .B(KEYINPUT127), .ZN(n693) );
  XNOR2_X1 U766 ( .A(n694), .B(G119), .ZN(G21) );
  XOR2_X1 U767 ( .A(G110), .B(KEYINPUT119), .Z(n696) );
  XNOR2_X1 U768 ( .A(n695), .B(n696), .ZN(G12) );
  XNOR2_X1 U769 ( .A(KEYINPUT125), .B(KEYINPUT59), .ZN(n697) );
  NOR2_X1 U770 ( .A1(n701), .A2(n700), .ZN(n705) );
  XNOR2_X1 U771 ( .A(KEYINPUT117), .B(KEYINPUT62), .ZN(n702) );
  XNOR2_X1 U772 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U773 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U774 ( .A1(n706), .A2(n780), .ZN(n708) );
  XNOR2_X1 U775 ( .A(KEYINPUT85), .B(KEYINPUT63), .ZN(n707) );
  XNOR2_X1 U776 ( .A(n708), .B(n707), .ZN(G57) );
  NAND2_X1 U777 ( .A1(n466), .A2(G217), .ZN(n710) );
  XNOR2_X1 U778 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U779 ( .A1(n711), .A2(n780), .ZN(G66) );
  XOR2_X1 U780 ( .A(G101), .B(n712), .Z(G3) );
  NAND2_X1 U781 ( .A1(n714), .A2(n725), .ZN(n713) );
  XNOR2_X1 U782 ( .A(n713), .B(n475), .ZN(G6) );
  XNOR2_X1 U783 ( .A(G107), .B(KEYINPUT118), .ZN(n718) );
  XOR2_X1 U784 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n716) );
  NAND2_X1 U785 ( .A1(n727), .A2(n714), .ZN(n715) );
  XNOR2_X1 U786 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U787 ( .A(n718), .B(n717), .ZN(G9) );
  XOR2_X1 U788 ( .A(KEYINPUT120), .B(KEYINPUT29), .Z(n720) );
  NAND2_X1 U789 ( .A1(n727), .A2(n723), .ZN(n719) );
  XNOR2_X1 U790 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U791 ( .A(n368), .B(n721), .ZN(G30) );
  XOR2_X1 U792 ( .A(G143), .B(n722), .Z(G45) );
  NAND2_X1 U793 ( .A1(n723), .A2(n725), .ZN(n724) );
  XNOR2_X1 U794 ( .A(n724), .B(n341), .ZN(G48) );
  NAND2_X1 U795 ( .A1(n728), .A2(n725), .ZN(n726) );
  XNOR2_X1 U796 ( .A(n726), .B(G113), .ZN(G15) );
  NAND2_X1 U797 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U798 ( .A(n729), .B(G116), .ZN(G18) );
  XNOR2_X1 U799 ( .A(KEYINPUT121), .B(KEYINPUT37), .ZN(n731) );
  XNOR2_X1 U800 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U801 ( .A(G125), .B(n732), .ZN(G27) );
  XNOR2_X1 U802 ( .A(n733), .B(G140), .ZN(n734) );
  XNOR2_X1 U803 ( .A(KEYINPUT122), .B(n734), .ZN(G42) );
  NAND2_X1 U804 ( .A1(n735), .A2(KEYINPUT80), .ZN(n736) );
  XNOR2_X1 U805 ( .A(n736), .B(KEYINPUT2), .ZN(n737) );
  NAND2_X1 U806 ( .A1(n737), .A2(n796), .ZN(n770) );
  XOR2_X1 U807 ( .A(KEYINPUT50), .B(n739), .Z(n745) );
  NAND2_X1 U808 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U809 ( .A(n742), .B(KEYINPUT49), .ZN(n743) );
  NOR2_X1 U810 ( .A1(n611), .A2(n743), .ZN(n744) );
  NAND2_X1 U811 ( .A1(n745), .A2(n744), .ZN(n747) );
  AND2_X1 U812 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U813 ( .A(KEYINPUT51), .B(n748), .Z(n749) );
  NOR2_X1 U814 ( .A1(n765), .A2(n749), .ZN(n760) );
  BUF_X1 U815 ( .A(n750), .Z(n764) );
  NOR2_X1 U816 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U817 ( .A1(n754), .A2(n753), .ZN(n757) );
  NOR2_X1 U818 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U819 ( .A1(n764), .A2(n758), .ZN(n759) );
  NOR2_X1 U820 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U821 ( .A(KEYINPUT52), .B(n761), .Z(n762) );
  NAND2_X1 U822 ( .A1(n763), .A2(n762), .ZN(n767) );
  OR2_X1 U823 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U824 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U825 ( .A(KEYINPUT123), .B(n768), .Z(n769) );
  NOR2_X1 U826 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U827 ( .A(KEYINPUT53), .B(n771), .ZN(G75) );
  NAND2_X1 U828 ( .A1(n466), .A2(G469), .ZN(n774) );
  XOR2_X1 U829 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n772) );
  XNOR2_X1 U830 ( .A(n774), .B(n773), .ZN(n775) );
  NOR2_X1 U831 ( .A1(n780), .A2(n775), .ZN(G54) );
  NAND2_X1 U832 ( .A1(n466), .A2(G478), .ZN(n778) );
  NOR2_X1 U833 ( .A1(n780), .A2(n779), .ZN(G63) );
  BUF_X1 U834 ( .A(n781), .Z(n782) );
  XNOR2_X1 U835 ( .A(n782), .B(G101), .ZN(n784) );
  NAND2_X1 U836 ( .A1(n784), .A2(n783), .ZN(n791) );
  NOR2_X1 U837 ( .A1(n430), .A2(G953), .ZN(n789) );
  NAND2_X1 U838 ( .A1(G953), .A2(G224), .ZN(n785) );
  XOR2_X1 U839 ( .A(KEYINPUT61), .B(n785), .Z(n786) );
  NOR2_X1 U840 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U841 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U842 ( .A(n791), .B(n790), .ZN(G69) );
  XNOR2_X1 U843 ( .A(n793), .B(n792), .ZN(n794) );
  XNOR2_X1 U844 ( .A(n795), .B(n794), .ZN(n798) );
  NAND2_X1 U845 ( .A1(n797), .A2(n796), .ZN(n802) );
  XNOR2_X1 U846 ( .A(G227), .B(n798), .ZN(n799) );
  NAND2_X1 U847 ( .A1(n799), .A2(G900), .ZN(n800) );
  NAND2_X1 U848 ( .A1(G953), .A2(n800), .ZN(n801) );
  NAND2_X1 U849 ( .A1(n802), .A2(n801), .ZN(G72) );
  XNOR2_X1 U850 ( .A(n803), .B(G122), .ZN(G24) );
endmodule

