//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT65), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(G101), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n462), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n474), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n475), .A2(new_n463), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n466), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT67), .Z(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  OAI211_X1 g057(.A(G2105), .B(new_n469), .C1(new_n462), .C2(new_n470), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n467), .A2(KEYINPUT65), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n468), .B1(new_n487), .B2(KEYINPUT3), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n463), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  OAI221_X1 g065(.A(new_n481), .B1(new_n482), .B2(new_n483), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND2_X1  g067(.A1(new_n463), .A2(G138), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n469), .B(new_n494), .C1(new_n462), .C2(new_n470), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(new_n474), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n504));
  INV_X1    g079(.A(G126), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT68), .B1(new_n483), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n488), .A2(new_n507), .A3(G126), .A4(G2105), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n502), .A2(new_n504), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(new_n515), .B1(new_n512), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(G651), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n519), .A2(new_n521), .B1(new_n518), .B2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n520), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n527), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT72), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT72), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n516), .A2(new_n522), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(G89), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n523), .A2(new_n543), .B1(new_n525), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n520), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(G171));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT73), .B(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n537), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n522), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n520), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n549), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n555), .A2(new_n520), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n558), .A2(KEYINPUT74), .A3(new_n553), .A4(new_n551), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  XNOR2_X1  g141(.A(new_n523), .B(KEYINPUT76), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G91), .ZN(new_n568));
  NOR2_X1   g143(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n569));
  AND2_X1   g144(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n552), .B(G53), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n552), .A2(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n569), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n520), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n568), .A2(new_n573), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  NAND2_X1  g152(.A1(new_n567), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n552), .A2(G49), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n516), .A2(G61), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n520), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n522), .A2(G48), .A3(G543), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n523), .B(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(G305));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n523), .A2(new_n592), .B1(new_n525), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n520), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n594), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT10), .B1(new_n589), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n516), .A2(G66), .ZN(new_n601));
  INV_X1    g176(.A(G79), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n514), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n552), .B2(G54), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n567), .A2(new_n605), .A3(G92), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n600), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n598), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n598), .B1(new_n608), .B2(G868), .ZN(G321));
  MUX2_X1   g185(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g186(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n608), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n608), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n472), .A2(G135), .ZN(new_n619));
  INV_X1    g194(.A(new_n483), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n619), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT78), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2096), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n474), .A2(new_n462), .A3(new_n463), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XOR2_X1   g203(.A(KEYINPUT13), .B(G2100), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT80), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2451), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2435), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2438), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n635), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT81), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n646), .A2(G14), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT82), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT17), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n650), .B2(new_n651), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n653), .B1(new_n652), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  AOI22_X1  g247(.A1(new_n670), .A2(new_n671), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  OR3_X1    g248(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n674), .C1(new_n671), .C2(new_n670), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G1981), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G229));
  NOR2_X1   g256(.A1(G29), .A2(G33), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT89), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT25), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n472), .A2(G139), .ZN(new_n686));
  AOI22_X1  g261(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(new_n463), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n682), .B1(new_n690), .B2(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G2072), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT91), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n620), .A2(G129), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n695));
  NAND3_X1  g270(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n462), .A2(G105), .A3(new_n463), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT93), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n702));
  INV_X1    g277(.A(G141), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n489), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n472), .A2(KEYINPUT92), .A3(G141), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G32), .B(new_n707), .S(G29), .Z(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G26), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  OR2_X1    g289(.A1(G104), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n716));
  INV_X1    g291(.A(G140), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n489), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G128), .B2(new_n620), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n714), .B1(new_n719), .B2(new_n712), .ZN(new_n720));
  INV_X1    g295(.A(G2067), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n712), .A2(G35), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G162), .B2(new_n712), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT29), .B(G2090), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n693), .A2(new_n710), .A3(new_n722), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT24), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(G34), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(G34), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n729), .A2(new_n730), .A3(new_n712), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n478), .B2(new_n712), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT90), .B(G2084), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT23), .ZN(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI22_X1  g312(.A1(G299), .A2(G16), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1956), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n727), .A2(new_n734), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n736), .A2(G5), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G171), .B2(new_n736), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1961), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G29), .B2(new_n625), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n712), .A2(G27), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G164), .B2(new_n712), .ZN(new_n747));
  INV_X1    g322(.A(G2078), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT30), .B(G28), .Z(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(G29), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G19), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n560), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1341), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n691), .A2(G2072), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n751), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G286), .A2(new_n736), .ZN(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G21), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n757), .A2(KEYINPUT95), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(KEYINPUT95), .B2(new_n757), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n741), .A2(new_n745), .A3(new_n756), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G24), .ZN(new_n764));
  INV_X1    g339(.A(G290), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT85), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1986), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n712), .A2(G25), .ZN(new_n769));
  INV_X1    g344(.A(G131), .ZN(new_n770));
  NOR2_X1   g345(.A1(G95), .A2(G2105), .ZN(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n489), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G119), .B2(new_n620), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n769), .B1(new_n774), .B2(new_n712), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT35), .B(G1991), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n768), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n736), .A2(G23), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G288), .B2(G16), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(KEYINPUT87), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT33), .B(G1976), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n785), .B(new_n780), .C1(G288), .C2(G16), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n783), .A2(new_n784), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n736), .A2(G22), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G166), .B2(new_n736), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1971), .Z(new_n791));
  INV_X1    g366(.A(new_n784), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n782), .B2(new_n786), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n736), .A2(G6), .ZN(new_n794));
  INV_X1    g369(.A(G305), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n736), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n788), .A2(new_n791), .A3(new_n793), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n779), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT36), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n779), .B(new_n805), .C1(new_n801), .C2(new_n802), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n763), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n736), .A2(G4), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n608), .B2(new_n736), .ZN(new_n809));
  INV_X1    g384(.A(G1348), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n760), .A2(new_n761), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT96), .Z(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT31), .B(G11), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n807), .A2(new_n811), .A3(new_n813), .A4(new_n814), .ZN(G150));
  NAND2_X1  g390(.A1(G150), .A2(KEYINPUT97), .ZN(new_n816));
  INV_X1    g391(.A(new_n814), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n817), .B(new_n763), .C1(new_n804), .C2(new_n806), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n818), .A2(new_n819), .A3(new_n811), .A4(new_n813), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n816), .A2(new_n820), .ZN(G311));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  INV_X1    g397(.A(G55), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n523), .A2(new_n822), .B1(new_n525), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n520), .ZN(new_n826));
  OAI21_X1  g401(.A(G860), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NOR2_X1   g403(.A1(new_n824), .A2(new_n826), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n557), .B2(new_n559), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n558), .A2(new_n553), .A3(new_n551), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n829), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n608), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n828), .B1(new_n840), .B2(G860), .ZN(G145));
  XOR2_X1   g416(.A(new_n774), .B(new_n628), .Z(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n719), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n707), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n719), .A2(new_n701), .A3(new_n706), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(G164), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(G164), .B1(new_n845), .B2(new_n846), .ZN(new_n849));
  OAI211_X1 g424(.A(KEYINPUT99), .B(new_n690), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n472), .A2(G142), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n620), .A2(G130), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n855), .B(new_n856), .C1(G118), .C2(new_n463), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n851), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n845), .A2(new_n846), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n509), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n690), .A2(KEYINPUT99), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n690), .A2(KEYINPUT99), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n847), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n850), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n858), .B1(new_n850), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n843), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n850), .A2(new_n863), .ZN(new_n867));
  INV_X1    g442(.A(new_n858), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n850), .A2(new_n858), .A3(new_n863), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n869), .A2(new_n842), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n866), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(G162), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n866), .A2(new_n871), .A3(new_n872), .A4(new_n491), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n478), .B(new_n625), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  INV_X1    g454(.A(new_n877), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(new_n880), .A3(new_n875), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT40), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n878), .A2(new_n884), .A3(new_n879), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(G395));
  XNOR2_X1  g461(.A(new_n836), .B(new_n615), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n608), .A2(G299), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n607), .A2(new_n575), .A3(new_n568), .A4(new_n573), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n890), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(new_n894), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n888), .A2(KEYINPUT41), .A3(new_n889), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(KEYINPUT102), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n887), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n892), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G288), .B(G166), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n765), .ZN(new_n902));
  XNOR2_X1  g477(.A(G288), .B(G303), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G290), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G305), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n904), .A3(new_n795), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n900), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n892), .A2(new_n909), .A3(new_n899), .A4(new_n911), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(G868), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT103), .B1(new_n829), .B2(G868), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n913), .A2(KEYINPUT103), .A3(G868), .A4(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(G295));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n917), .A2(new_n920), .A3(new_n918), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n917), .B2(new_n918), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(G331));
  AOI21_X1  g498(.A(G301), .B1(new_n834), .B2(new_n835), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n830), .A2(new_n833), .ZN(new_n925));
  AOI211_X1 g500(.A(new_n831), .B(new_n829), .C1(new_n557), .C2(new_n559), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n925), .A2(new_n926), .A3(G171), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n924), .A2(new_n927), .A3(G286), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n834), .A2(G301), .A3(new_n835), .ZN(new_n929));
  OAI21_X1  g504(.A(G171), .B1(new_n925), .B2(new_n926), .ZN(new_n930));
  AOI21_X1  g505(.A(G168), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n895), .B(new_n898), .C1(new_n928), .C2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(G286), .B1(new_n924), .B2(new_n927), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(G168), .A3(new_n930), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n890), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n908), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n879), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n896), .A2(new_n897), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n928), .B2(new_n931), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n908), .B1(new_n939), .B2(new_n935), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n908), .B1(new_n932), .B2(new_n935), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(KEYINPUT105), .B(KEYINPUT43), .C1(new_n937), .C2(new_n940), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n943), .A2(new_n947), .A3(KEYINPUT44), .A4(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n937), .B2(new_n944), .ZN(new_n950));
  INV_X1    g525(.A(new_n940), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(new_n946), .A3(new_n879), .A4(new_n936), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(KEYINPUT44), .B2(new_n953), .ZN(G397));
  INV_X1    g529(.A(KEYINPUT118), .ZN(new_n955));
  AND4_X1   g530(.A1(G40), .A2(new_n466), .A3(new_n473), .A4(new_n476), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n497), .B1(new_n488), .B2(new_n494), .ZN(new_n959));
  INV_X1    g534(.A(new_n501), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n504), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n506), .A2(new_n508), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n509), .A2(new_n965), .A3(new_n958), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n957), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT58), .B(G1341), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n955), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n509), .A2(new_n965), .A3(new_n958), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n965), .B1(new_n509), .B2(new_n958), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n956), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n968), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(KEYINPUT118), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT45), .B(new_n958), .C1(new_n961), .C2(new_n962), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n956), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT45), .B1(new_n509), .B2(new_n958), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1996), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR4_X1   g556(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT117), .A4(G1996), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n969), .B(new_n974), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT59), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n983), .B(new_n560), .C1(KEYINPUT119), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n560), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n964), .A2(new_n966), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n957), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n992));
  AOI211_X1 g567(.A(new_n992), .B(new_n990), .C1(new_n509), .C2(new_n958), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT109), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(G1348), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n972), .A2(G2067), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n608), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n990), .B1(new_n970), .B2(new_n971), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(new_n956), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n810), .ZN(new_n1001));
  INV_X1    g576(.A(new_n997), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n607), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n985), .A2(new_n988), .B1(new_n1004), .B2(KEYINPUT60), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n1006));
  OR3_X1    g581(.A1(G299), .A2(KEYINPUT116), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT116), .B1(G299), .B2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n568), .A2(new_n575), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n568), .A2(KEYINPUT115), .A3(new_n575), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n573), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n1006), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n964), .A2(KEYINPUT50), .A3(new_n966), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n990), .B(new_n958), .C1(new_n961), .C2(new_n962), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT111), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n509), .A2(new_n1020), .A3(new_n990), .A4(new_n958), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(new_n1022), .A3(new_n956), .ZN(new_n1023));
  INV_X1    g598(.A(G1956), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n979), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1016), .A2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1023), .A2(new_n1024), .B1(new_n979), .B2(new_n1026), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(KEYINPUT120), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT61), .ZN(new_n1034));
  OR3_X1    g609(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT120), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OR4_X1    g611(.A1(KEYINPUT60), .A2(new_n996), .A3(new_n607), .A4(new_n997), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1032), .A2(KEYINPUT121), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1030), .A2(new_n1031), .A3(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1038), .A2(KEYINPUT61), .A3(new_n1029), .A4(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1005), .A2(new_n1036), .A3(new_n1037), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1029), .A2(new_n998), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n1032), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G2090), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1017), .A2(new_n1022), .A3(new_n1046), .A4(new_n956), .ZN(new_n1047));
  XOR2_X1   g622(.A(KEYINPUT107), .B(G1971), .Z(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n977), .B2(new_n978), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G8), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G303), .A2(G8), .ZN(new_n1052));
  XOR2_X1   g627(.A(new_n1052), .B(KEYINPUT55), .Z(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n995), .A2(new_n1046), .A3(new_n956), .A4(new_n999), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1049), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(G8), .A3(new_n1053), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n578), .A2(G1976), .A3(new_n579), .A4(new_n580), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n972), .A2(G8), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT52), .ZN(new_n1061));
  INV_X1    g636(.A(G1981), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(new_n587), .C1(new_n589), .C2(new_n590), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n516), .A2(new_n522), .A3(G86), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT110), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1064), .A2(new_n585), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1064), .B2(new_n585), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n584), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1063), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1063), .B(KEYINPUT49), .C1(new_n1062), .C2(new_n1068), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(G8), .A3(new_n972), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1976), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n972), .A2(new_n1075), .A3(G8), .A4(new_n1059), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1061), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1055), .A2(new_n1058), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1055), .A2(new_n1058), .A3(KEYINPUT124), .A4(new_n1077), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT45), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n761), .B1(new_n1083), .B2(new_n977), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1000), .B2(G2084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G286), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1084), .B(G168), .C1(new_n1000), .C2(G2084), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1086), .A2(KEYINPUT51), .A3(G8), .A4(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(G8), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT122), .B(G1961), .Z(new_n1092));
  NAND2_X1  g667(.A1(new_n1000), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  INV_X1    g669(.A(new_n979), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(G2078), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1083), .A2(new_n977), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n748), .A2(KEYINPUT53), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1093), .B(new_n1096), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G171), .B(KEYINPUT54), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1088), .A2(new_n1091), .A3(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1093), .B(KEYINPUT123), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n979), .A2(KEYINPUT53), .A3(new_n748), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(new_n1100), .A3(new_n1096), .A4(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1082), .A2(new_n1103), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1045), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1058), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1085), .A2(G8), .A3(G168), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT113), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1057), .A2(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1054), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1112), .B1(new_n1114), .B2(new_n1077), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1053), .B1(new_n1057), .B2(G8), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1061), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1116), .A2(KEYINPUT113), .A3(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(KEYINPUT63), .B(new_n1111), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT114), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT112), .B(KEYINPUT63), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1078), .B2(new_n1110), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1114), .A2(new_n1112), .A3(new_n1077), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT113), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(KEYINPUT63), .A4(new_n1111), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1120), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1063), .B1(new_n1129), .B2(G288), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(G8), .A3(new_n972), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1058), .B2(new_n1117), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1088), .A2(new_n1091), .A3(KEYINPUT62), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT62), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1099), .A2(G171), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1108), .A2(new_n1128), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n978), .A2(new_n956), .ZN(new_n1140));
  INV_X1    g715(.A(new_n776), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n774), .A2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n774), .A2(new_n1141), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT45), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n963), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n957), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n980), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT106), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT106), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1150), .A3(new_n980), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n706), .A3(new_n701), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n719), .B(new_n721), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(G1996), .B2(new_n707), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1140), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G290), .B(G1986), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n1144), .B(new_n1156), .C1(new_n1147), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1139), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT46), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1152), .B(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1147), .B1(new_n1154), .B2(new_n707), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT126), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1161), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT47), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1142), .B(KEYINPUT125), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1156), .A2(new_n1170), .B1(G2067), .B2(new_n844), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1156), .A2(new_n1144), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1140), .A2(G1986), .A3(G290), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT48), .Z(new_n1174));
  AOI22_X1  g749(.A1(new_n1171), .A2(new_n1147), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1164), .A2(KEYINPUT47), .A3(new_n1166), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1169), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1169), .A2(new_n1175), .A3(KEYINPUT127), .A4(new_n1176), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1159), .A2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g757(.A(new_n460), .B(G229), .C1(new_n950), .C2(new_n952), .ZN(new_n1184));
  NOR2_X1   g758(.A1(new_n647), .A2(G227), .ZN(new_n1185));
  AND3_X1   g759(.A1(new_n1184), .A2(new_n882), .A3(new_n1185), .ZN(G308));
  NAND3_X1  g760(.A1(new_n1184), .A2(new_n882), .A3(new_n1185), .ZN(G225));
endmodule


