//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n442, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n577, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n641, new_n644, new_n645, new_n647,
    new_n648, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1241, new_n1242;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G108), .ZN(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(new_n442), .A2(G57), .A3(G69), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT69), .Z(G319));
  NAND2_X1  g036(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(KEYINPUT72), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n463), .A2(new_n467), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n472), .B1(new_n479), .B2(G125), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT71), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n483));
  INV_X1    g058(.A(G125), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n474), .B2(new_n478), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n483), .B(G2105), .C1(new_n485), .C2(new_n472), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n470), .B1(new_n482), .B2(new_n486), .ZN(G160));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n466), .B2(G136), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n481), .B1(new_n464), .B2(new_n465), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(new_n465), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT3), .B1(KEYINPUT72), .B2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n481), .A2(G114), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n498), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n503), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n479), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n481), .B1(new_n496), .B2(new_n497), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n506), .B2(new_n503), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n505), .B2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT73), .B(KEYINPUT6), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT74), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n513), .B(G651), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(G543), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n519), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n511), .A2(new_n512), .A3(new_n518), .A4(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n510), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n511), .A2(G543), .A3(new_n518), .A4(new_n512), .ZN(new_n530));
  INV_X1    g105(.A(G50), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G166));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n525), .A2(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n526), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G51), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n530), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n522), .A2(G543), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n519), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n545));
  AOI21_X1  g120(.A(KEYINPUT75), .B1(new_n519), .B2(KEYINPUT5), .ZN(new_n546));
  OAI211_X1 g121(.A(G64), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(G77), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI221_X1 g127(.A(new_n550), .B1(new_n530), .B2(new_n551), .C1(new_n552), .C2(new_n526), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  OAI211_X1 g129(.A(G56), .B(new_n544), .C1(new_n545), .C2(new_n546), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n555), .A2(KEYINPUT76), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT76), .B1(new_n555), .B2(new_n556), .ZN(new_n558));
  NOR3_X1   g133(.A1(new_n557), .A2(new_n558), .A3(new_n510), .ZN(new_n559));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  OAI22_X1  g136(.A1(new_n560), .A2(new_n530), .B1(new_n526), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT77), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n558), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n555), .A2(KEYINPUT76), .A3(new_n556), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(G651), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n530), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G43), .ZN(new_n568));
  INV_X1    g143(.A(new_n526), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G81), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n566), .A2(new_n568), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n563), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  AND3_X1   g149(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G36), .ZN(G176));
  NAND2_X1  g151(.A1(G1), .A2(G3), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT8), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT78), .ZN(G188));
  NAND2_X1  g155(.A1(new_n569), .A2(G91), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n510), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n530), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n584), .B1(new_n586), .B2(G53), .ZN(new_n587));
  INV_X1    g162(.A(G53), .ZN(new_n588));
  NOR4_X1   g163(.A1(new_n530), .A2(new_n585), .A3(KEYINPUT9), .A4(new_n588), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n581), .B(new_n583), .C1(new_n587), .C2(new_n589), .ZN(G299));
  NAND2_X1  g165(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n513), .B1(new_n593), .B2(G651), .ZN(new_n594));
  AOI211_X1 g169(.A(KEYINPUT74), .B(new_n510), .C1(new_n591), .C2(new_n592), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n596), .A2(G51), .A3(G543), .A4(new_n512), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n596), .A2(G89), .A3(new_n512), .A4(new_n525), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT80), .A4(new_n538), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n540), .B2(new_n542), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(G286));
  OR2_X1    g177(.A1(new_n529), .A2(new_n532), .ZN(G303));
  AND2_X1   g178(.A1(new_n567), .A2(G49), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n605));
  INV_X1    g180(.A(G87), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n526), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G288));
  NAND2_X1  g184(.A1(G73), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n611));
  INV_X1    g186(.A(G61), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G651), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT81), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n613), .A2(new_n616), .A3(G651), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G48), .ZN(new_n619));
  INV_X1    g194(.A(G86), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n619), .A2(new_n530), .B1(new_n526), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n622), .ZN(G305));
  AND2_X1   g198(.A1(new_n569), .A2(G85), .ZN(new_n624));
  INV_X1    g199(.A(G47), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n626));
  OAI22_X1  g201(.A1(new_n530), .A2(new_n625), .B1(new_n626), .B2(new_n510), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(G290));
  NAND2_X1  g204(.A1(G301), .A2(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(G79), .A2(G543), .ZN(new_n631));
  INV_X1    g206(.A(G66), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n611), .B2(new_n632), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n567), .A2(G54), .B1(G651), .B2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G92), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n526), .A2(KEYINPUT10), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT10), .B1(new_n526), .B2(new_n635), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n630), .B1(new_n638), .B2(G868), .ZN(G284));
  OAI21_X1  g214(.A(new_n630), .B1(new_n638), .B2(G868), .ZN(G321));
  INV_X1    g215(.A(G868), .ZN(new_n641));
  MUX2_X1   g216(.A(G286), .B(G299), .S(new_n641), .Z(G297));
  MUX2_X1   g217(.A(G286), .B(G299), .S(new_n641), .Z(G280));
  XNOR2_X1  g218(.A(KEYINPUT82), .B(G559), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n638), .B1(G860), .B2(new_n645), .ZN(G148));
  NAND2_X1  g221(.A1(new_n638), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G868), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(G868), .B2(new_n573), .ZN(G323));
  XNOR2_X1  g224(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g225(.A1(new_n479), .A2(new_n468), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT12), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n492), .A2(G123), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n466), .A2(G135), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n481), .A2(G111), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n655), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(G2096), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n660), .ZN(G156));
  XNOR2_X1  g236(.A(G2427), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT85), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2451), .B(G2454), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1341), .B(G1348), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  AND2_X1   g251(.A1(new_n676), .A2(G14), .ZN(G401));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  XOR2_X1   g254(.A(G2067), .B(G2678), .Z(new_n680));
  AOI21_X1  g255(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n679), .B(KEYINPUT17), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n681), .B1(new_n683), .B2(new_n680), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT86), .Z(new_n685));
  INV_X1    g260(.A(new_n679), .ZN(new_n686));
  INV_X1    g261(.A(new_n680), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(new_n687), .A3(new_n678), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT18), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n683), .A2(new_n678), .A3(new_n680), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n685), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G2096), .B(G2100), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G227));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT87), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n695), .A2(KEYINPUT88), .A3(new_n696), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n695), .A2(new_n696), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n708), .A2(new_n697), .A3(new_n701), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n706), .B(new_n709), .C1(new_n701), .C2(new_n708), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  INV_X1    g288(.A(G1981), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1986), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n712), .B(new_n716), .ZN(G229));
  XNOR2_X1  g292(.A(KEYINPUT31), .B(G11), .ZN(new_n718));
  NAND2_X1  g293(.A1(G299), .A2(G16), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n720), .A2(KEYINPUT23), .A3(G20), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT23), .ZN(new_n722));
  INV_X1    g297(.A(G20), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(G16), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1956), .ZN(new_n726));
  OAI21_X1  g301(.A(KEYINPUT94), .B1(G5), .B2(G16), .ZN(new_n727));
  OR3_X1    g302(.A1(KEYINPUT94), .A2(G5), .A3(G16), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n727), .B(new_n728), .C1(G301), .C2(new_n720), .ZN(new_n729));
  INV_X1    g304(.A(G1961), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G26), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n492), .A2(G128), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT93), .Z(new_n736));
  NOR2_X1   g311(.A1(new_n481), .A2(G116), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n466), .B2(G140), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n734), .B1(new_n741), .B2(G29), .ZN(new_n742));
  MUX2_X1   g317(.A(new_n734), .B(new_n742), .S(KEYINPUT28), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2067), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n745), .ZN(new_n747));
  MUX2_X1   g322(.A(new_n746), .B(new_n747), .S(KEYINPUT95), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n720), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n720), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n749), .A2(G2090), .B1(G1966), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(G1966), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(G164), .A2(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G27), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n466), .A2(G139), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n468), .A2(G103), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  AOI22_X1  g336(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n759), .B(new_n761), .C1(new_n762), .C2(new_n481), .ZN(new_n763));
  MUX2_X1   g338(.A(G33), .B(new_n763), .S(G29), .Z(new_n764));
  AOI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(G2072), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n766), .A2(new_n745), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G160), .B2(new_n745), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(G2084), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n764), .A2(G2072), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n765), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n744), .A2(new_n752), .A3(new_n754), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(G2084), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n492), .A2(G129), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT26), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n466), .A2(G141), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n468), .A2(G105), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n775), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G32), .B(new_n780), .S(G29), .Z(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT27), .B(G1996), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n756), .A2(new_n757), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(G28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(G28), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n786), .A2(new_n787), .A3(new_n745), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n774), .A2(new_n783), .A3(new_n784), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G19), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n573), .B2(G16), .ZN(new_n791));
  INV_X1    g366(.A(G1341), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n794), .A2(new_n795), .B1(new_n749), .B2(G2090), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n732), .A2(new_n773), .A3(new_n789), .A4(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n720), .B1(new_n618), .B2(new_n622), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n720), .A2(G6), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(KEYINPUT92), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n799), .A2(KEYINPUT92), .A3(new_n801), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT32), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT32), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n799), .A2(KEYINPUT92), .A3(new_n801), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n802), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n714), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G23), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n608), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT33), .B(G1976), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n720), .A2(G22), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G166), .B2(new_n720), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1971), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT32), .B1(new_n803), .B2(new_n804), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n807), .A2(new_n802), .A3(new_n806), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n818), .A2(new_n819), .A3(G1981), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n809), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT34), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n809), .A2(new_n817), .A3(KEYINPUT34), .A4(new_n820), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n745), .A2(G25), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n492), .A2(G119), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n466), .A2(G131), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n481), .A2(G107), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT90), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n826), .B1(new_n835), .B2(new_n745), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT35), .B(G1991), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT91), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G16), .A2(G24), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n628), .B2(G16), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(G1986), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(G1986), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n798), .B1(new_n825), .B2(new_n845), .ZN(new_n846));
  AOI211_X1 g421(.A(KEYINPUT36), .B(new_n844), .C1(new_n823), .C2(new_n824), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n718), .B(new_n797), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n720), .A2(G4), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n638), .B2(new_n720), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G1348), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n659), .A2(new_n745), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(G311));
  INV_X1    g428(.A(new_n797), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n825), .A2(new_n845), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT36), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n825), .A2(new_n798), .A3(new_n845), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n851), .ZN(new_n859));
  INV_X1    g434(.A(new_n852), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n718), .ZN(G150));
  NAND2_X1  g436(.A1(new_n569), .A2(G93), .ZN(new_n862));
  AND2_X1   g437(.A1(G80), .A2(G543), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n525), .B2(G67), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(new_n510), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n596), .A2(G55), .A3(G543), .A4(new_n512), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n862), .A2(new_n866), .A3(KEYINPUT97), .A4(new_n865), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n869));
  INV_X1    g444(.A(G55), .ZN(new_n870));
  OAI22_X1  g445(.A1(new_n530), .A2(new_n870), .B1(new_n510), .B2(new_n864), .ZN(new_n871));
  INV_X1    g446(.A(G93), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n526), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n566), .A2(new_n568), .A3(new_n570), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n573), .A2(new_n867), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n638), .A2(G559), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT98), .Z(new_n884));
  AOI21_X1  g459(.A(G860), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n868), .A2(new_n874), .A3(G860), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(KEYINPUT37), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(G145));
  XNOR2_X1  g464(.A(new_n741), .B(G164), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n763), .B(new_n780), .Z(new_n891));
  XOR2_X1   g466(.A(new_n890), .B(new_n891), .Z(new_n892));
  INV_X1    g467(.A(new_n652), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n835), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n833), .A2(new_n834), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n652), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT99), .B1(new_n481), .B2(G118), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n481), .A2(KEYINPUT99), .A3(G118), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n899), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n466), .A2(G142), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n492), .A2(G130), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n894), .A2(new_n896), .A3(new_n907), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  OR3_X1    g488(.A1(new_n892), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n659), .B(new_n494), .ZN(new_n915));
  XOR2_X1   g490(.A(G160), .B(new_n915), .Z(new_n916));
  OAI21_X1  g491(.A(new_n892), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G37), .ZN(new_n919));
  INV_X1    g494(.A(new_n892), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n920), .B(new_n921), .C1(new_n912), .C2(new_n913), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n912), .B2(new_n913), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n892), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n918), .B(new_n919), .C1(new_n925), .C2(new_n916), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g502(.A1(G290), .A2(new_n608), .ZN(new_n928));
  NAND2_X1  g503(.A1(G288), .A2(new_n628), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n932));
  XNOR2_X1  g507(.A(G305), .B(G166), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(new_n930), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n933), .A3(KEYINPUT105), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT42), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n573), .A2(new_n867), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n875), .A2(new_n876), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(new_n647), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n567), .A2(KEYINPUT79), .A3(G53), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT9), .ZN(new_n945));
  INV_X1    g520(.A(new_n589), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n638), .A2(new_n947), .A3(new_n581), .A4(new_n583), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n949));
  NAND2_X1  g524(.A1(G299), .A2(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n948), .A2(KEYINPUT41), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT41), .B1(new_n948), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n943), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT104), .ZN(new_n955));
  INV_X1    g530(.A(new_n943), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n948), .A2(new_n950), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n943), .A2(new_n959), .A3(new_n953), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n955), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n939), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n939), .A2(new_n961), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n641), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n964), .A2(new_n966), .B1(new_n641), .B2(new_n875), .ZN(G295));
  AOI22_X1  g542(.A1(new_n964), .A2(new_n966), .B1(new_n641), .B2(new_n875), .ZN(G331));
  XOR2_X1   g543(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n969));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n971), .B(G301), .C1(new_n601), .C2(new_n599), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT109), .B1(G286), .B2(G171), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G301), .A2(G168), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(G301), .A2(G168), .A3(KEYINPUT108), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n877), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(G286), .A2(G171), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n971), .ZN(new_n982));
  NAND3_X1  g557(.A1(G286), .A2(KEYINPUT109), .A3(G171), .ZN(new_n983));
  AND4_X1   g558(.A1(new_n877), .A2(new_n982), .A3(new_n983), .A4(new_n979), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n953), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n936), .A2(new_n937), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(new_n983), .A3(new_n979), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n942), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n974), .A2(new_n877), .A3(new_n979), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n957), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(KEYINPUT110), .A3(new_n953), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n987), .A2(new_n988), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n995), .A2(new_n919), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n987), .A2(new_n992), .A3(new_n994), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n938), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n970), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n992), .B1(new_n985), .B2(KEYINPUT111), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n993), .B2(new_n953), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n938), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AND4_X1   g578(.A1(new_n970), .A2(new_n1003), .A3(new_n919), .A4(new_n995), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n969), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n996), .A2(new_n970), .A3(new_n998), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1003), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n995), .A2(new_n919), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT43), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1009), .A3(KEYINPUT44), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1005), .A2(new_n1010), .ZN(G397));
  INV_X1    g586(.A(G2067), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n741), .B(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1996), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n780), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n895), .A2(new_n837), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n895), .A2(new_n837), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(G290), .A2(G1986), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G290), .A2(G1986), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT113), .B(G40), .Z(new_n1023));
  AOI211_X1 g598(.A(new_n470), .B(new_n1023), .C1(new_n482), .C2(new_n486), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n501), .A2(new_n500), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n492), .B2(G126), .ZN(new_n1026));
  INV_X1    g601(.A(new_n504), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n474), .B2(new_n478), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT4), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n466), .B2(G138), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1026), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT112), .B(G1384), .Z(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1024), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1022), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G164), .A2(G1384), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1024), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(G288), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n608), .A2(KEYINPUT117), .A3(G1976), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT52), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n618), .A2(new_n622), .A3(new_n714), .ZN(new_n1047));
  INV_X1    g622(.A(new_n614), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n621), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1047), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1040), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1043), .A2(new_n1040), .A3(new_n1055), .A4(new_n1044), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1046), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT114), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n1060));
  NAND4_X1  g635(.A1(G303), .A2(new_n1060), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1063), .A2(KEYINPUT115), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(KEYINPUT115), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1023), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT45), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(G164), .B2(G1384), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1031), .A2(KEYINPUT45), .A3(new_n1033), .ZN(new_n1070));
  NAND4_X1  g645(.A1(G160), .A2(new_n1067), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1971), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n1074));
  INV_X1    g649(.A(G1384), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1031), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1031), .B2(new_n1075), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G2090), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1024), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1038), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1066), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1066), .A2(KEYINPUT116), .A3(new_n1082), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1057), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1066), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1024), .A2(new_n1079), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1080), .B1(new_n1090), .B2(KEYINPUT118), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n479), .A2(G125), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n471), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n483), .B1(new_n1093), .B2(G2105), .ZN(new_n1094));
  INV_X1    g669(.A(new_n486), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n469), .B(new_n1067), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1076), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1089), .B(new_n1073), .C1(new_n1091), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G8), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1090), .A2(KEYINPUT118), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n1080), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1089), .B1(new_n1106), .B2(new_n1073), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1088), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1087), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G2084), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1039), .A2(KEYINPUT45), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1111), .A2(G160), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1112));
  INV_X1    g687(.A(G1966), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1099), .A2(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT51), .B1(new_n1114), .B2(G168), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1038), .B1(new_n1114), .B2(G168), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1116), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT126), .B(KEYINPUT54), .Z(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1071), .B2(G2078), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1090), .A2(new_n730), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(G160), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1121), .A2(G2078), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1111), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(G301), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1070), .A2(new_n469), .ZN(new_n1129));
  INV_X1    g704(.A(G40), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1034), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1093), .A2(G2105), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .A4(new_n1126), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1122), .A2(new_n1123), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(G171), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1120), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1124), .A2(G301), .A3(new_n1127), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(G171), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(KEYINPUT54), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1119), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT56), .B(G2072), .Z(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1125), .A2(new_n1141), .A3(new_n1070), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G1956), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1090), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT121), .B1(new_n1071), .B2(new_n1142), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(KEYINPUT57), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1149), .A2(KEYINPUT57), .ZN(new_n1151));
  OR3_X1    g726(.A1(G299), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n1153));
  NAND3_X1  g728(.A1(G299), .A2(new_n1149), .A3(KEYINPUT57), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1153), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1148), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT124), .ZN(new_n1158));
  AOI21_X1  g733(.A(G1348), .B1(new_n1024), .B2(new_n1079), .ZN(new_n1159));
  NAND4_X1  g734(.A1(G160), .A2(new_n1012), .A3(new_n1067), .A4(new_n1039), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT122), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(G1348), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1164), .A2(new_n1165), .A3(new_n1160), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(new_n638), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1168), .B(new_n1148), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1158), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1148), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n638), .A2(KEYINPUT125), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1164), .A2(new_n1165), .A3(new_n1160), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1165), .B1(new_n1164), .B2(new_n1160), .ZN(new_n1176));
  OAI211_X1 g751(.A(KEYINPUT60), .B(new_n1174), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n638), .A2(KEYINPUT125), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  OR3_X1    g755(.A1(new_n1175), .A2(new_n1176), .A3(KEYINPUT60), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1182), .A2(KEYINPUT60), .A3(new_n1178), .A4(new_n1174), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1125), .A2(new_n1014), .A3(new_n1070), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1024), .A2(new_n1039), .ZN(new_n1186));
  XOR2_X1   g761(.A(KEYINPUT58), .B(G1341), .Z(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1185), .A2(new_n1188), .B1(new_n563), .B2(new_n572), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT59), .Z(new_n1190));
  AND2_X1   g765(.A1(new_n1148), .A2(new_n1171), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1172), .B1(new_n1191), .B2(KEYINPUT61), .ZN(new_n1192));
  OR3_X1    g767(.A1(new_n1148), .A2(new_n1171), .A3(KEYINPUT61), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1184), .A2(new_n1190), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI211_X1 g769(.A(new_n1109), .B(new_n1140), .C1(new_n1173), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1057), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1114), .A2(new_n1038), .A3(G286), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT63), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1073), .B1(new_n1091), .B2(new_n1101), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT119), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1201), .A2(G8), .A3(new_n1102), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1199), .B1(new_n1202), .B2(new_n1088), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1196), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1196), .B(new_n1197), .C1(new_n1082), .C2(new_n1066), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1054), .A2(new_n1042), .A3(new_n608), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1047), .ZN(new_n1208));
  AOI22_X1  g783(.A1(new_n1206), .A2(KEYINPUT63), .B1(new_n1040), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1119), .A2(KEYINPUT62), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1210), .A2(new_n1108), .A3(new_n1087), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1128), .B1(new_n1119), .B2(KEYINPUT62), .ZN(new_n1212));
  OAI211_X1 g787(.A(new_n1205), .B(new_n1209), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1037), .B1(new_n1195), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1035), .A2(G1996), .ZN(new_n1215));
  OR2_X1    g790(.A1(new_n1215), .A2(KEYINPUT46), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1013), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1036), .B1(new_n1217), .B2(new_n780), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1215), .A2(KEYINPUT46), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1216), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT47), .Z(new_n1221));
  NOR2_X1   g796(.A1(new_n1020), .A2(new_n1035), .ZN(new_n1222));
  XOR2_X1   g797(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1223));
  XNOR2_X1  g798(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(new_n1019), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1224), .B1(new_n1225), .B2(new_n1036), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1013), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n736), .A2(new_n1012), .A3(new_n740), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1035), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NOR3_X1   g804(.A1(new_n1221), .A2(new_n1226), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1214), .A2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g806(.A(G319), .ZN(new_n1233));
  OR2_X1    g807(.A1(G229), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g808(.A(G227), .B1(new_n676), .B2(G14), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n926), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g810(.A(new_n998), .ZN(new_n1237));
  OAI21_X1  g811(.A(KEYINPUT43), .B1(new_n1237), .B2(new_n1008), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n996), .A2(new_n970), .A3(new_n1003), .ZN(new_n1239));
  AOI211_X1 g813(.A(new_n1234), .B(new_n1236), .C1(new_n1238), .C2(new_n1239), .ZN(G308));
  AOI21_X1  g814(.A(new_n1234), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1241));
  INV_X1    g815(.A(new_n1236), .ZN(new_n1242));
  NAND2_X1  g816(.A1(new_n1241), .A2(new_n1242), .ZN(G225));
endmodule


