//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1188, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  INV_X1    g0029(.A(G238), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n228), .B1(new_n202), .B2(new_n229), .C1(new_n203), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n213), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n216), .B(new_n221), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n229), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT64), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G223), .A2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G222), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n256), .B(new_n257), .C1(new_n258), .C2(G1698), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n259), .B(new_n260), .C1(G77), .C2(new_n256), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n263), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(G226), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G190), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(G200), .B2(new_n268), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n219), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n210), .B2(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G50), .ZN(new_n275));
  INV_X1    g0075(.A(G13), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(G50), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n204), .A2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(G150), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n253), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n280), .B1(new_n281), .B2(new_n283), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n279), .B1(new_n273), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT9), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n271), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT10), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n268), .A2(G179), .ZN(new_n293));
  AOI21_X1  g0093(.A(G169), .B1(new_n261), .B2(new_n267), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n293), .A2(new_n288), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G238), .A2(G1698), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n256), .B(new_n298), .C1(new_n229), .C2(G1698), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n260), .C1(G107), .C2(new_n256), .ZN(new_n300));
  INV_X1    g0100(.A(new_n264), .ZN(new_n301));
  INV_X1    g0101(.A(new_n266), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n300), .B(new_n301), .C1(new_n224), .C2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT65), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G200), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n274), .A2(G77), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G77), .B2(new_n278), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT15), .B(G87), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n283), .B2(new_n284), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n307), .B1(new_n273), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n305), .B(new_n312), .C1(new_n269), .C2(new_n304), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n304), .A2(G179), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n304), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n297), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n264), .B1(G232), .B2(new_n266), .ZN(new_n319));
  INV_X1    g0119(.A(new_n260), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT67), .B(G33), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(KEYINPUT3), .ZN(new_n323));
  MUX2_X1   g0123(.A(G223), .B(G226), .S(G1698), .Z(new_n324));
  AOI22_X1  g0124(.A1(new_n323), .A2(new_n324), .B1(G33), .B2(G87), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n319), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G87), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n320), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n301), .B1(new_n302), .B2(new_n229), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT69), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT69), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n319), .B(new_n333), .C1(new_n320), .C2(new_n325), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n327), .B1(new_n335), .B2(new_n315), .ZN(new_n336));
  XNOR2_X1  g0136(.A(G58), .B(G68), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(G20), .B1(G159), .B2(new_n282), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT67), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT3), .ZN(new_n342));
  AOI21_X1  g0142(.A(G20), .B1(new_n342), .B2(new_n252), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n323), .A2(KEYINPUT7), .A3(G20), .ZN(new_n346));
  OAI211_X1 g0146(.A(KEYINPUT16), .B(new_n338), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n338), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n254), .B1(new_n322), .B2(KEYINPUT3), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n344), .A2(G20), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT68), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n251), .A2(G33), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n211), .B1(new_n321), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n354), .B2(new_n344), .ZN(new_n355));
  AOI21_X1  g0155(.A(G20), .B1(new_n252), .B2(new_n254), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n356), .A2(KEYINPUT68), .A3(KEYINPUT7), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n351), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n348), .B1(new_n358), .B2(G68), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n273), .B(new_n347), .C1(new_n359), .C2(KEYINPUT16), .ZN(new_n360));
  INV_X1    g0160(.A(new_n284), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(new_n278), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n274), .B2(new_n361), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n336), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT18), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n332), .A2(new_n368), .A3(new_n334), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n326), .A2(G190), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n360), .B(new_n363), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n301), .B1(new_n302), .B2(new_n230), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G97), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n229), .A2(G1698), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(G226), .B2(G1698), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n375), .B1(new_n377), .B2(new_n255), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n374), .B1(new_n260), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT13), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n379), .B(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n381), .A2(G200), .ZN(new_n382));
  NAND2_X1  g0182(.A1(KEYINPUT66), .A2(KEYINPUT13), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n379), .A2(new_n383), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n384), .A2(G190), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n203), .A2(G20), .ZN(new_n387));
  OAI221_X1 g0187(.A(new_n387), .B1(new_n283), .B2(new_n201), .C1(new_n286), .C2(new_n223), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n273), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT11), .ZN(new_n391));
  INV_X1    g0191(.A(new_n278), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n277), .A2(KEYINPUT12), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n391), .B1(KEYINPUT12), .B2(new_n392), .C1(new_n387), .C2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT12), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n274), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n390), .B2(KEYINPUT11), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n382), .A2(new_n386), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT14), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n381), .A2(new_n402), .A3(G169), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n384), .A2(G179), .A3(new_n385), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n402), .B1(new_n381), .B2(G169), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n399), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n318), .A2(new_n373), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n278), .A2(G97), .ZN(new_n410));
  INV_X1    g0210(.A(new_n273), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n210), .A2(G33), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n278), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n414), .B2(G97), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G97), .A2(G107), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n208), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT6), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT70), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n208), .A2(KEYINPUT70), .A3(new_n418), .A4(new_n416), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n420), .A2(G20), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n282), .A2(G77), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n358), .B2(G107), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n415), .B1(new_n426), .B2(new_n411), .ZN(new_n427));
  INV_X1    g0227(.A(G41), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n428), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT72), .B1(new_n428), .B2(KEYINPUT5), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n210), .B(G45), .C1(new_n428), .C2(KEYINPUT5), .ZN(new_n432));
  OAI211_X1 g0232(.A(G257), .B(new_n320), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT72), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT5), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(G41), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n428), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n260), .A2(new_n262), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT73), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n433), .A2(KEYINPUT73), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n224), .A2(G1698), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(KEYINPUT4), .B1(G250), .B2(G1698), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n448), .B2(new_n255), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n342), .A2(new_n252), .A3(new_n447), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n452), .B2(KEYINPUT71), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT71), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(new_n454), .A3(new_n451), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n320), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n445), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n427), .B1(G190), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT74), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n445), .B2(new_n456), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n452), .A2(KEYINPUT71), .ZN(new_n461));
  INV_X1    g0261(.A(new_n449), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n455), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n260), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n433), .A2(KEYINPUT73), .A3(new_n440), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT73), .B1(new_n433), .B2(new_n440), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n467), .A3(KEYINPUT74), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n460), .A2(new_n468), .A3(G200), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n458), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G179), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n457), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n464), .A2(new_n467), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n315), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n474), .A3(new_n427), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n323), .A2(new_n211), .A3(G68), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT19), .B1(new_n285), .B2(G97), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n225), .A2(new_n206), .A3(new_n207), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT19), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n375), .B2(new_n211), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(new_n273), .B1(new_n392), .B2(new_n308), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n413), .A2(new_n225), .ZN(new_n485));
  XOR2_X1   g0285(.A(new_n485), .B(KEYINPUT76), .Z(new_n486));
  NOR2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G238), .A2(G1698), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n224), .B2(G1698), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n323), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n339), .A2(new_n341), .ZN(new_n491));
  INV_X1    g0291(.A(G116), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT75), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT75), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n320), .B1(new_n490), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n210), .A2(G45), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(G274), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n260), .B(new_n500), .C1(new_n226), .C2(new_n499), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n368), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n498), .A2(new_n269), .A3(new_n501), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(G179), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n315), .B2(new_n502), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n483), .B1(new_n308), .B2(new_n413), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n487), .A2(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n470), .A2(new_n475), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT24), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT78), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n323), .A2(new_n512), .A3(new_n211), .A4(G87), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n342), .A2(new_n211), .A3(G87), .A4(new_n252), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT78), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT22), .ZN(new_n516));
  NOR4_X1   g0316(.A1(new_n255), .A2(KEYINPUT22), .A3(G20), .A4(new_n225), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT79), .B1(new_n211), .B2(G107), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n491), .A2(new_n496), .B1(KEYINPUT79), .B2(KEYINPUT23), .ZN(new_n524));
  OAI221_X1 g0324(.A(new_n522), .B1(new_n207), .B2(new_n523), .C1(new_n524), .C2(G20), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n511), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n514), .B2(KEYINPUT78), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n517), .B1(new_n529), .B2(new_n513), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n530), .A2(KEYINPUT24), .A3(new_n525), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n273), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT80), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT25), .ZN(new_n534));
  AOI211_X1 g0334(.A(G107), .B(new_n278), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n537), .A2(new_n538), .B1(new_n414), .B2(G107), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n342), .A2(new_n252), .ZN(new_n540));
  INV_X1    g0340(.A(G257), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G1698), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(G250), .B2(G1698), .ZN(new_n543));
  INV_X1    g0343(.A(G294), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n540), .A2(new_n543), .B1(new_n544), .B2(new_n322), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n260), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT81), .ZN(new_n547));
  INV_X1    g0347(.A(G264), .ZN(new_n548));
  NOR4_X1   g0348(.A1(new_n438), .A2(new_n547), .A3(new_n548), .A4(new_n260), .ZN(new_n549));
  INV_X1    g0349(.A(new_n432), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n436), .A2(new_n437), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n260), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT81), .B1(new_n552), .B2(G264), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n546), .B(new_n440), .C1(new_n549), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G200), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(G264), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n547), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n552), .A2(KEYINPUT81), .A3(G264), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n557), .A2(new_n558), .B1(new_n260), .B2(new_n545), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(G190), .A3(new_n440), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n532), .A2(new_n539), .A3(new_n555), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n554), .A2(new_n315), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n558), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n471), .A3(new_n440), .A4(new_n546), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n519), .A2(new_n511), .A3(new_n526), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT24), .B1(new_n530), .B2(new_n525), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n411), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n539), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n446), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n273), .B(new_n572), .C1(new_n496), .C2(new_n211), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n573), .B(new_n574), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n413), .A2(new_n492), .B1(new_n278), .B2(new_n496), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G179), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n548), .A2(G1698), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G257), .B2(G1698), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n540), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G303), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n256), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n260), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n552), .A2(G270), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT77), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT77), .B1(new_n552), .B2(G270), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n440), .B(new_n585), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n579), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n315), .B1(new_n575), .B2(new_n577), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT21), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT21), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n590), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n591), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n578), .B1(new_n590), .B2(G200), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n269), .B2(new_n590), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n571), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n409), .A2(new_n510), .A3(new_n601), .ZN(G372));
  INV_X1    g0402(.A(KEYINPUT82), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n570), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n565), .B(KEYINPUT82), .C1(new_n568), .C2(new_n569), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n597), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT83), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n470), .A2(new_n561), .A3(new_n509), .A4(new_n475), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n590), .A2(new_n595), .A3(new_n592), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n595), .B1(new_n590), .B2(new_n592), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n612), .A2(new_n613), .B1(new_n590), .B2(new_n579), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n604), .B2(new_n605), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT83), .B1(new_n615), .B2(new_n609), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n505), .A2(new_n487), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n507), .A2(new_n508), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT26), .B1(new_n619), .B2(new_n475), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n474), .A2(new_n427), .ZN(new_n621));
  XNOR2_X1  g0421(.A(KEYINPUT84), .B(KEYINPUT26), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n509), .A2(new_n621), .A3(new_n472), .A4(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n620), .A2(new_n623), .A3(new_n618), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n611), .A2(new_n616), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n409), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n407), .B1(new_n400), .B2(new_n317), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n372), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n367), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n295), .B1(new_n629), .B2(new_n292), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(G369));
  NAND2_X1  g0431(.A1(new_n277), .A2(new_n211), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n575), .B2(new_n577), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n614), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n600), .B2(new_n639), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G330), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n638), .B1(new_n532), .B2(new_n539), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n571), .A2(new_n645), .B1(new_n570), .B2(new_n638), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n604), .A2(new_n605), .A3(new_n638), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n597), .A2(new_n637), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n570), .A3(new_n561), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(G399));
  NAND2_X1  g0451(.A1(new_n214), .A2(new_n428), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n210), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n478), .A2(G116), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n654), .A2(new_n655), .B1(new_n218), .B2(new_n653), .ZN(new_n656));
  XOR2_X1   g0456(.A(new_n656), .B(KEYINPUT28), .Z(new_n657));
  INV_X1    g0457(.A(KEYINPUT87), .ZN(new_n658));
  INV_X1    g0458(.A(new_n622), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n619), .B2(new_n475), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n509), .A2(new_n621), .A3(new_n661), .A4(new_n472), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n660), .A2(new_n662), .A3(new_n618), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n562), .A2(new_n564), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n532), .B2(new_n539), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT85), .B1(new_n665), .B2(new_n614), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT85), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n597), .A2(new_n570), .A3(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n510), .A2(new_n561), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n663), .B1(new_n669), .B2(KEYINPUT86), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT86), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n610), .A2(new_n671), .A3(new_n668), .A4(new_n666), .ZN(new_n672));
  AOI211_X1 g0472(.A(new_n658), .B(new_n637), .C1(new_n670), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(KEYINPUT86), .ZN(new_n674));
  INV_X1    g0474(.A(new_n663), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT87), .B1(new_n676), .B2(new_n638), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT29), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n625), .A2(new_n638), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n601), .A2(new_n510), .A3(new_n638), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n588), .A2(new_n589), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n498), .A2(new_n471), .A3(new_n501), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n585), .A2(new_n440), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n559), .A4(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT30), .ZN(new_n688));
  OR3_X1    g0488(.A1(new_n687), .A2(new_n688), .A3(new_n473), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n687), .B2(new_n473), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n502), .A2(G179), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n473), .A2(new_n590), .A3(new_n554), .A4(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n637), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n683), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n682), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n657), .B1(new_n701), .B2(G1), .ZN(G364));
  XOR2_X1   g0502(.A(new_n644), .B(KEYINPUT88), .Z(new_n703));
  INV_X1    g0503(.A(G45), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n276), .A2(new_n704), .A3(G20), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT89), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT89), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n654), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n703), .B(new_n708), .C1(G330), .C2(new_n641), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n219), .B1(G20), .B2(new_n315), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT91), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G190), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT33), .B(G317), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n211), .A2(new_n269), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n471), .A2(G200), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n714), .A2(new_n715), .B1(G322), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT92), .Z(new_n721));
  INV_X1    g0521(.A(G283), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n211), .A2(G190), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n368), .A2(G179), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n717), .A2(new_n723), .ZN(new_n726));
  INV_X1    g0526(.A(G311), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n722), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G179), .A2(G200), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n211), .B1(new_n729), .B2(G190), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n716), .A2(new_n724), .ZN(new_n731));
  OAI221_X1 g0531(.A(new_n255), .B1(new_n730), .B2(new_n544), .C1(new_n583), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n723), .A2(new_n729), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n728), .B(new_n732), .C1(G329), .C2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G326), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n713), .A2(new_n269), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n721), .B(new_n735), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n731), .A2(new_n225), .ZN(new_n740));
  INV_X1    g0540(.A(new_n730), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n255), .B(new_n740), .C1(G97), .C2(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(G50), .A2(new_n737), .B1(new_n714), .B2(G68), .ZN(new_n743));
  INV_X1    g0543(.A(G159), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n733), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT32), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n718), .A2(new_n202), .B1(new_n725), .B2(new_n207), .ZN(new_n747));
  INV_X1    g0547(.A(new_n726), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n747), .B1(G77), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n742), .A2(new_n743), .A3(new_n746), .A4(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n711), .B1(new_n739), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n710), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n214), .A2(new_n540), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n704), .B2(new_n218), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(new_n246), .B2(new_n704), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n214), .A2(new_n256), .ZN(new_n760));
  INV_X1    g0560(.A(G355), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n761), .B1(G116), .B2(new_n214), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT90), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n756), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n751), .A2(new_n708), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n754), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n641), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n709), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(G396));
  INV_X1    g0569(.A(new_n708), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n317), .A2(new_n637), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n313), .B1(new_n312), .B2(new_n638), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n771), .B1(new_n772), .B2(new_n317), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n679), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n625), .A2(new_n638), .A3(new_n773), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n770), .B1(new_n777), .B2(new_n699), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n699), .B2(new_n777), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G143), .A2(new_n719), .B1(new_n748), .B2(G159), .ZN(new_n780));
  INV_X1    g0580(.A(new_n714), .ZN(new_n781));
  INV_X1    g0581(.A(G137), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n780), .B1(new_n781), .B2(new_n281), .C1(new_n782), .C2(new_n738), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT34), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n725), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G68), .ZN(new_n787));
  INV_X1    g0587(.A(G132), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n787), .B1(new_n201), .B2(new_n731), .C1(new_n788), .C2(new_n733), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n540), .B(new_n789), .C1(G58), .C2(new_n741), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n783), .A2(new_n784), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n785), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n255), .B1(new_n725), .B2(new_n225), .ZN(new_n793));
  INV_X1    g0593(.A(new_n496), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n794), .A2(new_n726), .B1(new_n731), .B2(new_n207), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n793), .B(new_n795), .C1(G311), .C2(new_n734), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n714), .A2(G283), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n718), .A2(new_n544), .B1(new_n730), .B2(new_n206), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT93), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n737), .A2(G303), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n792), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n711), .B1(new_n803), .B2(KEYINPUT94), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(KEYINPUT94), .B2(new_n803), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n710), .A2(new_n752), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n708), .B1(new_n223), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n805), .B(new_n807), .C1(new_n773), .C2(new_n753), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n779), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G384));
  AND3_X1   g0610(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT35), .ZN(new_n813));
  OAI211_X1 g0613(.A(G116), .B(new_n220), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT36), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n218), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n201), .A2(G68), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n210), .B(G13), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n407), .A2(new_n637), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT98), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n347), .A2(new_n273), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n338), .B1(new_n345), .B2(new_n346), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT95), .ZN(new_n826));
  OR2_X1    g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT16), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT96), .ZN(new_n830));
  INV_X1    g0630(.A(new_n363), .ZN(new_n831));
  OR3_X1    g0631(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n635), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n830), .B1(new_n829), .B2(new_n831), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n832), .A2(new_n336), .A3(new_n834), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n836), .A3(new_n371), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT37), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n365), .A2(new_n371), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n364), .A2(new_n833), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n839), .A2(KEYINPUT97), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n365), .A2(new_n841), .A3(new_n840), .A4(new_n371), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT97), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n838), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n835), .B1(new_n367), .B2(new_n372), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT39), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n845), .B2(new_n842), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n841), .B1(new_n367), .B2(new_n372), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n837), .A2(KEYINPUT37), .B1(new_n842), .B2(new_n845), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n852), .B1(new_n858), .B2(new_n848), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n851), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n823), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n771), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n776), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n850), .A2(new_n859), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n398), .A2(new_n638), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n408), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n401), .B(new_n407), .C1(new_n398), .C2(new_n638), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n863), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n367), .A2(new_n833), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n861), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n678), .A2(new_n409), .A3(new_n681), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n630), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n871), .B(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n868), .A2(new_n698), .A3(new_n773), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n864), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n850), .A2(new_n856), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(KEYINPUT40), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n409), .A2(new_n698), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(G330), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT99), .ZN(new_n887));
  OAI21_X1  g0687(.A(G1), .B1(new_n276), .B2(G20), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n887), .B(new_n888), .C1(new_n874), .C2(new_n885), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n886), .A2(KEYINPUT99), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n820), .B1(new_n889), .B2(new_n890), .ZN(G367));
  NAND3_X1  g0691(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT104), .Z(new_n893));
  NOR2_X1   g0693(.A1(new_n475), .A2(new_n638), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT101), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n470), .A2(new_n475), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n427), .A2(new_n637), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n650), .A2(new_n648), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT44), .Z(new_n901));
  NOR2_X1   g0701(.A1(new_n898), .A2(new_n899), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT45), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(new_n647), .Z(new_n905));
  OAI21_X1  g0705(.A(new_n650), .B1(new_n646), .B2(new_n649), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n906), .A2(new_n643), .A3(new_n642), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n703), .B2(new_n906), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n682), .A2(new_n699), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OR3_X1    g0710(.A1(new_n905), .A2(KEYINPUT103), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT103), .B1(new_n905), .B2(new_n910), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n700), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n652), .B(KEYINPUT41), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n893), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n487), .A2(new_n638), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT100), .Z(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n508), .A3(new_n507), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n619), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT102), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n898), .A2(new_n650), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT42), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n898), .A2(new_n570), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n472), .B2(new_n621), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n923), .B1(new_n637), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n921), .A3(new_n927), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n920), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n920), .A3(new_n930), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n647), .A2(new_n898), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n915), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n919), .A2(new_n766), .ZN(new_n938));
  INV_X1    g0738(.A(new_n241), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n755), .B1(new_n214), .B2(new_n308), .C1(new_n939), .C2(new_n757), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n770), .A2(new_n940), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n256), .B1(new_n730), .B2(new_n203), .C1(new_n223), .C2(new_n725), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n718), .A2(new_n281), .B1(new_n726), .B2(new_n201), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n731), .A2(new_n202), .B1(new_n733), .B2(new_n782), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n737), .A2(G143), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n945), .B(new_n946), .C1(new_n744), .C2(new_n781), .ZN(new_n947));
  INV_X1    g0747(.A(new_n731), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT46), .B1(new_n948), .B2(new_n496), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(G107), .B2(new_n741), .ZN(new_n950));
  XNOR2_X1  g0750(.A(KEYINPUT105), .B(G317), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n725), .A2(new_n206), .B1(new_n733), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(G283), .B2(new_n748), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n948), .A2(KEYINPUT46), .A3(G116), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G303), .B2(new_n719), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n950), .A2(new_n540), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n544), .A2(new_n781), .B1(new_n738), .B2(new_n727), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n947), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n941), .B1(new_n959), .B2(new_n710), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n938), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n937), .A2(new_n961), .ZN(G387));
  XOR2_X1   g0762(.A(new_n652), .B(KEYINPUT109), .Z(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n909), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n701), .B2(new_n908), .ZN(new_n966));
  INV_X1    g0766(.A(new_n893), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n646), .A2(new_n766), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n760), .A2(new_n655), .B1(G107), .B2(new_n214), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT106), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n238), .A2(G45), .ZN(new_n971));
  INV_X1    g0771(.A(new_n655), .ZN(new_n972));
  AOI211_X1 g0772(.A(G45), .B(new_n972), .C1(G68), .C2(G77), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n284), .A2(G50), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT50), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n757), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n970), .B1(new_n971), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n770), .B1(new_n977), .B2(new_n756), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n794), .A2(new_n725), .B1(new_n733), .B2(new_n736), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n737), .A2(G322), .ZN(new_n980));
  INV_X1    g0780(.A(new_n951), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n719), .A2(new_n981), .B1(new_n748), .B2(G303), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(new_n781), .C2(new_n727), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT48), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n948), .A2(G294), .B1(new_n741), .B2(G283), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT49), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n323), .B(new_n979), .C1(new_n990), .C2(KEYINPUT108), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(KEYINPUT108), .B2(new_n990), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n714), .A2(new_n361), .B1(G68), .B2(new_n748), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT107), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G50), .A2(new_n719), .B1(new_n734), .B2(G150), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n223), .B2(new_n731), .C1(new_n206), .C2(new_n725), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n540), .B(new_n996), .C1(new_n309), .C2(new_n741), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n744), .B2(new_n738), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n992), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n978), .B1(new_n999), .B2(new_n710), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n908), .A2(new_n967), .B1(new_n968), .B2(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n966), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT110), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(KEYINPUT110), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(G393));
  OAI221_X1 g0805(.A(new_n755), .B1(new_n206), .B2(new_n214), .C1(new_n249), .C2(new_n757), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G283), .A2(new_n948), .B1(new_n734), .B2(G322), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n544), .B2(new_n726), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n256), .B(new_n1008), .C1(G107), .C2(new_n786), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n781), .A2(new_n583), .B1(new_n794), .B2(new_n730), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(KEYINPUT111), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(KEYINPUT111), .B2(new_n1010), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n737), .A2(G317), .B1(G311), .B2(new_n719), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT52), .Z(new_n1014));
  AOI22_X1  g0814(.A1(new_n737), .A2(G150), .B1(G159), .B2(new_n719), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT51), .Z(new_n1016));
  AOI22_X1  g0816(.A1(G87), .A2(new_n786), .B1(new_n734), .B2(G143), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n203), .B2(new_n731), .C1(new_n284), .C2(new_n726), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n781), .A2(new_n201), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n730), .A2(new_n223), .ZN(new_n1020));
  NOR4_X1   g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n540), .A4(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1012), .A2(new_n1014), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n770), .B(new_n1006), .C1(new_n1022), .C2(new_n711), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n898), .B2(new_n754), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n904), .B(new_n647), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n967), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n964), .B1(new_n911), .B2(new_n912), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1025), .A2(new_n909), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT112), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  AND3_X1   g0830(.A1(new_n1027), .A2(KEYINPUT113), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT113), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1026), .B1(new_n1031), .B2(new_n1032), .ZN(G390));
  NAND2_X1  g0833(.A1(new_n676), .A2(new_n638), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n658), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n676), .A2(KEYINPUT87), .A3(new_n638), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n1036), .A3(new_n862), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n772), .A2(new_n317), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n868), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n879), .A2(new_n822), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n863), .A2(new_n868), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n822), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n857), .A2(new_n860), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n868), .A2(G330), .A3(new_n698), .A4(new_n773), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1042), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1047), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1049), .A2(new_n1050), .A3(new_n893), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1045), .A2(new_n752), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n806), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1053), .A2(new_n361), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(KEYINPUT54), .B(G143), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n256), .B1(new_n730), .B2(new_n744), .C1(new_n726), .C2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G132), .A2(new_n719), .B1(new_n734), .B2(G125), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n201), .B2(new_n725), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(G128), .C2(new_n737), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n731), .A2(new_n281), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT53), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT116), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1061), .A2(new_n1062), .B1(G137), .B2(new_n714), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1059), .B(new_n1063), .C1(new_n1062), .C2(new_n1061), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n714), .A2(G107), .B1(G97), .B2(new_n748), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n722), .B2(new_n738), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT117), .Z(new_n1067));
  OAI221_X1 g0867(.A(new_n787), .B1(new_n492), .B2(new_n718), .C1(new_n544), .C2(new_n733), .ZN(new_n1068));
  OR4_X1    g0868(.A1(new_n256), .A2(new_n1068), .A3(new_n740), .A4(new_n1020), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1064), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n708), .B(new_n1054), .C1(new_n1070), .C2(new_n710), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1051), .B1(new_n1052), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n698), .A2(G330), .A3(new_n773), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n867), .A3(new_n866), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n1047), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n774), .A2(KEYINPUT115), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1073), .B(new_n1078), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1076), .A2(KEYINPUT114), .A3(new_n863), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT114), .B1(new_n1076), .B2(new_n863), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n409), .A2(G330), .A3(new_n698), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n872), .A2(new_n630), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1047), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1038), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n673), .A2(new_n677), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n862), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1040), .B1(new_n1093), .B2(new_n868), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1090), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1089), .A2(new_n1096), .A3(new_n1048), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1088), .A2(new_n1097), .A3(new_n963), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1072), .A2(new_n1098), .ZN(G378));
  NOR2_X1   g0899(.A1(new_n323), .A2(G41), .ZN(new_n1100));
  AOI211_X1 g0900(.A(G50), .B(new_n1100), .C1(new_n253), .C2(new_n428), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n223), .A2(new_n731), .B1(new_n718), .B2(new_n207), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n309), .A2(new_n748), .B1(new_n786), .B2(G58), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n722), .B2(new_n733), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1102), .B(new_n1104), .C1(G68), .C2(new_n741), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G97), .A2(new_n714), .B1(new_n737), .B2(G116), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1100), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT58), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1101), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n726), .A2(new_n782), .ZN(new_n1110));
  INV_X1    g0910(.A(G128), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1111), .A2(new_n718), .B1(new_n731), .B2(new_n1055), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(G150), .C2(new_n741), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n737), .A2(G125), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(new_n788), .C2(new_n781), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1115), .A2(KEYINPUT59), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(KEYINPUT59), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n786), .A2(G159), .ZN(new_n1118));
  AOI211_X1 g0918(.A(G33), .B(G41), .C1(new_n734), .C2(G124), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1109), .B1(new_n1108), .B2(new_n1107), .C1(new_n1116), .C2(new_n1120), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1121), .A2(new_n710), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n770), .B1(G50), .B2(new_n1053), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n297), .B(KEYINPUT118), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n288), .A2(new_n635), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT119), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1124), .B(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1127), .B(new_n1128), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1122), .B(new_n1123), .C1(new_n1129), .C2(new_n752), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n878), .A2(G330), .A3(new_n880), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n871), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1135), .A2(KEYINPUT120), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1134), .B(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1130), .B1(new_n1137), .B2(new_n967), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1097), .A2(new_n1086), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT121), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT121), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1097), .A2(new_n1141), .A3(new_n1086), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT57), .B1(new_n1143), .B2(new_n1137), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT57), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1133), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n1135), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n871), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1097), .A2(new_n1141), .A3(new_n1086), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1141), .B1(new_n1097), .B2(new_n1086), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n963), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1138), .B1(new_n1144), .B2(new_n1154), .ZN(G375));
  AND2_X1   g0955(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1085), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n914), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n1087), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n770), .B1(G68), .B2(new_n1053), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n731), .A2(new_n744), .B1(new_n725), .B2(new_n202), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n540), .B(new_n1161), .C1(G50), .C2(new_n741), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G150), .A2(new_n748), .B1(new_n734), .B2(G128), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n782), .C2(new_n718), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n788), .A2(new_n738), .B1(new_n781), .B2(new_n1055), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n255), .B1(new_n730), .B2(new_n308), .C1(new_n223), .C2(new_n725), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n726), .A2(new_n207), .B1(new_n733), .B2(new_n583), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n206), .A2(new_n731), .B1(new_n718), .B2(new_n722), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n544), .B2(new_n738), .C1(new_n794), .C2(new_n781), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1166), .B1(KEYINPUT123), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(KEYINPUT123), .B2(new_n1171), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1160), .B1(new_n1173), .B2(new_n710), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n868), .B2(new_n753), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n893), .B(KEYINPUT122), .Z(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(new_n1156), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1159), .A2(new_n1178), .ZN(G381));
  AOI22_X1  g0979(.A1(new_n915), .A2(new_n936), .B1(new_n938), .B2(new_n960), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n1026), .C1(new_n1032), .C2(new_n1031), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1003), .A2(new_n768), .A3(new_n1004), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n1181), .A2(G384), .A3(G381), .A4(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT124), .B1(new_n1072), .B2(new_n1098), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1072), .A2(KEYINPUT124), .A3(new_n1098), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(G375), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(G407));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1183), .B2(new_n636), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(G213), .ZN(G409));
  OAI211_X1 g0989(.A(G378), .B(new_n1138), .C1(new_n1144), .C2(new_n1154), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1185), .A2(new_n1184), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1137), .B(new_n1158), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1176), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(new_n1130), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1190), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n636), .A2(G213), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1089), .A2(new_n964), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT125), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1157), .A2(new_n1201), .A3(KEYINPUT60), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT60), .B1(new_n1157), .B2(new_n1201), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1200), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1178), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n809), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(G384), .A3(new_n1178), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n636), .A2(G213), .A3(G2897), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT61), .B1(new_n1199), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1197), .A2(new_n1215), .A3(new_n1198), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT126), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT62), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1197), .A2(KEYINPUT62), .A3(new_n1215), .A4(new_n1198), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT126), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1190), .A2(new_n1196), .B1(G213), .B2(new_n636), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT62), .B1(new_n1222), .B2(new_n1215), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1213), .B(new_n1219), .C1(new_n1221), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G387), .A2(G390), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G393), .A2(G396), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1182), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1181), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1181), .B2(new_n1225), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1222), .A2(KEYINPUT63), .A3(new_n1215), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT63), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1216), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .A4(new_n1213), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1231), .A2(new_n1236), .ZN(G405));
  INV_X1    g1037(.A(new_n1190), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G375), .A2(new_n1191), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT127), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(G375), .A2(KEYINPUT127), .A3(new_n1191), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1214), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1241), .A2(new_n1214), .A3(new_n1242), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1230), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1243), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1241), .A2(new_n1214), .A3(new_n1242), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1232), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(G402));
endmodule


