

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(n726), .ZN(n744) );
  NOR2_X2 U551 ( .A1(n741), .A2(n740), .ZN(n752) );
  BUF_X1 U552 ( .A(n687), .Z(n577) );
  INV_X1 U553 ( .A(G2105), .ZN(n556) );
  NOR2_X2 U554 ( .A1(n707), .A2(n799), .ZN(n699) );
  NOR2_X1 U555 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U556 ( .A1(G651), .A2(n651), .ZN(n650) );
  NOR2_X1 U557 ( .A1(G651), .A2(G543), .ZN(n643) );
  XOR2_X1 U558 ( .A(KEYINPUT73), .B(n606), .Z(n519) );
  OR2_X1 U559 ( .A1(n834), .A2(n833), .ZN(n520) );
  NOR2_X1 U560 ( .A1(n764), .A2(n834), .ZN(n521) );
  NAND2_X1 U561 ( .A1(n831), .A2(n834), .ZN(n522) );
  OR2_X1 U562 ( .A1(n706), .A2(n988), .ZN(n705) );
  XNOR2_X1 U563 ( .A(n734), .B(KEYINPUT30), .ZN(n735) );
  NAND2_X1 U564 ( .A1(n695), .A2(n769), .ZN(n696) );
  INV_X1 U565 ( .A(KEYINPUT68), .ZN(n525) );
  XNOR2_X1 U566 ( .A(n525), .B(KEYINPUT1), .ZN(n526) );
  NOR2_X2 U567 ( .A1(G2104), .A2(n556), .ZN(n894) );
  AND2_X2 U568 ( .A1(n556), .A2(G2104), .ZN(n891) );
  XNOR2_X1 U569 ( .A(n614), .B(n613), .ZN(n988) );
  INV_X1 U570 ( .A(KEYINPUT66), .ZN(n562) );
  XNOR2_X1 U571 ( .A(n563), .B(n562), .ZN(n694) );
  XNOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n523), .B(KEYINPUT67), .ZN(n651) );
  NAND2_X1 U574 ( .A1(n650), .A2(G51), .ZN(n524) );
  XNOR2_X1 U575 ( .A(n524), .B(KEYINPUT78), .ZN(n529) );
  INV_X1 U576 ( .A(G651), .ZN(n533) );
  NOR2_X1 U577 ( .A1(G543), .A2(n533), .ZN(n527) );
  XNOR2_X2 U578 ( .A(n527), .B(n526), .ZN(n655) );
  NAND2_X1 U579 ( .A1(G63), .A2(n655), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U581 ( .A(KEYINPUT6), .B(n530), .ZN(n539) );
  NAND2_X1 U582 ( .A1(G89), .A2(n643), .ZN(n531) );
  XNOR2_X1 U583 ( .A(n531), .B(KEYINPUT4), .ZN(n532) );
  XNOR2_X1 U584 ( .A(n532), .B(KEYINPUT76), .ZN(n535) );
  NOR2_X1 U585 ( .A1(n651), .A2(n533), .ZN(n640) );
  NAND2_X1 U586 ( .A1(G76), .A2(n640), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U588 ( .A(KEYINPUT5), .B(n536), .ZN(n537) );
  XNOR2_X1 U589 ( .A(KEYINPUT77), .B(n537), .ZN(n538) );
  NOR2_X1 U590 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U591 ( .A(KEYINPUT7), .B(n540), .Z(G168) );
  NAND2_X1 U592 ( .A1(n643), .A2(G91), .ZN(n542) );
  NAND2_X1 U593 ( .A1(G65), .A2(n655), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U595 ( .A1(G78), .A2(n640), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G53), .A2(n650), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U598 ( .A1(n546), .A2(n545), .ZN(G299) );
  NAND2_X1 U599 ( .A1(G85), .A2(n643), .ZN(n548) );
  NAND2_X1 U600 ( .A1(G72), .A2(n640), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U602 ( .A1(n650), .A2(G47), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G60), .A2(n655), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  OR2_X1 U605 ( .A1(n552), .A2(n551), .ZN(G290) );
  NOR2_X1 U606 ( .A1(G2105), .A2(G2104), .ZN(n553) );
  XOR2_X1 U607 ( .A(KEYINPUT17), .B(n553), .Z(n687) );
  NAND2_X1 U608 ( .A1(n687), .A2(G137), .ZN(n561) );
  NAND2_X1 U609 ( .A1(G125), .A2(n894), .ZN(n555) );
  AND2_X1 U610 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  NAND2_X1 U611 ( .A1(G113), .A2(n895), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G101), .A2(n891), .ZN(n557) );
  XNOR2_X1 U614 ( .A(KEYINPUT23), .B(n557), .ZN(n558) );
  NOR2_X1 U615 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(n563) );
  BUF_X1 U617 ( .A(n694), .Z(G160) );
  XOR2_X1 U618 ( .A(G2446), .B(G2451), .Z(n565) );
  XNOR2_X1 U619 ( .A(G2454), .B(KEYINPUT107), .ZN(n564) );
  XNOR2_X1 U620 ( .A(n565), .B(n564), .ZN(n572) );
  XOR2_X1 U621 ( .A(G2438), .B(G2430), .Z(n567) );
  XNOR2_X1 U622 ( .A(G2435), .B(G2443), .ZN(n566) );
  XNOR2_X1 U623 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U624 ( .A(n568), .B(G2427), .Z(n570) );
  XNOR2_X1 U625 ( .A(G1348), .B(G1341), .ZN(n569) );
  XNOR2_X1 U626 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U627 ( .A(n572), .B(n571), .ZN(n573) );
  AND2_X1 U628 ( .A1(n573), .A2(G14), .ZN(G401) );
  NAND2_X1 U629 ( .A1(G123), .A2(n894), .ZN(n574) );
  XNOR2_X1 U630 ( .A(n574), .B(KEYINPUT18), .ZN(n582) );
  NAND2_X1 U631 ( .A1(G99), .A2(n891), .ZN(n576) );
  NAND2_X1 U632 ( .A1(G111), .A2(n895), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U634 ( .A1(G135), .A2(n577), .ZN(n578) );
  XNOR2_X1 U635 ( .A(KEYINPUT79), .B(n578), .ZN(n579) );
  NOR2_X1 U636 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U637 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U638 ( .A(KEYINPUT80), .B(n583), .ZN(n921) );
  XNOR2_X1 U639 ( .A(n921), .B(G2096), .ZN(n584) );
  OR2_X1 U640 ( .A1(G2100), .A2(n584), .ZN(G156) );
  INV_X1 U641 ( .A(G57), .ZN(G237) );
  INV_X1 U642 ( .A(G132), .ZN(G219) );
  INV_X1 U643 ( .A(G82), .ZN(G220) );
  NAND2_X1 U644 ( .A1(G94), .A2(G452), .ZN(n585) );
  XOR2_X1 U645 ( .A(KEYINPUT70), .B(n585), .Z(G173) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n586) );
  XNOR2_X1 U647 ( .A(n586), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U648 ( .A(G223), .B(KEYINPUT71), .ZN(n841) );
  NAND2_X1 U649 ( .A1(n841), .A2(G567), .ZN(n587) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n587), .Z(G234) );
  XOR2_X1 U651 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n589) );
  NAND2_X1 U652 ( .A1(G56), .A2(n655), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n595) );
  NAND2_X1 U654 ( .A1(n643), .A2(G81), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(KEYINPUT12), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G68), .A2(n640), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U658 ( .A(KEYINPUT13), .B(n593), .Z(n594) );
  NOR2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U660 ( .A1(n650), .A2(G43), .ZN(n596) );
  NAND2_X1 U661 ( .A1(n597), .A2(n596), .ZN(n978) );
  INV_X1 U662 ( .A(G860), .ZN(n619) );
  OR2_X1 U663 ( .A1(n978), .A2(n619), .ZN(G153) );
  NAND2_X1 U664 ( .A1(n640), .A2(G77), .ZN(n598) );
  XOR2_X1 U665 ( .A(KEYINPUT69), .B(n598), .Z(n600) );
  NAND2_X1 U666 ( .A1(n643), .A2(G90), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U668 ( .A(KEYINPUT9), .B(n601), .ZN(n605) );
  NAND2_X1 U669 ( .A1(n655), .A2(G64), .ZN(n603) );
  NAND2_X1 U670 ( .A1(n650), .A2(G52), .ZN(n602) );
  AND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(G301) );
  NAND2_X1 U673 ( .A1(G868), .A2(G301), .ZN(n616) );
  NAND2_X1 U674 ( .A1(G66), .A2(n655), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n643), .A2(G92), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n519), .A2(n607), .ZN(n608) );
  XNOR2_X1 U677 ( .A(KEYINPUT74), .B(n608), .ZN(n612) );
  NAND2_X1 U678 ( .A1(G79), .A2(n640), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G54), .A2(n650), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n614) );
  XNOR2_X1 U682 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n613) );
  OR2_X1 U683 ( .A1(n988), .A2(G868), .ZN(n615) );
  NAND2_X1 U684 ( .A1(n616), .A2(n615), .ZN(G284) );
  XOR2_X1 U685 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U686 ( .A(G868), .ZN(n667) );
  NOR2_X1 U687 ( .A1(G286), .A2(n667), .ZN(n618) );
  NOR2_X1 U688 ( .A1(G868), .A2(G299), .ZN(n617) );
  NOR2_X1 U689 ( .A1(n618), .A2(n617), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n619), .A2(G559), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n620), .A2(n988), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n621), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(G868), .A2(n978), .ZN(n624) );
  NAND2_X1 U694 ( .A1(G868), .A2(n988), .ZN(n622) );
  NOR2_X1 U695 ( .A1(G559), .A2(n622), .ZN(n623) );
  NOR2_X1 U696 ( .A1(n624), .A2(n623), .ZN(G282) );
  NAND2_X1 U697 ( .A1(n988), .A2(G559), .ZN(n665) );
  XNOR2_X1 U698 ( .A(n978), .B(n665), .ZN(n625) );
  NOR2_X1 U699 ( .A1(n625), .A2(G860), .ZN(n632) );
  NAND2_X1 U700 ( .A1(n643), .A2(G93), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G67), .A2(n655), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U703 ( .A1(G80), .A2(n640), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G55), .A2(n650), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n630) );
  OR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n668) );
  XOR2_X1 U707 ( .A(n632), .B(n668), .Z(G145) );
  NAND2_X1 U708 ( .A1(n650), .A2(G50), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G62), .A2(n655), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U711 ( .A(KEYINPUT83), .B(n635), .ZN(n639) );
  NAND2_X1 U712 ( .A1(G88), .A2(n643), .ZN(n637) );
  NAND2_X1 U713 ( .A1(G75), .A2(n640), .ZN(n636) );
  AND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(G303) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n642) );
  NAND2_X1 U717 ( .A1(G73), .A2(n640), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n642), .B(n641), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n643), .A2(G86), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G61), .A2(n655), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n650), .A2(G48), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(G305) );
  NAND2_X1 U725 ( .A1(n650), .A2(G49), .ZN(n657) );
  NAND2_X1 U726 ( .A1(G87), .A2(n651), .ZN(n653) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U731 ( .A(KEYINPUT81), .B(n658), .Z(G288) );
  XNOR2_X1 U732 ( .A(KEYINPUT19), .B(n668), .ZN(n659) );
  XNOR2_X1 U733 ( .A(G299), .B(n659), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(G290), .ZN(n663) );
  XNOR2_X1 U735 ( .A(G303), .B(G305), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(G288), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n664), .B(n978), .ZN(n868) );
  XOR2_X1 U739 ( .A(n868), .B(n665), .Z(n666) );
  NAND2_X1 U740 ( .A1(G868), .A2(n666), .ZN(n670) );
  NAND2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n670), .A2(n669), .ZN(G295) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n672) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n672), .B(n671), .ZN(n673) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U748 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n676) );
  XNOR2_X1 U751 ( .A(KEYINPUT22), .B(n676), .ZN(n677) );
  NAND2_X1 U752 ( .A1(n677), .A2(G96), .ZN(n678) );
  NOR2_X1 U753 ( .A1(n678), .A2(G218), .ZN(n679) );
  XNOR2_X1 U754 ( .A(n679), .B(KEYINPUT85), .ZN(n847) );
  NAND2_X1 U755 ( .A1(G2106), .A2(n847), .ZN(n683) );
  NAND2_X1 U756 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U757 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U758 ( .A1(G108), .A2(n681), .ZN(n846) );
  NAND2_X1 U759 ( .A1(G567), .A2(n846), .ZN(n682) );
  NAND2_X1 U760 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U761 ( .A(KEYINPUT86), .B(n684), .Z(G319) );
  INV_X1 U762 ( .A(G319), .ZN(n686) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n685) );
  NOR2_X1 U764 ( .A1(n686), .A2(n685), .ZN(n845) );
  NAND2_X1 U765 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U766 ( .A1(G102), .A2(n891), .ZN(n689) );
  NAND2_X1 U767 ( .A1(G138), .A2(n687), .ZN(n688) );
  NAND2_X1 U768 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U769 ( .A1(G126), .A2(n894), .ZN(n691) );
  NAND2_X1 U770 ( .A1(G114), .A2(n895), .ZN(n690) );
  NAND2_X1 U771 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U772 ( .A1(n693), .A2(n692), .ZN(G164) );
  INV_X1 U773 ( .A(G303), .ZN(G166) );
  NAND2_X1 U774 ( .A1(n694), .A2(G40), .ZN(n768) );
  INV_X1 U775 ( .A(n768), .ZN(n695) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n769) );
  XNOR2_X2 U777 ( .A(n696), .B(KEYINPUT64), .ZN(n707) );
  NAND2_X1 U778 ( .A1(n707), .A2(G8), .ZN(n834) );
  NOR2_X1 U779 ( .A1(G1976), .A2(G288), .ZN(n975) );
  NAND2_X1 U780 ( .A1(n975), .A2(KEYINPUT33), .ZN(n697) );
  OR2_X1 U781 ( .A1(n834), .A2(n697), .ZN(n809) );
  INV_X1 U782 ( .A(G1996), .ZN(n799) );
  XNOR2_X1 U783 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n698) );
  XNOR2_X1 U784 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U785 ( .A1(n707), .A2(G1341), .ZN(n700) );
  NAND2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n703) );
  INV_X1 U787 ( .A(KEYINPUT95), .ZN(n702) );
  XNOR2_X1 U788 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U789 ( .A1(n704), .A2(n978), .ZN(n706) );
  XNOR2_X1 U790 ( .A(n705), .B(KEYINPUT96), .ZN(n713) );
  NAND2_X1 U791 ( .A1(n706), .A2(n988), .ZN(n711) );
  INV_X1 U792 ( .A(n707), .ZN(n726) );
  NOR2_X1 U793 ( .A1(G2067), .A2(n744), .ZN(n709) );
  NOR2_X1 U794 ( .A1(G1348), .A2(n726), .ZN(n708) );
  NOR2_X1 U795 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U797 ( .A1(n713), .A2(n712), .ZN(n719) );
  NAND2_X1 U798 ( .A1(G2072), .A2(n726), .ZN(n714) );
  XOR2_X1 U799 ( .A(KEYINPUT27), .B(n714), .Z(n716) );
  NAND2_X1 U800 ( .A1(n744), .A2(G1956), .ZN(n715) );
  NAND2_X1 U801 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U802 ( .A1(G299), .A2(n720), .ZN(n717) );
  XNOR2_X1 U803 ( .A(n717), .B(KEYINPUT97), .ZN(n718) );
  NAND2_X1 U804 ( .A1(n719), .A2(n718), .ZN(n724) );
  NAND2_X1 U805 ( .A1(n720), .A2(G299), .ZN(n721) );
  XNOR2_X1 U806 ( .A(n721), .B(KEYINPUT28), .ZN(n722) );
  XNOR2_X1 U807 ( .A(KEYINPUT94), .B(n722), .ZN(n723) );
  NAND2_X1 U808 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U809 ( .A(n725), .B(KEYINPUT29), .ZN(n731) );
  XOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .Z(n958) );
  NAND2_X1 U811 ( .A1(n958), .A2(n726), .ZN(n728) );
  NAND2_X1 U812 ( .A1(n744), .A2(G1961), .ZN(n727) );
  NAND2_X1 U813 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U814 ( .A1(G301), .A2(n732), .ZN(n729) );
  XOR2_X1 U815 ( .A(KEYINPUT93), .B(n729), .Z(n730) );
  NOR2_X1 U816 ( .A1(n731), .A2(n730), .ZN(n741) );
  AND2_X1 U817 ( .A1(G301), .A2(n732), .ZN(n737) );
  NOR2_X1 U818 ( .A1(G1966), .A2(n834), .ZN(n753) );
  NOR2_X1 U819 ( .A1(n744), .A2(G2084), .ZN(n754) );
  NOR2_X1 U820 ( .A1(n753), .A2(n754), .ZN(n733) );
  NAND2_X1 U821 ( .A1(G8), .A2(n733), .ZN(n734) );
  NOR2_X1 U822 ( .A1(n735), .A2(G168), .ZN(n736) );
  NOR2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U824 ( .A(KEYINPUT98), .B(n738), .ZN(n739) );
  XNOR2_X1 U825 ( .A(KEYINPUT31), .B(n739), .ZN(n740) );
  INV_X1 U826 ( .A(n752), .ZN(n742) );
  NAND2_X1 U827 ( .A1(n742), .A2(G286), .ZN(n743) );
  XNOR2_X1 U828 ( .A(n743), .B(KEYINPUT100), .ZN(n749) );
  NOR2_X1 U829 ( .A1(n744), .A2(G2090), .ZN(n746) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n834), .ZN(n745) );
  NOR2_X1 U831 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n747), .A2(G303), .ZN(n748) );
  NAND2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U834 ( .A1(n750), .A2(G8), .ZN(n751) );
  XNOR2_X1 U835 ( .A(n751), .B(KEYINPUT32), .ZN(n826) );
  NOR2_X1 U836 ( .A1(n753), .A2(n752), .ZN(n756) );
  NAND2_X1 U837 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U838 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U839 ( .A(KEYINPUT99), .B(n757), .Z(n825) );
  NAND2_X1 U840 ( .A1(n826), .A2(n825), .ZN(n762) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U842 ( .A1(n975), .A2(n758), .ZN(n760) );
  INV_X1 U843 ( .A(KEYINPUT33), .ZN(n759) );
  AND2_X1 U844 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U845 ( .A1(n762), .A2(n761), .ZN(n766) );
  NAND2_X1 U846 ( .A1(G288), .A2(G1976), .ZN(n763) );
  XOR2_X1 U847 ( .A(KEYINPUT101), .B(n763), .Z(n981) );
  INV_X1 U848 ( .A(n981), .ZN(n764) );
  OR2_X1 U849 ( .A1(KEYINPUT33), .A2(n521), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U851 ( .A(n767), .B(KEYINPUT102), .ZN(n807) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n970) );
  XNOR2_X1 U853 ( .A(G1986), .B(G290), .ZN(n974) );
  NOR2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n821) );
  AND2_X1 U855 ( .A1(n974), .A2(n821), .ZN(n805) );
  XNOR2_X1 U856 ( .A(KEYINPUT37), .B(G2067), .ZN(n817) );
  NAND2_X1 U857 ( .A1(n891), .A2(G104), .ZN(n770) );
  XOR2_X1 U858 ( .A(KEYINPUT87), .B(n770), .Z(n772) );
  NAND2_X1 U859 ( .A1(n577), .A2(G140), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U861 ( .A(KEYINPUT34), .B(n773), .ZN(n779) );
  NAND2_X1 U862 ( .A1(n894), .A2(G128), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n774), .B(KEYINPUT88), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G116), .A2(n895), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U866 ( .A(KEYINPUT35), .B(n777), .Z(n778) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U868 ( .A(KEYINPUT36), .B(n780), .ZN(n912) );
  NOR2_X1 U869 ( .A1(n817), .A2(n912), .ZN(n936) );
  NAND2_X1 U870 ( .A1(n821), .A2(n936), .ZN(n815) );
  NAND2_X1 U871 ( .A1(G95), .A2(n891), .ZN(n781) );
  XOR2_X1 U872 ( .A(KEYINPUT90), .B(n781), .Z(n786) );
  NAND2_X1 U873 ( .A1(G119), .A2(n894), .ZN(n783) );
  NAND2_X1 U874 ( .A1(G107), .A2(n895), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U876 ( .A(KEYINPUT89), .B(n784), .Z(n785) );
  NOR2_X1 U877 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n577), .A2(G131), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n909) );
  NAND2_X1 U880 ( .A1(G1991), .A2(n909), .ZN(n789) );
  XNOR2_X1 U881 ( .A(n789), .B(KEYINPUT91), .ZN(n801) );
  NAND2_X1 U882 ( .A1(G117), .A2(n895), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G141), .A2(n577), .ZN(n791) );
  NAND2_X1 U884 ( .A1(G129), .A2(n894), .ZN(n790) );
  NAND2_X1 U885 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n891), .A2(G105), .ZN(n792) );
  XOR2_X1 U887 ( .A(KEYINPUT38), .B(n792), .Z(n793) );
  NOR2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U890 ( .A(n797), .B(KEYINPUT92), .ZN(n904) );
  INV_X1 U891 ( .A(n904), .ZN(n798) );
  NOR2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n926) );
  INV_X1 U894 ( .A(n821), .ZN(n802) );
  NOR2_X1 U895 ( .A1(n926), .A2(n802), .ZN(n812) );
  INV_X1 U896 ( .A(n812), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n815), .A2(n803), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n835) );
  NAND2_X1 U899 ( .A1(n970), .A2(n835), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n824) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n904), .ZN(n928) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n909), .ZN(n924) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n924), .A2(n810), .ZN(n811) );
  NOR2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U906 ( .A1(n928), .A2(n813), .ZN(n814) );
  XNOR2_X1 U907 ( .A(KEYINPUT39), .B(n814), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n912), .A2(n817), .ZN(n818) );
  XNOR2_X1 U910 ( .A(n818), .B(KEYINPUT104), .ZN(n942) );
  NAND2_X1 U911 ( .A1(n819), .A2(n942), .ZN(n820) );
  XOR2_X1 U912 ( .A(KEYINPUT105), .B(n820), .Z(n822) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U914 ( .A1(n824), .A2(n823), .ZN(n838) );
  AND2_X1 U915 ( .A1(n826), .A2(n825), .ZN(n829) );
  NAND2_X1 U916 ( .A1(G166), .A2(G8), .ZN(n827) );
  NOR2_X1 U917 ( .A1(G2090), .A2(n827), .ZN(n828) );
  NOR2_X1 U918 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U919 ( .A(n830), .B(KEYINPUT103), .ZN(n831) );
  NOR2_X1 U920 ( .A1(G1981), .A2(G305), .ZN(n832) );
  XOR2_X1 U921 ( .A(n832), .B(KEYINPUT24), .Z(n833) );
  NAND2_X1 U922 ( .A1(n522), .A2(n520), .ZN(n836) );
  NAND2_X1 U923 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U924 ( .A1(n838), .A2(n837), .ZN(n840) );
  XNOR2_X1 U925 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n839) );
  XNOR2_X1 U926 ( .A(n840), .B(n839), .ZN(G329) );
  NAND2_X1 U927 ( .A1(n841), .A2(G2106), .ZN(n842) );
  XNOR2_X1 U928 ( .A(n842), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U930 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U932 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XOR2_X1 U939 ( .A(G1976), .B(G1971), .Z(n849) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1956), .ZN(n848) );
  XNOR2_X1 U941 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U942 ( .A(n850), .B(G2474), .Z(n852) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U944 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U945 ( .A(KEYINPUT41), .B(G1981), .Z(n854) );
  XNOR2_X1 U946 ( .A(G1966), .B(G1961), .ZN(n853) );
  XNOR2_X1 U947 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U948 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U949 ( .A(KEYINPUT109), .B(G2072), .Z(n858) );
  XNOR2_X1 U950 ( .A(G2084), .B(G2078), .ZN(n857) );
  XNOR2_X1 U951 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U952 ( .A(n859), .B(G2100), .Z(n861) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2090), .ZN(n860) );
  XNOR2_X1 U954 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U955 ( .A(G2096), .B(KEYINPUT43), .Z(n863) );
  XNOR2_X1 U956 ( .A(G2678), .B(KEYINPUT42), .ZN(n862) );
  XNOR2_X1 U957 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U958 ( .A(n865), .B(n864), .Z(G227) );
  INV_X1 U959 ( .A(G301), .ZN(G171) );
  XOR2_X1 U960 ( .A(KEYINPUT115), .B(G286), .Z(n867) );
  XNOR2_X1 U961 ( .A(G171), .B(n988), .ZN(n866) );
  XNOR2_X1 U962 ( .A(n867), .B(n866), .ZN(n869) );
  XNOR2_X1 U963 ( .A(n869), .B(n868), .ZN(n870) );
  NOR2_X1 U964 ( .A1(G37), .A2(n870), .ZN(n871) );
  XNOR2_X1 U965 ( .A(KEYINPUT116), .B(n871), .ZN(G397) );
  NAND2_X1 U966 ( .A1(G112), .A2(n895), .ZN(n872) );
  XNOR2_X1 U967 ( .A(n872), .B(KEYINPUT110), .ZN(n875) );
  NAND2_X1 U968 ( .A1(G124), .A2(n894), .ZN(n873) );
  XNOR2_X1 U969 ( .A(n873), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U970 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U971 ( .A1(G100), .A2(n891), .ZN(n877) );
  NAND2_X1 U972 ( .A1(G136), .A2(n577), .ZN(n876) );
  NAND2_X1 U973 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U974 ( .A1(n879), .A2(n878), .ZN(G162) );
  NAND2_X1 U975 ( .A1(G106), .A2(n891), .ZN(n881) );
  NAND2_X1 U976 ( .A1(G142), .A2(n577), .ZN(n880) );
  NAND2_X1 U977 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U978 ( .A(n882), .B(KEYINPUT45), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G130), .A2(n894), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G118), .A2(n895), .ZN(n885) );
  XNOR2_X1 U982 ( .A(KEYINPUT111), .B(n885), .ZN(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n908) );
  XOR2_X1 U984 ( .A(KEYINPUT113), .B(KEYINPUT48), .Z(n889) );
  XNOR2_X1 U985 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U987 ( .A(n890), .B(KEYINPUT112), .Z(n902) );
  NAND2_X1 U988 ( .A1(G103), .A2(n891), .ZN(n893) );
  NAND2_X1 U989 ( .A1(G139), .A2(n577), .ZN(n892) );
  NAND2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U991 ( .A1(G127), .A2(n894), .ZN(n897) );
  NAND2_X1 U992 ( .A1(G115), .A2(n895), .ZN(n896) );
  NAND2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U995 ( .A1(n900), .A2(n899), .ZN(n931) );
  XNOR2_X1 U996 ( .A(G164), .B(n931), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n921), .B(n903), .ZN(n906) );
  XNOR2_X1 U999 ( .A(G160), .B(n904), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n911) );
  XNOR2_X1 U1002 ( .A(n909), .B(G162), .ZN(n910) );
  XNOR2_X1 U1003 ( .A(n911), .B(n910), .ZN(n913) );
  XNOR2_X1 U1004 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n914), .ZN(G395) );
  NOR2_X1 U1006 ( .A1(G229), .A2(G227), .ZN(n915) );
  XOR2_X1 U1007 ( .A(KEYINPUT49), .B(n915), .Z(n916) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n916), .ZN(n917) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n917), .ZN(n920) );
  NOR2_X1 U1010 ( .A1(G397), .A2(G395), .ZN(n918) );
  XOR2_X1 U1011 ( .A(KEYINPUT117), .B(n918), .Z(n919) );
  NAND2_X1 U1012 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(KEYINPUT55), .ZN(n945) );
  XNOR2_X1 U1016 ( .A(G2084), .B(G160), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1019 ( .A1(n926), .A2(n925), .ZN(n940) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1021 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1022 ( .A(KEYINPUT118), .B(n929), .Z(n930) );
  XNOR2_X1 U1023 ( .A(KEYINPUT51), .B(n930), .ZN(n938) );
  XOR2_X1 U1024 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n934), .Z(n935) );
  NOR2_X1 U1028 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1030 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1031 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1032 ( .A(KEYINPUT52), .B(n943), .Z(n944) );
  NAND2_X1 U1033 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1034 ( .A1(n946), .A2(G29), .ZN(n998) );
  XNOR2_X1 U1035 ( .A(G2084), .B(G34), .ZN(n947) );
  XNOR2_X1 U1036 ( .A(n947), .B(KEYINPUT54), .ZN(n949) );
  XNOR2_X1 U1037 ( .A(G35), .B(G2090), .ZN(n948) );
  NOR2_X1 U1038 ( .A1(n949), .A2(n948), .ZN(n964) );
  XNOR2_X1 U1039 ( .A(G2067), .B(G26), .ZN(n951) );
  XNOR2_X1 U1040 ( .A(G32), .B(G1996), .ZN(n950) );
  NOR2_X1 U1041 ( .A1(n951), .A2(n950), .ZN(n957) );
  XOR2_X1 U1042 ( .A(G2072), .B(G33), .Z(n952) );
  NAND2_X1 U1043 ( .A1(n952), .A2(G28), .ZN(n955) );
  XOR2_X1 U1044 ( .A(G25), .B(G1991), .Z(n953) );
  XNOR2_X1 U1045 ( .A(KEYINPUT119), .B(n953), .ZN(n954) );
  NOR2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1047 ( .A1(n957), .A2(n956), .ZN(n960) );
  XNOR2_X1 U1048 ( .A(G27), .B(n958), .ZN(n959) );
  NOR2_X1 U1049 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1050 ( .A(n961), .B(KEYINPUT120), .Z(n962) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n962), .ZN(n963) );
  NAND2_X1 U1052 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1053 ( .A(KEYINPUT55), .B(n965), .ZN(n966) );
  NOR2_X1 U1054 ( .A1(G29), .A2(n966), .ZN(n967) );
  XNOR2_X1 U1055 ( .A(n967), .B(KEYINPUT121), .ZN(n968) );
  NAND2_X1 U1056 ( .A1(G11), .A2(n968), .ZN(n996) );
  XOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .Z(n994) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(n969), .B(KEYINPUT122), .ZN(n971) );
  NAND2_X1 U1060 ( .A1(n971), .A2(n970), .ZN(n973) );
  XOR2_X1 U1061 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n972) );
  XNOR2_X1 U1062 ( .A(n973), .B(n972), .ZN(n987) );
  NOR2_X1 U1063 ( .A1(n975), .A2(n974), .ZN(n977) );
  XOR2_X1 U1064 ( .A(G1956), .B(G299), .Z(n976) );
  NAND2_X1 U1065 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1066 ( .A(G1341), .B(n978), .ZN(n979) );
  NOR2_X1 U1067 ( .A1(n980), .A2(n979), .ZN(n982) );
  NAND2_X1 U1068 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1069 ( .A(G1971), .B(G166), .Z(n983) );
  XNOR2_X1 U1070 ( .A(KEYINPUT124), .B(n983), .ZN(n984) );
  NOR2_X1 U1071 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1072 ( .A1(n987), .A2(n986), .ZN(n992) );
  XNOR2_X1 U1073 ( .A(G1348), .B(n988), .ZN(n990) );
  XNOR2_X1 U1074 ( .A(G171), .B(G1961), .ZN(n989) );
  NAND2_X1 U1075 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1076 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1077 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1078 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1079 ( .A1(n998), .A2(n997), .ZN(n1024) );
  XOR2_X1 U1080 ( .A(KEYINPUT125), .B(G16), .Z(n1022) );
  XOR2_X1 U1081 ( .A(G1961), .B(G5), .Z(n1008) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .ZN(n999) );
  XNOR2_X1 U1083 ( .A(n999), .B(G4), .ZN(n1003) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n1000) );
  NOR2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1088 ( .A(G20), .B(G1956), .ZN(n1004) );
  NOR2_X1 U1089 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1091 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  XNOR2_X1 U1092 ( .A(G21), .B(G1966), .ZN(n1009) );
  NOR2_X1 U1093 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(KEYINPUT126), .B(n1011), .Z(n1019) );
  XOR2_X1 U1095 ( .A(G1976), .B(G23), .Z(n1014) );
  XNOR2_X1 U1096 ( .A(G1986), .B(KEYINPUT127), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(n1012), .B(G24), .ZN(n1013) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(G22), .B(G1971), .ZN(n1015) );
  NOR2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1017), .Z(n1018) );
  NOR2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1020), .Z(n1021) );
  NOR2_X1 U1104 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1105 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1106 ( .A(n1025), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

