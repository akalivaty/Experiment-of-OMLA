//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  OAI21_X1  g0007(.A(G50), .B1(G58), .B2(G68), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(G20), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT65), .B(G77), .Z(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT67), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n213), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n216), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(G33), .A2(G87), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT68), .B(G1698), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n249), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI211_X1 g0055(.A(KEYINPUT81), .B(new_n248), .C1(new_n250), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT81), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G1698), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n261), .A3(G223), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G226), .A2(G1698), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n255), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n248), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n257), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n256), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n267), .A2(new_n273), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n274), .B1(new_n276), .B2(new_n233), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n268), .A2(G179), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n267), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n248), .B1(new_n250), .B2(new_n255), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(new_n257), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n277), .B1(new_n282), .B2(new_n256), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n279), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT18), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT70), .ZN(new_n287));
  INV_X1    g0087(.A(G58), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT69), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT8), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n288), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT69), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n289), .A2(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(new_n210), .ZN(new_n297));
  INV_X1    g0097(.A(G20), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(G1), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G13), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(G1), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G20), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n291), .A2(new_n294), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(KEYINPUT3), .B(G33), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT7), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n306), .A2(new_n307), .A3(G20), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT7), .B1(new_n255), .B2(new_n298), .ZN(new_n309));
  OAI21_X1  g0109(.A(G68), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n288), .A2(new_n219), .ZN(new_n311));
  NOR2_X1   g0111(.A1(G58), .A2(G68), .ZN(new_n312));
  OAI21_X1  g0112(.A(G20), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(G20), .A2(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G159), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n310), .A2(KEYINPUT16), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n297), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n307), .A2(G20), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT80), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n254), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n252), .A2(KEYINPUT80), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n307), .B1(new_n306), .B2(G20), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G68), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n322), .B1(new_n330), .B2(new_n317), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n305), .B1(new_n320), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n285), .A2(new_n286), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n286), .B1(new_n285), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT15), .B(G87), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT72), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n253), .A2(G20), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n220), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT8), .B(G58), .Z(new_n342));
  AOI22_X1  g0142(.A1(new_n341), .A2(G20), .B1(new_n314), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n297), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n299), .A2(new_n202), .B1(new_n341), .B2(new_n303), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n259), .A2(new_n261), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n306), .B1(new_n218), .B2(new_n258), .C1(new_n233), .C2(new_n347), .ZN(new_n348));
  OR2_X1    g0148(.A1(KEYINPUT71), .A2(G107), .ZN(new_n349));
  NAND2_X1  g0149(.A1(KEYINPUT71), .A2(G107), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n348), .B(new_n267), .C1(new_n306), .C2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n273), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n353), .A2(new_n267), .A3(new_n269), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(G244), .B2(new_n275), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n346), .B1(new_n358), .B2(KEYINPUT73), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT73), .B1(new_n356), .B2(G169), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n357), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n306), .A2(G223), .A3(G1698), .ZN(new_n364));
  INV_X1    g0164(.A(G222), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n252), .A2(new_n254), .A3(new_n259), .A4(new_n261), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n364), .B1(new_n220), .B2(new_n306), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n267), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n354), .B1(G226), .B2(new_n275), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n284), .ZN(new_n371));
  MUX2_X1   g0171(.A(new_n303), .B(new_n299), .S(G50), .Z(new_n372));
  INV_X1    g0172(.A(G150), .ZN(new_n373));
  INV_X1    g0173(.A(new_n314), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(new_n201), .B2(new_n298), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n295), .B2(new_n339), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n372), .B1(new_n376), .B2(new_n297), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n371), .B(new_n377), .C1(G179), .C2(new_n370), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n356), .A2(G190), .ZN(new_n379));
  INV_X1    g0179(.A(G200), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n379), .B(new_n346), .C1(new_n380), .C2(new_n356), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n363), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n298), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n328), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n316), .B1(new_n384), .B2(G68), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n297), .B1(new_n385), .B2(KEYINPUT16), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n219), .B1(new_n327), .B2(new_n328), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n321), .B1(new_n387), .B2(new_n316), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G190), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n268), .A2(new_n390), .A3(new_n278), .ZN(new_n391));
  AOI21_X1  g0191(.A(G200), .B1(new_n268), .B2(new_n278), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n389), .B(new_n305), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  XOR2_X1   g0193(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n268), .A2(new_n390), .A3(new_n278), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n283), .B2(G200), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n386), .A2(new_n388), .B1(new_n304), .B2(new_n300), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT82), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n398), .B(new_n399), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n377), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT9), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n368), .A2(G190), .A3(new_n369), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT9), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n377), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n370), .A2(G200), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n405), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n410), .A2(KEYINPUT10), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(KEYINPUT10), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND4_X1   g0213(.A1(new_n335), .A2(new_n382), .A3(new_n403), .A4(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G238), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n274), .B1(new_n276), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n259), .A2(new_n261), .A3(G226), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G232), .A2(G1698), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n255), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n253), .A2(new_n204), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n267), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(KEYINPUT74), .B(new_n267), .C1(new_n419), .C2(new_n420), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n416), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XOR2_X1   g0225(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n426), .ZN(new_n428));
  AOI211_X1 g0228(.A(new_n428), .B(new_n416), .C1(new_n423), .C2(new_n424), .ZN(new_n429));
  OAI21_X1  g0229(.A(G169), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT14), .ZN(new_n431));
  INV_X1    g0231(.A(new_n429), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n425), .A2(KEYINPUT76), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT13), .B1(new_n425), .B2(KEYINPUT76), .ZN(new_n434));
  OAI211_X1 g0234(.A(G179), .B(new_n432), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n436), .B(G169), .C1(new_n427), .C2(new_n429), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT78), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n431), .A2(new_n435), .A3(KEYINPUT78), .A4(new_n437), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT12), .ZN(new_n443));
  INV_X1    g0243(.A(new_n303), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(new_n219), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n303), .A2(KEYINPUT12), .A3(G68), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n445), .A2(new_n446), .B1(new_n219), .B2(new_n299), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n314), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n298), .A2(G33), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(new_n202), .B2(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n450), .A2(KEYINPUT11), .A3(new_n319), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT11), .B1(new_n450), .B2(new_n319), .ZN(new_n452));
  OR3_X1    g0252(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n442), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n425), .B(new_n426), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n455), .B2(G200), .ZN(new_n456));
  OAI211_X1 g0256(.A(G190), .B(new_n432), .C1(new_n433), .C2(new_n434), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n456), .A2(KEYINPUT77), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT77), .B1(new_n456), .B2(new_n457), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n414), .A2(new_n454), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT4), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n252), .A2(new_n254), .A3(G244), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(new_n347), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n306), .A2(new_n249), .A3(KEYINPUT4), .A4(G244), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n306), .A2(G250), .A3(G1698), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n267), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT84), .B1(new_n472), .B2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT84), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(new_n271), .A3(KEYINPUT5), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G1), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n477), .B(G45), .C1(new_n271), .C2(KEYINPUT5), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n267), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n473), .B2(new_n475), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n480), .A2(G257), .B1(new_n270), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n471), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT85), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT85), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n471), .A2(new_n485), .A3(new_n482), .ZN(new_n486));
  AOI21_X1  g0286(.A(G169), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G97), .A2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n206), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT6), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n491), .A2(KEYINPUT83), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n491), .A2(KEYINPUT83), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n492), .A2(new_n493), .B1(new_n204), .B2(G107), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n495), .A2(new_n298), .B1(new_n202), .B2(new_n374), .ZN(new_n496));
  INV_X1    g0296(.A(new_n351), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n327), .B2(new_n328), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n319), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n303), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n477), .A2(G33), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n297), .A2(new_n303), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n502), .B2(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(G179), .B2(new_n483), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT86), .B1(new_n487), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n471), .A2(new_n485), .A3(new_n482), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n485), .B1(new_n471), .B2(new_n482), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G190), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n504), .B1(G200), .B2(new_n483), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n284), .B1(new_n507), .B2(new_n508), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT86), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n476), .A2(new_n479), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(G257), .A3(new_n280), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n481), .A2(new_n270), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(new_n267), .B2(new_n470), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n357), .B1(new_n499), .B2(new_n503), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n513), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n506), .A2(new_n512), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n502), .A2(KEYINPUT87), .A3(G87), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT87), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n297), .A2(new_n303), .A3(new_n501), .ZN(new_n525));
  INV_X1    g0325(.A(G87), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n306), .A2(new_n298), .A3(G68), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n449), .A2(new_n204), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(KEYINPUT19), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G87), .A2(G97), .ZN(new_n532));
  NAND3_X1  g0332(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n497), .A2(new_n532), .B1(new_n298), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n319), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n337), .A2(new_n444), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n528), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n306), .A2(G244), .A3(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G116), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n538), .B(new_n539), .C1(new_n415), .C2(new_n366), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n267), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n272), .A2(G1), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n280), .A2(G274), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G250), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n280), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(new_n546), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(new_n267), .B2(new_n540), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n537), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n284), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n535), .B(new_n536), .C1(new_n337), .C2(new_n525), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n357), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n252), .A2(new_n254), .A3(G257), .A4(G1698), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G294), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n366), .C2(new_n544), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n267), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n480), .A2(G264), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n517), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n380), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n562), .A2(new_n390), .A3(new_n563), .A4(new_n517), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n298), .A2(G107), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n302), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g0369(.A(new_n569), .B(KEYINPUT25), .Z(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n205), .B2(new_n525), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n252), .A2(new_n254), .A3(new_n298), .A4(G87), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n306), .A2(KEYINPUT22), .A3(new_n298), .A4(G87), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n349), .A2(G20), .A3(new_n350), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT23), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT23), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n568), .B1(new_n339), .B2(G116), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n574), .A2(new_n575), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT24), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n205), .A2(G20), .ZN(new_n582));
  INV_X1    g0382(.A(G116), .ZN(new_n583));
  OAI22_X1  g0383(.A1(KEYINPUT23), .A2(new_n582), .B1(new_n449), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(KEYINPUT23), .B2(new_n576), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT24), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n574), .A4(new_n575), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n571), .B1(new_n588), .B2(new_n319), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT91), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n567), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n567), .B2(new_n589), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n558), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n306), .A2(new_n249), .A3(G257), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n306), .A2(G264), .A3(G1698), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n255), .A2(G303), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT88), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT88), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n594), .A2(new_n595), .A3(new_n599), .A4(new_n596), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n267), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n480), .A2(G270), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n517), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n296), .A2(new_n210), .B1(G20), .B2(new_n583), .ZN(new_n606));
  AOI21_X1  g0406(.A(G20), .B1(G33), .B2(G283), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n253), .A2(G97), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT89), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n607), .B2(new_n608), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n606), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(KEYINPUT20), .B(new_n606), .C1(new_n610), .C2(new_n611), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n303), .A2(G116), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n502), .B2(G116), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n284), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n605), .A2(new_n619), .A3(KEYINPUT21), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT21), .B1(new_n605), .B2(new_n619), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n601), .A2(new_n604), .A3(G179), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n616), .A2(new_n618), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT90), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n280), .B1(new_n597), .B2(KEYINPUT88), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n603), .B1(new_n627), .B2(new_n600), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n624), .A4(G179), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n605), .A2(G200), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n632), .B(new_n625), .C1(new_n390), .C2(new_n605), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n564), .A2(new_n284), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n297), .B1(new_n581), .B2(new_n587), .ZN(new_n635));
  OAI221_X1 g0435(.A(new_n634), .B1(G179), .B2(new_n564), .C1(new_n635), .C2(new_n571), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n622), .A2(new_n631), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  NOR4_X1   g0437(.A1(new_n463), .A2(new_n522), .A3(new_n593), .A4(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n378), .ZN(new_n639));
  INV_X1    g0439(.A(new_n459), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n456), .A2(KEYINPUT77), .A3(new_n457), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n363), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n453), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n440), .B2(new_n441), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n403), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n335), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT92), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n413), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n411), .A2(KEYINPUT92), .A3(new_n412), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n639), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n513), .A2(new_n514), .A3(new_n520), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n514), .B1(new_n513), .B2(new_n520), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n553), .A2(new_n557), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n567), .A2(new_n589), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT91), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n567), .A2(new_n589), .A3(new_n590), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n622), .A2(new_n631), .A3(new_n636), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n654), .A2(new_n512), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n558), .B1(new_n652), .B2(new_n653), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT26), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n655), .A2(new_n487), .A3(new_n505), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n661), .A2(new_n663), .A3(new_n557), .A4(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n651), .B1(new_n668), .B2(new_n463), .ZN(G369));
  NAND2_X1  g0469(.A1(new_n622), .A2(new_n631), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n302), .A2(new_n298), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G343), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n624), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n622), .A2(new_n631), .A3(new_n633), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(KEYINPUT93), .B(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n589), .A2(new_n676), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n657), .B2(new_n658), .ZN(new_n686));
  INV_X1    g0486(.A(new_n636), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n676), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n684), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n686), .A2(new_n670), .A3(new_n636), .A4(new_n676), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(new_n689), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n214), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n209), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n477), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n497), .A2(new_n583), .A3(new_n532), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n655), .B1(new_n506), .B2(new_n521), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT97), .B1(new_n704), .B2(KEYINPUT26), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT97), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n662), .A2(new_n706), .A3(new_n665), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n664), .A2(KEYINPUT26), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n557), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n522), .A2(new_n593), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n660), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n677), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT29), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n667), .A2(new_n676), .ZN(new_n715));
  XOR2_X1   g0515(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n601), .A2(new_n604), .A3(G179), .ZN(new_n719));
  AND4_X1   g0519(.A1(new_n563), .A2(new_n541), .A3(new_n562), .A4(new_n547), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(new_n484), .A3(new_n486), .A4(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n548), .A2(new_n357), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT94), .B1(new_n724), .B2(new_n628), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT94), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n605), .A2(new_n726), .A3(new_n357), .A4(new_n548), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n725), .A2(new_n727), .A3(new_n483), .A4(new_n564), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n509), .A2(KEYINPUT30), .A3(new_n719), .A4(new_n720), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n723), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT31), .B1(new_n730), .B2(new_n677), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT95), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n677), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT95), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n738), .A3(new_n731), .ZN(new_n739));
  OR4_X1    g0539(.A1(new_n522), .A2(new_n637), .A3(new_n593), .A4(new_n677), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n734), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n683), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n718), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n703), .B1(new_n743), .B2(G1), .ZN(G364));
  INV_X1    g0544(.A(new_n684), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n681), .A2(new_n683), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n301), .A2(G20), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G45), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT98), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n700), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n745), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT99), .ZN(new_n752));
  INV_X1    g0552(.A(new_n750), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n210), .B1(G20), .B2(new_n284), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n298), .B1(new_n756), .B2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n204), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n298), .A2(new_n357), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(new_n390), .A3(new_n380), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR4_X1   g0561(.A1(new_n298), .A2(new_n357), .A3(new_n380), .A4(G190), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n761), .A2(new_n341), .B1(new_n762), .B2(G68), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(G190), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n763), .B1(new_n288), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n764), .A2(new_n380), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n758), .B(new_n767), .C1(G50), .C2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT102), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n298), .B2(G190), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n380), .A2(G179), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n390), .A2(KEYINPUT102), .A3(G20), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G107), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n772), .A2(G20), .A3(G190), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n776), .B(new_n306), .C1(new_n526), .C2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT103), .Z(new_n779));
  NAND3_X1  g0579(.A1(new_n771), .A2(new_n773), .A3(new_n756), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n769), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT104), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n757), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n761), .A2(G311), .B1(new_n787), .B2(G294), .ZN(new_n788));
  INV_X1    g0588(.A(new_n768), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT105), .B(G326), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT106), .Z(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT33), .B(G317), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n306), .B1(new_n762), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G303), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n797), .B2(new_n777), .C1(new_n766), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n780), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n794), .B(new_n799), .C1(G329), .C2(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n784), .A2(new_n785), .B1(new_n792), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n755), .B1(new_n786), .B2(new_n802), .ZN(new_n803));
  OR3_X1    g0603(.A1(KEYINPUT101), .A2(G13), .A3(G33), .ZN(new_n804));
  OAI21_X1  g0604(.A(KEYINPUT101), .B1(G13), .B2(G33), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n754), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n696), .A2(new_n255), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n810), .A2(G355), .B1(new_n583), .B2(new_n696), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n246), .A2(G45), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT100), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n696), .A2(new_n306), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(G45), .B2(new_n208), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n811), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n753), .B(new_n803), .C1(new_n809), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n808), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n681), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n752), .A2(new_n819), .ZN(G396));
  OAI21_X1  g0620(.A(new_n381), .B1(new_n346), .B2(new_n676), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n363), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n363), .A2(new_n677), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n715), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n667), .A2(new_n676), .A3(new_n824), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n750), .B1(new_n828), .B2(new_n742), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n742), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n830), .A2(KEYINPUT108), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(KEYINPUT108), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n806), .A2(new_n754), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n750), .B1(G77), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n789), .A2(new_n797), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n758), .B(new_n837), .C1(G294), .C2(new_n765), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n800), .A2(G311), .ZN(new_n839));
  INV_X1    g0639(.A(new_n762), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n840), .A2(new_n793), .B1(new_n205), .B2(new_n777), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n306), .B(new_n841), .C1(G116), .C2(new_n761), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n774), .A2(new_n526), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n838), .A2(new_n839), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n761), .A2(G159), .B1(new_n762), .B2(G150), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n765), .A2(G143), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n789), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n775), .A2(G68), .ZN(new_n853));
  INV_X1    g0653(.A(G50), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n306), .B1(new_n757), .B2(new_n288), .C1(new_n777), .C2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(G132), .B2(new_n800), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n845), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n836), .B1(new_n858), .B2(new_n754), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n824), .B2(new_n807), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT107), .Z(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n833), .A2(new_n862), .ZN(G384));
  NOR3_X1   g0663(.A1(new_n210), .A2(new_n298), .A3(new_n583), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT35), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(new_n495), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n865), .B2(new_n495), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT36), .ZN(new_n868));
  OR3_X1    g0668(.A1(new_n220), .A2(new_n208), .A3(new_n311), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n854), .A2(G68), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n477), .B(G13), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n385), .A2(new_n322), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n305), .B1(new_n320), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n675), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n335), .B2(new_n403), .ZN(new_n877));
  INV_X1    g0677(.A(new_n279), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n284), .B1(new_n268), .B2(new_n278), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n332), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n332), .A2(new_n675), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n880), .A2(new_n393), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(KEYINPUT110), .B(KEYINPUT37), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n285), .A2(new_n875), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n393), .A3(new_n876), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n882), .A2(new_n883), .B1(new_n885), .B2(KEYINPUT37), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n873), .B1(new_n877), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n876), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n400), .A2(new_n401), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n393), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n880), .A2(KEYINPUT18), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n285), .A2(new_n286), .A3(new_n332), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n888), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n885), .A2(KEYINPUT37), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n880), .A2(new_n393), .A3(new_n881), .A4(new_n883), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n887), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT111), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT111), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n887), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n643), .A2(new_n676), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n454), .A2(new_n461), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n906), .B1(new_n644), .B2(new_n460), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n823), .B(KEYINPUT109), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n827), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n905), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n454), .A2(new_n677), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n887), .A2(new_n900), .A3(KEYINPUT39), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT112), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n883), .B1(new_n881), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n880), .A2(new_n393), .A3(new_n881), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n882), .A2(new_n918), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n881), .B1(new_n335), .B2(new_n403), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n873), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n925), .A2(new_n900), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n915), .B(new_n916), .C1(new_n926), .C2(KEYINPUT39), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n895), .A2(new_n674), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n914), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n714), .A2(new_n462), .A3(new_n717), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n651), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT40), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n732), .A2(new_n733), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n825), .B1(new_n935), .B2(new_n740), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n907), .B1(new_n454), .B2(new_n461), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n644), .A2(new_n460), .A3(new_n906), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n887), .A2(new_n900), .A3(new_n903), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n903), .B1(new_n887), .B2(new_n900), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n934), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n934), .B1(new_n925), .B2(new_n900), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n936), .B(new_n944), .C1(new_n937), .C2(new_n938), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n935), .A2(new_n740), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n462), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n682), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n946), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n933), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n477), .B2(new_n747), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n933), .A2(new_n950), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n872), .B1(new_n952), .B2(new_n953), .ZN(G367));
  INV_X1    g0754(.A(KEYINPUT117), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n537), .A2(new_n676), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n558), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n557), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n504), .A2(new_n677), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n654), .A2(new_n512), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n513), .A2(new_n520), .A3(new_n677), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n693), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT42), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n636), .B1(new_n963), .B2(new_n964), .ZN(new_n968));
  INV_X1    g0768(.A(new_n654), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n676), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n965), .A2(new_n966), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n967), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n961), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n963), .A2(new_n964), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n691), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n972), .A2(new_n961), .A3(new_n973), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n978), .B1(new_n975), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n749), .A2(new_n477), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n694), .B2(new_n976), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n693), .A2(new_n689), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n988), .A2(KEYINPUT44), .A3(new_n963), .A4(new_n964), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n991));
  NAND3_X1  g0791(.A1(new_n694), .A2(new_n976), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n694), .A2(new_n976), .ZN(new_n993));
  INV_X1    g0793(.A(new_n991), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n990), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n691), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n692), .A2(new_n990), .A3(new_n992), .A4(new_n995), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n670), .A2(new_n676), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n690), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n693), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n745), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n684), .A3(new_n693), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n718), .A2(new_n1005), .A3(new_n742), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n743), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n697), .B(KEYINPUT41), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n985), .B1(new_n1010), .B2(KEYINPUT114), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n743), .A2(new_n1005), .A3(new_n997), .A4(new_n998), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1008), .B1(new_n1012), .B2(new_n743), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT114), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n983), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n814), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n809), .B1(new_n239), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n696), .B2(new_n338), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n760), .A2(new_n854), .B1(new_n777), .B2(new_n288), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n255), .B(new_n1020), .C1(G159), .C2(new_n762), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n848), .B2(new_n780), .C1(new_n220), .C2(new_n774), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n757), .A2(new_n219), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n768), .B2(G143), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n373), .B2(new_n766), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n777), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1027), .A2(KEYINPUT115), .B1(G97), .B2(new_n775), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(KEYINPUT115), .B2(new_n1027), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT46), .B1(new_n1026), .B2(G116), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n351), .B2(new_n787), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G303), .A2(new_n765), .B1(new_n768), .B2(G311), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n800), .A2(G317), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n255), .B1(new_n760), .B2(new_n793), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G294), .B2(new_n762), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1022), .A2(new_n1025), .B1(new_n1029), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(KEYINPUT116), .B(KEYINPUT47), .Z(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n753), .B(new_n1019), .C1(new_n1039), .C2(new_n754), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n957), .A2(new_n808), .A3(new_n958), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n955), .B1(new_n1016), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n984), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1010), .A2(KEYINPUT114), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n982), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1047), .A2(KEYINPUT117), .A3(new_n1042), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(G387));
  OR2_X1    g0850(.A1(new_n236), .A2(new_n272), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1051), .A2(new_n814), .B1(new_n701), .B2(new_n810), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n342), .A2(new_n854), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n272), .B1(new_n219), .B2(new_n202), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1054), .A2(new_n701), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1052), .A2(new_n1056), .B1(G107), .B2(new_n214), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n753), .B1(new_n1057), .B2(new_n809), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n306), .B1(new_n775), .B2(G116), .ZN(new_n1059));
  INV_X1    g0859(.A(G294), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n777), .A2(new_n1060), .B1(new_n757), .B2(new_n793), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n761), .A2(G303), .B1(new_n762), .B2(G311), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n765), .A2(G317), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n798), .C2(new_n789), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT48), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1061), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT49), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1059), .B1(new_n780), .B2(new_n790), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n338), .A2(new_n787), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n854), .B2(new_n766), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT118), .Z(new_n1073));
  OAI22_X1  g0873(.A1(new_n204), .A2(new_n774), .B1(new_n780), .B2(new_n373), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n255), .B1(new_n761), .B2(G68), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n341), .A2(new_n1026), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n781), .C2(new_n789), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1074), .B(new_n1077), .C1(new_n295), .C2(new_n762), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1070), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1058), .B1(new_n1079), .B2(new_n755), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n690), .B2(new_n808), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1005), .B2(new_n985), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n697), .B(KEYINPUT119), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1006), .A2(KEYINPUT120), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n743), .B2(new_n1005), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT120), .B1(new_n1006), .B2(new_n1083), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1082), .B1(new_n1085), .B2(new_n1086), .ZN(G393));
  INV_X1    g0887(.A(KEYINPUT121), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n998), .A2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(new_n997), .Z(new_n1090));
  INV_X1    g0890(.A(new_n1006), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1012), .B(new_n1083), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n963), .A2(new_n808), .A3(new_n964), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n761), .A2(new_n342), .B1(new_n762), .B2(G50), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n202), .B2(new_n757), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT122), .Z(new_n1096));
  AOI22_X1  g0896(.A1(G150), .A2(new_n768), .B1(new_n765), .B2(G159), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT51), .Z(new_n1098));
  OAI21_X1  g0898(.A(new_n306), .B1(new_n777), .B2(new_n219), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1099), .B(new_n843), .C1(G143), .C2(new_n800), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n255), .B1(new_n777), .B2(new_n793), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n840), .A2(new_n797), .B1(new_n760), .B2(new_n1060), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(G116), .C2(new_n787), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G311), .A2(new_n765), .B1(new_n768), .B2(G317), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT123), .B(KEYINPUT52), .Z(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n800), .A2(G322), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1104), .A2(new_n1107), .A3(new_n776), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n755), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n243), .A2(new_n814), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n754), .B(new_n808), .C1(G97), .C2(new_n696), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n753), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1090), .A2(new_n985), .B1(new_n1093), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1092), .A2(new_n1114), .ZN(G390));
  OAI21_X1  g0915(.A(new_n916), .B1(new_n926), .B2(KEYINPUT39), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n908), .A2(new_n909), .B1(new_n827), .B2(new_n912), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n915), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n926), .A2(new_n915), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n911), .B1(new_n713), .B2(new_n824), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n937), .A2(new_n938), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n737), .A2(new_n731), .ZN(new_n1124));
  NOR4_X1   g0924(.A1(new_n522), .A2(new_n637), .A3(new_n593), .A4(new_n677), .ZN(new_n1125));
  OAI211_X1 g0925(.A(G330), .B(new_n824), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n908), .B2(new_n909), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n910), .A2(new_n683), .A3(new_n741), .A4(new_n824), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1118), .A2(new_n1122), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n462), .A2(G330), .A3(new_n947), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n651), .A2(new_n931), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1126), .A2(new_n908), .A3(new_n909), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1129), .A2(new_n1120), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n913), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n741), .A2(new_n683), .A3(new_n824), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1121), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n910), .A2(G330), .A3(new_n936), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1138), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1134), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1131), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1127), .B1(new_n1121), .B2(new_n1139), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1136), .B1(new_n1145), .B2(new_n1138), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1128), .A2(new_n1146), .A3(new_n1130), .A4(new_n1134), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1144), .A2(new_n1083), .A3(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1118), .A2(new_n1122), .A3(new_n1129), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1141), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1116), .A2(new_n806), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n750), .B1(new_n295), .B2(new_n835), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n306), .B1(new_n760), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1026), .A2(G150), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1156), .A2(KEYINPUT53), .B1(new_n781), .B2(new_n757), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G137), .C2(new_n762), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(KEYINPUT53), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G128), .A2(new_n768), .B1(new_n765), .B2(G132), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G50), .A2(new_n775), .B1(new_n800), .B2(G125), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT124), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n757), .A2(new_n202), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n789), .A2(new_n793), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(G116), .C2(new_n765), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n840), .A2(new_n497), .B1(new_n760), .B2(new_n204), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n306), .B(new_n1168), .C1(G87), .C2(new_n1026), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n800), .A2(G294), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n853), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1164), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1153), .B1(new_n1173), .B2(new_n754), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1151), .A2(new_n985), .B1(new_n1152), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1148), .A2(new_n1175), .ZN(G378));
  OAI21_X1  g0976(.A(new_n824), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n908), .B2(new_n909), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT40), .B1(new_n1178), .B2(new_n905), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n945), .A2(G330), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n648), .A2(new_n378), .A3(new_n649), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n404), .A2(new_n674), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1182), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n648), .A2(new_n378), .A3(new_n649), .A4(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1179), .A2(new_n1180), .A3(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1191));
  INV_X1    g0991(.A(G330), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1178), .B2(new_n944), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1191), .B1(new_n943), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n930), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1189), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n943), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n914), .A2(new_n929), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1189), .A2(new_n806), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n750), .B1(G50), .B2(new_n835), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n306), .A2(G41), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G50), .B(new_n1203), .C1(new_n253), .C2(new_n271), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n789), .A2(new_n583), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1023), .B(new_n1205), .C1(G107), .C2(new_n765), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1076), .B(new_n1203), .C1(new_n204), .C2(new_n840), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n338), .B2(new_n761), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n775), .A2(G58), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n800), .A2(G283), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1206), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1204), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n765), .A2(G128), .B1(G150), .B2(new_n787), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1154), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1026), .A2(new_n1216), .B1(new_n762), .B2(G132), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n848), .B2(new_n760), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1215), .B(new_n1218), .C1(G125), .C2(new_n768), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(KEYINPUT59), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n253), .B(new_n271), .C1(new_n774), .C2(new_n781), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G124), .B2(new_n800), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT59), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .C1(new_n1221), .C2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1202), .B1(new_n1226), .B2(new_n754), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1200), .A2(new_n985), .B1(new_n1201), .B2(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1198), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT57), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n913), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1133), .B1(new_n1233), .B2(new_n1136), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1133), .B1(new_n1151), .B2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1083), .B1(new_n1231), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1134), .B1(new_n1131), .B2(new_n1143), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1237), .B2(new_n1200), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1228), .B1(new_n1236), .B2(new_n1238), .ZN(G375));
  OAI211_X1 g1039(.A(new_n1133), .B(new_n1136), .C1(new_n1145), .C2(new_n1138), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1143), .A2(new_n1009), .A3(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT125), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1121), .A2(new_n806), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n750), .B1(G68), .B2(new_n835), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1071), .B1(new_n202), .B2(new_n774), .C1(new_n797), .C2(new_n780), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G283), .A2(new_n765), .B1(new_n768), .B2(G294), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n306), .B1(new_n1026), .B2(G97), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n761), .A2(new_n351), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n762), .A2(G116), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n768), .A2(G132), .B1(G50), .B2(new_n787), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n848), .B2(new_n766), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1026), .A2(G159), .B1(new_n762), .B2(new_n1216), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n255), .B1(new_n761), .B2(G150), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n800), .A2(G128), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1209), .A4(new_n1255), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1245), .A2(new_n1250), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1244), .B1(new_n1257), .B2(new_n754), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1146), .A2(new_n985), .B1(new_n1243), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1242), .A2(new_n1259), .ZN(G381));
  AND2_X1   g1060(.A1(new_n1092), .A2(new_n1114), .ZN(new_n1261));
  INV_X1    g1061(.A(G384), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(G396), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1264), .B(new_n1082), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1263), .A2(G381), .A3(G378), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G375), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1049), .A3(new_n1267), .ZN(G407));
  OR2_X1    g1068(.A1(G378), .A2(G343), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G375), .C2(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(G213), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(G343), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1240), .A2(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1233), .A2(KEYINPUT60), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1083), .A3(new_n1275), .A4(new_n1143), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(G384), .A3(new_n1259), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1276), .B2(new_n1259), .ZN(new_n1279));
  OAI211_X1 g1079(.A(G2897), .B(new_n1272), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1279), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1272), .A2(G2897), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1277), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G378), .B(new_n1228), .C1(new_n1236), .C2(new_n1238), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1152), .A2(new_n1174), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n1131), .B2(new_n984), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1083), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1151), .B2(new_n1234), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1144), .B2(new_n1290), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1237), .A2(new_n1200), .A3(new_n1009), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1201), .A2(new_n1227), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(new_n984), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1291), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1286), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1272), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT63), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1301), .B1(new_n1299), .B2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1044), .A2(new_n1048), .A3(new_n1261), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G393), .A2(G396), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1306), .A2(new_n1265), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1016), .A2(new_n1043), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1308), .B2(G390), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1306), .A2(KEYINPUT126), .A3(new_n1265), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT126), .B1(new_n1306), .B2(new_n1265), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1261), .A2(new_n1016), .A3(new_n1043), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G390), .B1(new_n1047), .B2(new_n1042), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1310), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1272), .B1(new_n1286), .B2(new_n1296), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(KEYINPUT63), .A3(new_n1302), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1300), .A2(new_n1304), .A3(new_n1317), .A4(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1318), .A2(new_n1321), .A3(new_n1302), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1323), .B1(new_n1318), .B2(new_n1284), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1321), .B1(new_n1318), .B2(new_n1302), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1322), .A2(new_n1324), .A3(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1320), .B1(new_n1326), .B2(new_n1317), .ZN(G405));
  INV_X1    g1127(.A(KEYINPUT127), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1317), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1310), .A2(KEYINPUT127), .A3(new_n1316), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(G375), .A2(new_n1291), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1303), .B1(new_n1331), .B2(new_n1286), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1331), .A2(new_n1303), .A3(new_n1286), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1329), .B(new_n1330), .C1(new_n1332), .C2(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1332), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1335), .A2(new_n1328), .A3(new_n1317), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1336), .ZN(G402));
endmodule


