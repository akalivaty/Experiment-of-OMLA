//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(G319));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n466), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(G101), .A3(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n469), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n468), .A2(G136), .ZN(new_n480));
  AND2_X1   g055(.A1(G112), .A2(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n481), .B1(G100), .B2(new_n476), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n464), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n485), .B(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n483), .B1(new_n487), .B2(G124), .ZN(G162));
  NAND3_X1  g063(.A1(new_n484), .A2(KEYINPUT4), .A3(G138), .ZN(new_n489));
  INV_X1    g064(.A(G102), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(new_n464), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n476), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n493), .A2(KEYINPUT71), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(KEYINPUT71), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n467), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n471), .A2(new_n466), .A3(G138), .A4(new_n476), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n498), .A2(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n509), .A2(new_n518), .ZN(G166));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(new_n522), .B1(new_n504), .B2(new_n505), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(new_n516), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(new_n506), .A2(G64), .ZN(new_n529));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n508), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n506), .A2(new_n520), .A3(G90), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n520), .A2(G52), .A3(G543), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n535), .B1(new_n533), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(G171));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT73), .B(G43), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n514), .A2(new_n540), .B1(new_n516), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(G56), .B1(new_n511), .B2(new_n510), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n508), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(new_n513), .ZN(new_n553));
  NAND2_X1  g128(.A1(KEYINPUT6), .A2(G651), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n553), .A2(new_n554), .B1(new_n504), .B2(new_n505), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G91), .ZN(new_n556));
  INV_X1    g131(.A(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n553), .B2(new_n554), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n558), .A2(new_n559), .A3(G53), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n559), .B1(new_n558), .B2(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n504), .A2(new_n564), .A3(new_n505), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT74), .B1(new_n511), .B2(new_n510), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n563), .B1(new_n567), .B2(G65), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n508), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(new_n565), .B2(new_n566), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT75), .B1(new_n572), .B2(new_n563), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n562), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G299));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n533), .A2(new_n534), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT72), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n576), .B1(new_n580), .B2(new_n532), .ZN(new_n581));
  AOI211_X1 g156(.A(KEYINPUT76), .B(new_n531), .C1(new_n578), .C2(new_n579), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G301));
  INV_X1    g158(.A(G168), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  AND3_X1   g160(.A1(new_n506), .A2(new_n520), .A3(G87), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT77), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n506), .A2(G74), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n558), .B2(G49), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n555), .A2(G86), .B1(new_n558), .B2(G48), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n506), .A2(G61), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT78), .B1(new_n594), .B2(G651), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n596));
  AOI211_X1 g171(.A(new_n596), .B(new_n508), .C1(new_n592), .C2(new_n593), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n591), .B1(new_n595), .B2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n508), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n514), .A2(new_n601), .B1(new_n516), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n600), .A2(new_n603), .ZN(G290));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n565), .B2(new_n566), .ZN(new_n606));
  AND2_X1   g181(.A1(G79), .A2(G543), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n555), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n514), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n558), .A2(G54), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n608), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G301), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n616), .ZN(G284));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(new_n616), .ZN(G321));
  NOR2_X1   g195(.A1(G286), .A2(new_n616), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n574), .B2(new_n616), .ZN(G297));
  AOI21_X1  g197(.A(new_n621), .B1(new_n574), .B2(new_n616), .ZN(G280));
  INV_X1    g198(.A(new_n615), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G860), .ZN(G148));
  NOR3_X1   g201(.A1(new_n542), .A2(G868), .A3(new_n545), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n615), .A2(G559), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(KEYINPUT81), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G111), .B2(new_n476), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(KEYINPUT81), .B2(new_n631), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n487), .A2(G123), .ZN(new_n635));
  AOI211_X1 g210(.A(new_n634), .B(new_n635), .C1(G135), .C2(new_n468), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(KEYINPUT80), .B2(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(KEYINPUT80), .A2(G2100), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n637), .A2(new_n644), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT15), .B(G2435), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2427), .ZN(new_n649));
  INV_X1    g224(.A(G2430), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n652), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT84), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n668), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n671), .B(new_n667), .C1(new_n664), .C2(new_n668), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n666), .A2(new_n664), .A3(new_n668), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2096), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n682), .A2(new_n683), .ZN(new_n690));
  INV_X1    g265(.A(new_n684), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n681), .B2(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n687), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n697), .B(new_n700), .ZN(G229));
  NAND2_X1  g276(.A1(G164), .A2(G29), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G27), .B2(G29), .ZN(new_n703));
  INV_X1    g278(.A(G2078), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G32), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n468), .A2(G141), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n476), .A2(G105), .A3(G2104), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT26), .Z(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n487), .B2(G129), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n707), .B1(new_n713), .B2(new_n706), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT27), .B(G1996), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n705), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n715), .B2(new_n716), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G19), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n546), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1341), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n636), .B2(G29), .ZN(new_n723));
  AND2_X1   g298(.A1(KEYINPUT24), .A2(G34), .ZN(new_n724));
  NOR2_X1   g299(.A1(KEYINPUT24), .A2(G34), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n706), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n478), .B2(new_n706), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2084), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n723), .B(new_n728), .C1(new_n704), .C2(new_n703), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT31), .B(G11), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT30), .B(G28), .Z(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G29), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G21), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G168), .B2(new_n733), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT94), .B(G1966), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n732), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n624), .A2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G4), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G1348), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n738), .B1(new_n735), .B2(new_n737), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n706), .A2(G33), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT25), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n471), .A2(new_n466), .A3(G127), .ZN(new_n746));
  NAND2_X1  g321(.A1(G115), .A2(G2104), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n476), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n745), .B(new_n748), .C1(G139), .C2(new_n468), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n749), .B2(new_n706), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G2072), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n740), .A2(new_n741), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n719), .A2(new_n729), .A3(new_n742), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n706), .A2(G26), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT28), .Z(new_n756));
  MUX2_X1   g331(.A(G104), .B(G116), .S(G2105), .Z(new_n757));
  AOI22_X1  g332(.A1(new_n468), .A2(G140), .B1(G2104), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n485), .B(KEYINPUT70), .ZN(new_n759));
  INV_X1    g334(.A(G128), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n756), .B1(new_n765), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT93), .B(G2067), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n754), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G2090), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT96), .Z(new_n774));
  NOR2_X1   g349(.A1(G5), .A2(G16), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G171), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT95), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n733), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1956), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n778), .B(new_n782), .C1(G2090), .C2(new_n772), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n769), .A2(new_n774), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n706), .A2(G25), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n487), .A2(G119), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT87), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n476), .A2(G95), .ZN(new_n789));
  NAND2_X1  g364(.A1(G107), .A2(G2105), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n464), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n468), .B2(G131), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT88), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n786), .B1(new_n794), .B2(new_n706), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT35), .B(G1991), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G16), .A2(G24), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n600), .A2(new_n603), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT89), .ZN(new_n801));
  INV_X1    g376(.A(G1986), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n733), .A2(G23), .ZN(new_n804));
  INV_X1    g379(.A(G288), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n733), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT90), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT33), .B(G1976), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G6), .B(G305), .S(G16), .Z(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT32), .B(G1981), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G22), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G166), .B2(G16), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1971), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n803), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n797), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n809), .A2(new_n816), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT91), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n820), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n785), .B1(new_n825), .B2(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n784), .ZN(G150));
  NOR2_X1   g405(.A1(new_n546), .A2(KEYINPUT99), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n555), .A2(G93), .B1(new_n558), .B2(G55), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n833));
  OAI21_X1  g408(.A(G67), .B1(new_n511), .B2(new_n510), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n833), .B1(new_n836), .B2(G651), .ZN(new_n837));
  AOI211_X1 g412(.A(KEYINPUT98), .B(new_n508), .C1(new_n834), .C2(new_n835), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n542), .A2(new_n840), .A3(new_n545), .ZN(new_n841));
  OAI21_X1  g416(.A(KEYINPUT100), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT98), .B1(new_n843), .B2(new_n508), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n836), .A2(new_n833), .A3(G651), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT100), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n555), .A2(G81), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n516), .A2(new_n541), .ZN(new_n849));
  INV_X1    g424(.A(G56), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n504), .B2(new_n505), .ZN(new_n851));
  INV_X1    g426(.A(new_n544), .ZN(new_n852));
  OAI21_X1  g427(.A(G651), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n848), .A2(new_n849), .A3(new_n853), .A4(KEYINPUT99), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n846), .A2(new_n847), .A3(new_n854), .A4(new_n832), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n831), .B1(new_n842), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n842), .A2(new_n831), .A3(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n615), .A2(new_n625), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n859), .B(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n839), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  INV_X1    g445(.A(new_n765), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G164), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n765), .A2(new_n502), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n713), .B(new_n749), .Z(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  MUX2_X1   g452(.A(G106), .B(G118), .S(G2105), .Z(new_n878));
  AOI22_X1  g453(.A1(new_n468), .A2(G142), .B1(G2104), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G130), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n759), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n639), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n793), .B(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(G162), .B(G160), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n636), .B(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n877), .A2(new_n884), .ZN(new_n889));
  INV_X1    g464(.A(new_n883), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n893), .A2(new_n894), .A3(new_n891), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n892), .B1(new_n895), .B2(new_n887), .ZN(new_n896));
  XNOR2_X1  g471(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(G395));
  AND3_X1   g473(.A1(new_n842), .A2(new_n831), .A3(new_n855), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n899), .A2(new_n856), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n628), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n568), .A2(new_n569), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(G651), .A3(new_n573), .ZN(new_n903));
  INV_X1    g478(.A(new_n562), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n615), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT103), .B1(new_n574), .B2(new_n615), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n574), .A2(new_n615), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n901), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n903), .A2(new_n904), .A3(new_n615), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(new_n914), .B2(new_n905), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n907), .A2(new_n908), .A3(KEYINPUT41), .A4(new_n909), .ZN(new_n918));
  OAI211_X1 g493(.A(KEYINPUT104), .B(new_n913), .C1(new_n914), .C2(new_n905), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n912), .B1(new_n901), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n912), .B(KEYINPUT42), .C1(new_n901), .C2(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  NAND2_X1  g502(.A1(G290), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n799), .A2(KEYINPUT105), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n928), .A2(G288), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G288), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G305), .B(G166), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n926), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR4_X1   g510(.A1(new_n933), .A2(new_n930), .A3(new_n931), .A4(KEYINPUT106), .ZN(new_n936));
  OAI22_X1  g511(.A1(new_n935), .A2(new_n936), .B1(new_n932), .B2(new_n934), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT107), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n925), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n938), .A4(new_n924), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(G868), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n839), .A2(G868), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT108), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n616), .B1(new_n940), .B2(new_n941), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n947), .A2(new_n948), .A3(new_n944), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n946), .A2(new_n949), .ZN(G295));
  NOR2_X1   g525(.A1(new_n947), .A2(new_n944), .ZN(G331));
  OAI21_X1  g526(.A(G168), .B1(new_n581), .B2(new_n582), .ZN(new_n952));
  NAND2_X1  g527(.A1(G286), .A2(new_n538), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(KEYINPUT109), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n538), .A2(KEYINPUT76), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n580), .A2(new_n576), .A3(new_n532), .ZN(new_n957));
  AOI21_X1  g532(.A(G286), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n953), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n900), .A2(new_n954), .A3(new_n960), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n960), .A2(new_n954), .B1(new_n858), .B2(new_n857), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n920), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n958), .A2(new_n955), .A3(new_n959), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT109), .B1(new_n952), .B2(new_n953), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n859), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n900), .A2(new_n960), .A3(new_n954), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n910), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n963), .A2(new_n937), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT111), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n963), .A2(new_n937), .A3(new_n968), .A4(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G37), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n905), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT41), .A3(new_n909), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n974), .A2(new_n909), .A3(KEYINPUT112), .A4(KEYINPUT41), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n977), .B(new_n978), .C1(new_n911), .C2(KEYINPUT41), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n961), .B2(new_n962), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n966), .A2(new_n981), .A3(new_n910), .A4(new_n967), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n968), .A2(KEYINPUT113), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n938), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n973), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n963), .A2(KEYINPUT110), .A3(new_n968), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT110), .B1(new_n963), .B2(new_n968), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n938), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n973), .A2(KEYINPUT43), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT44), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n970), .A2(new_n972), .ZN(new_n995));
  INV_X1    g570(.A(G37), .ZN(new_n996));
  AND4_X1   g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n985), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n994), .B1(new_n973), .B2(new_n985), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n973), .A2(new_n987), .A3(new_n991), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n993), .B1(new_n1001), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n502), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G160), .A2(G40), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n765), .A2(G2067), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n765), .A2(G2067), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1009), .B1(new_n1012), .B2(new_n713), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1009), .A2(G1996), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT46), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT47), .Z(new_n1017));
  NAND3_X1  g592(.A1(new_n794), .A2(KEYINPUT125), .A3(new_n796), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n713), .B(G1996), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1012), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT125), .B1(new_n794), .B2(new_n796), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1010), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n1008), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n793), .B(new_n796), .Z(new_n1025));
  OAI21_X1  g600(.A(new_n1008), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT126), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(KEYINPUT126), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1008), .A2(new_n802), .A3(new_n799), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT48), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1017), .A2(new_n1023), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1007), .B1(new_n1004), .B2(KEYINPUT50), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n492), .B2(new_n501), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(G2090), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1007), .B1(new_n1034), .B2(KEYINPUT45), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1971), .B1(new_n1006), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(G8), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  OAI211_X1 g617(.A(G303), .B(G8), .C1(new_n1042), .C2(KEYINPUT55), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(KEYINPUT55), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1043), .B(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1007), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(new_n1034), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G305), .B(G1981), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(KEYINPUT118), .A3(new_n1052), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n805), .A2(G1976), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1050), .A2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT117), .B(G1976), .Z(new_n1061));
  NOR2_X1   g636(.A1(new_n805), .A2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1060), .A2(KEYINPUT52), .A3(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1060), .A2(KEYINPUT52), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1058), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1040), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1036), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1034), .A2(KEYINPUT115), .A3(new_n1035), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1033), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1066), .B1(new_n1070), .B2(G2090), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(G8), .A3(new_n1045), .ZN(new_n1072));
  INV_X1    g647(.A(G2084), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1068), .A2(new_n1033), .A3(new_n1073), .A4(new_n1069), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1006), .A2(new_n1039), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n736), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1048), .B(G286), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1047), .A2(new_n1065), .A3(new_n1072), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT63), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1077), .A2(KEYINPUT63), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1071), .A2(G8), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1046), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1081), .A2(new_n1083), .A3(new_n1072), .A4(new_n1065), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1072), .ZN(new_n1086));
  OR2_X1    g661(.A1(G288), .A2(G1976), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1058), .A2(new_n1087), .B1(G1981), .B2(G305), .ZN(new_n1088));
  XOR2_X1   g663(.A(new_n1050), .B(KEYINPUT119), .Z(new_n1089));
  AOI22_X1  g664(.A1(new_n1086), .A2(new_n1065), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1074), .A2(new_n1076), .A3(G168), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT51), .ZN(new_n1093));
  AOI21_X1  g668(.A(G168), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  OAI211_X1 g670(.A(G8), .B(new_n1091), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1093), .A2(new_n1096), .A3(KEYINPUT62), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT62), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1047), .A2(new_n1065), .A3(new_n1072), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1070), .A2(KEYINPUT121), .ZN(new_n1101));
  INV_X1    g676(.A(G1961), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1068), .A2(new_n1033), .A3(new_n1103), .A4(new_n1069), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1101), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1006), .A2(new_n1039), .A3(new_n704), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  AOI211_X1 g682(.A(KEYINPUT123), .B(G301), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n618), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1100), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1085), .B(new_n1090), .C1(new_n1099), .C2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT120), .B1(new_n560), .B2(new_n561), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n574), .B(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1037), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1006), .A2(new_n1039), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1117), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1119), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT61), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1101), .A2(new_n741), .A3(new_n1104), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1049), .A2(new_n1034), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(G2067), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1127), .A2(new_n615), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n615), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT60), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n615), .A2(KEYINPUT60), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1127), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT58), .B(G1341), .Z(new_n1136));
  NAND2_X1  g711(.A1(new_n1128), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1075), .B2(G1996), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n546), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT59), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1126), .A2(new_n1133), .A3(new_n1135), .A4(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1124), .B1(new_n1132), .B2(new_n1122), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT122), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1111), .A2(new_n1108), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1006), .A2(new_n1039), .A3(KEYINPUT124), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1106), .B1(KEYINPUT53), .B2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1106), .A2(new_n1146), .A3(KEYINPUT53), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1105), .B(G301), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT54), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1105), .B1(new_n1148), .B2(new_n1147), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT54), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1110), .A2(new_n618), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1100), .B(new_n1151), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1113), .B1(new_n1144), .B2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n799), .B(G1986), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1026), .B1(new_n1009), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1032), .B1(new_n1158), .B2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g736(.A1(new_n662), .A2(G319), .ZN(new_n1163));
  NOR3_X1   g737(.A1(G227), .A2(G229), .A3(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g738(.A(new_n1164), .B(KEYINPUT127), .ZN(new_n1165));
  NAND4_X1  g739(.A1(new_n896), .A2(new_n1165), .A3(new_n988), .A4(new_n992), .ZN(G225));
  INV_X1    g740(.A(G225), .ZN(G308));
endmodule


