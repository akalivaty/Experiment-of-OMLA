//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  NAND2_X1  g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n191), .A2(KEYINPUT64), .A3(G146), .ZN(new_n192));
  AOI21_X1  g006(.A(KEYINPUT64), .B1(new_n191), .B2(G146), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n188), .B(new_n190), .C1(new_n192), .C2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(new_n195), .ZN(new_n196));
  OR2_X1    g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n187), .A3(new_n197), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n194), .A2(KEYINPUT68), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT68), .B1(new_n194), .B2(new_n198), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G134), .B(G137), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n203), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n202), .B1(G134), .B2(new_n208), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n207), .A2(G131), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(G134), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n202), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n212), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n199), .A2(new_n200), .B1(new_n210), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n211), .A3(new_n217), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n191), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g036(.A(G128), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n196), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n190), .B(new_n226), .C1(new_n192), .C2(new_n193), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n204), .A2(new_n211), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n220), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n219), .A2(KEYINPUT30), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT30), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n220), .A2(new_n228), .A3(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n194), .A2(new_n198), .ZN(new_n234));
  OAI21_X1  g048(.A(G131), .B1(new_n207), .B2(new_n209), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(new_n220), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n232), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G119), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT67), .B(G119), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT2), .A2(G113), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT2), .A3(G113), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT2), .A2(G113), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G119), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(KEYINPUT67), .ZN(new_n253));
  OAI21_X1  g067(.A(G116), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n247), .B1(new_n243), .B2(new_n245), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(new_n239), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n231), .A2(new_n237), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT31), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  INV_X1    g075(.A(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n257), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n219), .A2(new_n267), .A3(new_n230), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n258), .A2(new_n259), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n258), .A2(new_n266), .A3(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT31), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n270), .A3(KEYINPUT31), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n265), .B(KEYINPUT70), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n268), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n219), .A2(KEYINPUT28), .A3(new_n267), .A4(new_n230), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n257), .B1(new_n233), .B2(new_n236), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n274), .A2(new_n275), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(G472), .A2(G902), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT32), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(KEYINPUT32), .A3(new_n285), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n258), .A2(new_n268), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n265), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(KEYINPUT71), .A3(new_n265), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n276), .A2(new_n279), .A3(new_n280), .A4(new_n281), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n292), .A2(new_n293), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n200), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n194), .A2(new_n198), .A3(KEYINPUT68), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n297), .A2(new_n298), .B1(new_n235), .B2(new_n220), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n257), .B1(new_n299), .B2(new_n233), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n265), .A2(new_n293), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n279), .A2(new_n280), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n302), .A2(KEYINPUT72), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT72), .B1(new_n302), .B2(new_n303), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n296), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT73), .B1(new_n307), .B2(G472), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n309));
  INV_X1    g123(.A(G472), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n309), .B(new_n310), .C1(new_n296), .C2(new_n306), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n287), .B(new_n288), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G217), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(G234), .B2(new_n303), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT16), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(G125), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(G146), .B(new_n318), .C1(new_n322), .C2(new_n316), .ZN(new_n323));
  XNOR2_X1  g137(.A(G125), .B(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n189), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n251), .A2(G128), .ZN(new_n326));
  XOR2_X1   g140(.A(KEYINPUT67), .B(G119), .Z(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G128), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT23), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n327), .A2(KEYINPUT23), .A3(G128), .ZN(new_n330));
  AOI21_X1  g144(.A(G110), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT24), .B(G110), .Z(new_n332));
  NOR2_X1   g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n323), .B(new_n325), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(G110), .A3(new_n330), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n318), .B1(new_n322), .B2(new_n316), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n189), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n323), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n328), .A2(new_n332), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G137), .ZN(new_n341));
  INV_X1    g155(.A(G953), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(G221), .A3(G234), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n334), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(new_n334), .B2(new_n340), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT25), .A3(new_n303), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n334), .A2(new_n340), .ZN(new_n349));
  INV_X1    g163(.A(new_n344), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n334), .A2(new_n340), .A3(new_n344), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n303), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT25), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n315), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n314), .A2(G902), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n312), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT74), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G214), .B1(G237), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G104), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT3), .B1(new_n367), .B2(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(G107), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n370), .B(G101), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(G101), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n371), .A2(new_n372), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n262), .B(new_n366), .C1(new_n368), .C2(new_n369), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n257), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT5), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n327), .A2(new_n380), .A3(G116), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT5), .B(new_n239), .C1(new_n240), .C2(new_n238), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G113), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n365), .A2(G104), .ZN(new_n384));
  OAI21_X1  g198(.A(G101), .B1(new_n369), .B2(new_n384), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n376), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n256), .A3(new_n386), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n378), .A2(new_n379), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n379), .B1(new_n378), .B2(new_n387), .ZN(new_n389));
  XNOR2_X1  g203(.A(G110), .B(G122), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n378), .A2(new_n387), .A3(new_n390), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT6), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT80), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n224), .A2(new_n227), .A3(new_n320), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n395), .A2(KEYINPUT81), .B1(new_n234), .B2(G125), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n234), .A2(KEYINPUT81), .A3(G125), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G224), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G953), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n396), .B2(new_n397), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n378), .A2(new_n387), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT79), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n378), .A2(new_n379), .A3(new_n387), .ZN(new_n407));
  INV_X1    g221(.A(new_n390), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n410));
  INV_X1    g224(.A(new_n393), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n391), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n394), .A2(new_n404), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G210), .B1(G237), .B2(G902), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n390), .B(KEYINPUT8), .ZN(new_n417));
  INV_X1    g231(.A(new_n387), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n386), .B1(new_n383), .B2(new_n256), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n396), .B2(new_n397), .ZN(new_n422));
  AND4_X1   g236(.A1(new_n403), .A2(new_n420), .A3(new_n392), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n398), .A2(KEYINPUT7), .A3(new_n401), .ZN(new_n424));
  AOI21_X1  g238(.A(G902), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n415), .A2(new_n416), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n416), .B1(new_n415), .B2(new_n425), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n363), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT9), .B(G234), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n429), .A2(new_n313), .A3(G953), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n191), .B2(G128), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n225), .A2(KEYINPUT86), .A3(G143), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n191), .A2(G128), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G134), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n213), .A3(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G122), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT14), .B1(new_n441), .B2(G116), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT14), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n238), .A3(G122), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n441), .A2(G116), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G107), .ZN(new_n448));
  XNOR2_X1  g262(.A(G116), .B(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n365), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(G107), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT87), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n440), .A2(new_n448), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT13), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n435), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n437), .A2(new_n455), .A3(G134), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n435), .B(new_n436), .C1(new_n454), .C2(new_n213), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n449), .B(new_n365), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n431), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT88), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n453), .A2(new_n459), .A3(new_n431), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n303), .A4(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G478), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(KEYINPUT15), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n303), .A3(new_n463), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT88), .ZN(new_n469));
  INV_X1    g283(.A(new_n466), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n467), .B1(new_n471), .B2(new_n464), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n475));
  OAI21_X1  g289(.A(G131), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n477));
  INV_X1    g291(.A(G237), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n342), .A3(G214), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n191), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n211), .A3(new_n473), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n476), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT83), .ZN(new_n483));
  OAI211_X1 g297(.A(KEYINPUT17), .B(G131), .C1(new_n474), .C2(new_n475), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n337), .A2(new_n323), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT83), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n476), .A2(new_n486), .A3(new_n477), .A4(new_n481), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G113), .B(G122), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n367), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n322), .A2(G146), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n325), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n480), .A2(new_n473), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT18), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(new_n211), .ZN(new_n495));
  OAI221_X1 g309(.A(new_n492), .B1(new_n493), .B2(new_n495), .C1(new_n476), .C2(new_n494), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n488), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n476), .A2(new_n481), .ZN(new_n498));
  OR2_X1    g312(.A1(KEYINPUT82), .A2(KEYINPUT19), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n324), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n324), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n498), .B(new_n323), .C1(new_n502), .C2(G146), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n496), .ZN(new_n504));
  INV_X1    g318(.A(new_n490), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT84), .A3(KEYINPUT20), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT84), .ZN(new_n511));
  INV_X1    g325(.A(new_n508), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n497), .B2(new_n506), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n508), .B(KEYINPUT85), .Z(new_n516));
  NAND3_X1  g330(.A1(new_n507), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(G234), .A2(G237), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n519), .A2(G952), .A3(new_n342), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  XOR2_X1   g335(.A(KEYINPUT21), .B(G898), .Z(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT89), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n519), .A2(G902), .A3(G953), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n521), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT90), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n488), .A2(new_n496), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n490), .ZN(new_n529));
  OAI21_X1  g343(.A(G475), .B1(new_n529), .B2(G902), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n472), .A2(new_n518), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n518), .A2(new_n530), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n534), .A2(KEYINPUT91), .A3(new_n527), .A4(new_n472), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n428), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n235), .A2(new_n220), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n199), .A2(new_n200), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n377), .A2(new_n373), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n386), .A2(new_n228), .A3(KEYINPUT10), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n376), .A2(new_n385), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n190), .B1(new_n192), .B2(new_n193), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n223), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n227), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n541), .B1(new_n545), .B2(KEYINPUT10), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n537), .B1(new_n540), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n373), .B(new_n377), .C1(new_n199), .C2(new_n200), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT64), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n195), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n191), .A2(KEYINPUT64), .A3(G146), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n221), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n225), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n227), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n386), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n537), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n549), .A2(new_n558), .A3(new_n559), .A4(new_n541), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n547), .A2(new_n548), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n342), .A2(G227), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT75), .ZN(new_n563));
  XNOR2_X1  g377(.A(G110), .B(G140), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(KEYINPUT77), .B(new_n537), .C1(new_n540), .C2(new_n546), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n561), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT78), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n386), .A2(new_n228), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n537), .B1(new_n570), .B2(new_n545), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(KEYINPUT12), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT12), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n556), .B1(new_n228), .B2(new_n386), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(new_n537), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n565), .A3(new_n560), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT78), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n561), .A2(new_n578), .A3(new_n566), .A4(new_n567), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G469), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n303), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n303), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n565), .B1(new_n576), .B2(new_n560), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n561), .A2(new_n567), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n565), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G469), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n582), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G221), .B1(new_n429), .B2(G902), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n536), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n312), .A2(KEYINPUT74), .A3(new_n359), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n362), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  NAND2_X1  g410(.A1(new_n284), .A2(new_n285), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n284), .A2(new_n303), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G472), .ZN(new_n599));
  AND4_X1   g413(.A1(new_n597), .A2(new_n589), .A3(new_n590), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n415), .A2(new_n425), .ZN(new_n601));
  INV_X1    g415(.A(new_n416), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT92), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n415), .A2(new_n416), .A3(new_n425), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT93), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n453), .A2(new_n607), .A3(new_n459), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n430), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT93), .B1(new_n430), .B2(new_n609), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n453), .B2(new_n459), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT33), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT95), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT95), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n615), .B(KEYINPUT33), .C1(new_n610), .C2(new_n612), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n461), .A2(new_n617), .A3(new_n463), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n465), .A2(G902), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n614), .A2(new_n616), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n468), .A2(new_n465), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n518), .A2(new_n530), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n415), .A2(KEYINPUT92), .A3(new_n416), .A4(new_n425), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n625), .A2(new_n363), .ZN(new_n626));
  AND4_X1   g440(.A1(new_n527), .A2(new_n606), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n600), .A2(new_n627), .A3(new_n359), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n606), .A2(new_n626), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n599), .A2(new_n597), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n359), .A2(new_n527), .ZN(new_n634));
  INV_X1    g448(.A(new_n472), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n507), .A2(new_n514), .A3(new_n508), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n510), .A2(new_n515), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n530), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n632), .A2(new_n591), .A3(new_n633), .A4(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n350), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT96), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n349), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n357), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n348), .A2(new_n355), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(new_n315), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n600), .A2(new_n536), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G110), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n649), .B(new_n651), .ZN(G12));
  AND3_X1   g466(.A1(new_n589), .A2(new_n590), .A3(new_n648), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n521), .B1(new_n525), .B2(G900), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n638), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n312), .A2(new_n653), .A3(new_n632), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  XOR2_X1   g472(.A(KEYINPUT98), .B(KEYINPUT39), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n654), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n591), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n661), .A2(KEYINPUT40), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(KEYINPUT40), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n426), .A2(new_n427), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT38), .ZN(new_n665));
  INV_X1    g479(.A(new_n288), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n300), .A2(new_n268), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n272), .B1(new_n276), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n310), .B1(new_n668), .B2(new_n303), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n666), .A2(new_n286), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n648), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n534), .A2(new_n472), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n672), .A3(new_n363), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n665), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n662), .A2(new_n663), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  NAND2_X1  g490(.A1(new_n624), .A2(new_n654), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n312), .A2(new_n653), .A3(new_n632), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  NAND2_X1  g494(.A1(new_n580), .A2(new_n303), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n581), .A2(KEYINPUT99), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n682), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n580), .A2(new_n303), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n590), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n627), .A2(new_n312), .A3(new_n359), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NOR2_X1   g504(.A1(new_n631), .A2(new_n686), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n312), .A3(new_n639), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  AOI21_X1  g507(.A(new_n671), .B1(new_n535), .B2(new_n533), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n312), .A2(new_n632), .A3(new_n694), .A4(new_n687), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  AND4_X1   g510(.A1(new_n527), .A2(new_n606), .A3(new_n672), .A4(new_n626), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n279), .A2(new_n280), .A3(new_n300), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n273), .B(new_n269), .C1(new_n276), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n285), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n271), .A2(new_n273), .B1(new_n282), .B2(new_n277), .ZN(new_n701));
  AOI21_X1  g515(.A(G902), .B1(new_n701), .B2(new_n275), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT100), .B(G472), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n359), .B(new_n700), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n686), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n697), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  OAI211_X1 g522(.A(new_n648), .B(new_n700), .C1(new_n702), .C2(new_n704), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT101), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n598), .A2(new_n703), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n711), .A2(new_n712), .A3(new_n648), .A4(new_n700), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n678), .A3(new_n691), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  INV_X1    g530(.A(new_n363), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n426), .A2(new_n427), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n585), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(G469), .B(new_n721), .C1(new_n587), .C2(new_n720), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n582), .A2(new_n722), .A3(new_n584), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n718), .A2(new_n723), .A3(new_n590), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n312), .A3(new_n359), .A4(new_n678), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n295), .A2(new_n293), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT71), .B1(new_n289), .B2(new_n265), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n291), .B(new_n266), .C1(new_n258), .C2(new_n268), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n305), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n302), .A2(KEYINPUT72), .A3(new_n303), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(G472), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n309), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n307), .A2(KEYINPUT73), .A3(G472), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n287), .A2(KEYINPUT103), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n286), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n738), .A2(new_n739), .A3(new_n288), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n677), .A2(new_n726), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n359), .A3(new_n724), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n727), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  AND4_X1   g560(.A1(new_n312), .A2(new_n724), .A3(new_n359), .A4(new_n656), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n213), .ZN(G36));
  OAI21_X1  g562(.A(G469), .B1(new_n587), .B2(KEYINPUT45), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(KEYINPUT45), .B(new_n721), .C1(new_n587), .C2(new_n720), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n583), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OR3_X1    g566(.A1(new_n752), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT104), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT105), .B1(new_n752), .B2(KEYINPUT46), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n582), .B1(new_n754), .B2(new_n755), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n590), .B(new_n660), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n718), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n534), .A2(new_n622), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT43), .Z(new_n764));
  NAND2_X1  g578(.A1(new_n599), .A2(new_n597), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n765), .A3(new_n648), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n761), .B(new_n768), .C1(new_n767), .C2(new_n766), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT106), .B(G137), .Z(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G39));
  OAI21_X1  g585(.A(new_n590), .B1(new_n758), .B2(new_n759), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT47), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT47), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n312), .A2(new_n359), .A3(new_n762), .A4(new_n677), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  AND2_X1   g591(.A1(new_n764), .A2(new_n520), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n717), .A3(new_n665), .ZN(new_n779));
  INV_X1    g593(.A(new_n706), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT50), .B1(new_n781), .B2(KEYINPUT112), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n779), .A2(KEYINPUT112), .A3(new_n780), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n783), .B1(new_n782), .B2(new_n784), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n762), .A2(new_n686), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n359), .A2(new_n792), .A3(new_n520), .A4(new_n670), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n622), .A2(new_n623), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n714), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n778), .A2(new_n792), .ZN(new_n797));
  INV_X1    g611(.A(new_n590), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n683), .A2(new_n685), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT107), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n773), .A2(new_n774), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n705), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n778), .A2(new_n802), .A3(new_n718), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT111), .ZN(new_n804));
  OAI221_X1 g618(.A(new_n795), .B1(new_n796), .B2(new_n797), .C1(new_n801), .C2(new_n804), .ZN(new_n805));
  OR3_X1    g619(.A1(new_n790), .A2(new_n791), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n791), .B1(new_n790), .B2(new_n805), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n359), .A2(new_n778), .A3(new_n742), .A4(new_n792), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT48), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n778), .A2(new_n691), .A3(new_n802), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n342), .A2(G952), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n793), .B2(new_n624), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(KEYINPUT48), .B2(new_n808), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n806), .A2(new_n807), .A3(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n590), .A2(new_n723), .A3(new_n671), .A4(new_n654), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n606), .A2(new_n672), .A3(new_n626), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n666), .A2(new_n286), .A3(new_n669), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n715), .A2(new_n657), .A3(new_n679), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT52), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n589), .A2(new_n590), .A3(new_n648), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n666), .A2(new_n286), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n738), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n824), .B(new_n632), .C1(new_n656), .C2(new_n678), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n715), .A4(new_n819), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n688), .A2(new_n649), .A3(new_n692), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n472), .A2(new_n530), .A3(new_n518), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n527), .B(new_n830), .C1(new_n534), .C2(new_n622), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n428), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n591), .A2(new_n832), .A3(new_n633), .A4(new_n359), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n695), .A2(new_n833), .A3(new_n707), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n747), .B1(new_n727), .B2(new_n744), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n677), .B1(new_n710), .B2(new_n713), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n472), .A2(new_n637), .A3(new_n530), .A4(new_n654), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n762), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n837), .A2(new_n724), .B1(new_n824), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n835), .A2(new_n836), .A3(new_n595), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT109), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n828), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n359), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n361), .B(new_n844), .C1(new_n738), .C2(new_n823), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT74), .B1(new_n312), .B2(new_n359), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n845), .A2(new_n846), .A3(new_n592), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n847), .A2(new_n829), .A3(new_n834), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(KEYINPUT109), .A3(new_n836), .A4(new_n840), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n843), .A2(KEYINPUT53), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT53), .B1(new_n843), .B2(new_n849), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g667(.A(KEYINPUT110), .B(KEYINPUT53), .C1(new_n843), .C2(new_n849), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT54), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n747), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n745), .A2(new_n856), .A3(new_n840), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n688), .A2(new_n649), .A3(new_n692), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n695), .A2(new_n833), .A3(new_n707), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n595), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n842), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n828), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n849), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n841), .A2(new_n828), .A3(new_n864), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n855), .A2(new_n869), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n815), .A2(new_n870), .B1(G952), .B2(G953), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n800), .B(KEYINPUT49), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n763), .A2(new_n844), .A3(new_n798), .A4(new_n717), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n872), .A2(new_n670), .A3(new_n665), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT108), .Z(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(G75));
  AOI21_X1  g690(.A(new_n303), .B1(new_n865), .B2(new_n868), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(G210), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n877), .B2(G210), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n394), .A2(new_n412), .A3(new_n414), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(new_n404), .Z(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT114), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT55), .Z(new_n885));
  AND3_X1   g699(.A1(new_n880), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n881), .B1(new_n880), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n342), .A2(G952), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G51));
  OAI21_X1  g703(.A(KEYINPUT54), .B1(new_n851), .B2(new_n867), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n869), .A3(KEYINPUT116), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n865), .A2(new_n868), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT54), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n583), .B(KEYINPUT57), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n580), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n750), .A2(new_n751), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT117), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n877), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n888), .B1(new_n897), .B2(new_n900), .ZN(G54));
  INV_X1    g715(.A(new_n888), .ZN(new_n902));
  AND2_X1   g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  OAI211_X1 g717(.A(G902), .B(new_n903), .C1(new_n851), .C2(new_n867), .ZN(new_n904));
  INV_X1    g718(.A(new_n507), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT119), .B1(new_n904), .B2(new_n905), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n902), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n904), .B2(new_n905), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n507), .A4(new_n903), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT120), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n906), .B(new_n907), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n918), .A3(new_n902), .A4(new_n914), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(G60));
  NAND3_X1  g734(.A1(new_n614), .A2(new_n616), .A3(new_n618), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n465), .A2(new_n303), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n922), .B1(new_n870), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n921), .A2(new_n925), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n891), .A2(new_n894), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n902), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT122), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n851), .A2(KEYINPUT54), .A3(new_n867), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n865), .A2(KEYINPUT110), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n851), .A2(new_n852), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n934), .A3(new_n850), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n932), .B1(new_n935), .B2(KEYINPUT54), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n921), .B1(new_n936), .B2(new_n925), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n937), .A2(new_n938), .A3(new_n902), .A4(new_n929), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n931), .A2(new_n939), .ZN(G63));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT60), .Z(new_n942));
  NAND3_X1  g756(.A1(new_n892), .A2(new_n645), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n892), .A2(new_n942), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n902), .B(new_n943), .C1(new_n944), .C2(new_n347), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g760(.A(new_n342), .B1(new_n523), .B2(G224), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n860), .B2(new_n342), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT123), .Z(new_n949));
  INV_X1    g763(.A(G898), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n882), .B1(new_n950), .B2(G953), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n949), .B(new_n951), .ZN(G69));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n675), .B1(KEYINPUT124), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n825), .A2(new_n715), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n953), .A2(KEYINPUT124), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(new_n958));
  OAI21_X1  g772(.A(new_n830), .B1(new_n534), .B2(new_n622), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n661), .A2(new_n762), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n362), .A3(new_n594), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n776), .A2(new_n769), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n342), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n231), .A2(new_n237), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(new_n502), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(G900), .B2(G953), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n742), .A2(new_n359), .A3(new_n817), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n955), .B1(new_n761), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n776), .A2(new_n769), .A3(new_n836), .A4(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n967), .B1(new_n970), .B2(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n342), .B1(G227), .B2(G900), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT125), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n973), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n972), .B(new_n975), .Z(G72));
  NOR3_X1   g790(.A1(new_n958), .A2(new_n860), .A3(new_n962), .ZN(new_n977));
  NAND2_X1  g791(.A1(G472), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT127), .ZN(new_n979));
  XNOR2_X1  g793(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n266), .B(new_n289), .C1(new_n977), .C2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n970), .A2(new_n860), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(new_n981), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n258), .A2(new_n265), .A3(new_n268), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n982), .B(new_n902), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n729), .A2(new_n730), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n981), .B1(new_n987), .B2(new_n272), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n935), .B2(new_n988), .ZN(G57));
endmodule


