//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n577, new_n578, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT64), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT67), .B1(new_n464), .B2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(new_n462), .A3(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n463), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n473), .B1(G2105), .B2(new_n479), .ZN(G160));
  XNOR2_X1  g055(.A(new_n477), .B(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n462), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(KEYINPUT70), .A3(new_n462), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n481), .A2(G2105), .ZN(new_n488));
  MUX2_X1   g063(.A(G100), .B(G112), .S(G2105), .Z(new_n489));
  AOI22_X1  g064(.A1(new_n488), .A2(G124), .B1(G2104), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n487), .A2(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n475), .B2(new_n476), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n461), .A2(new_n495), .A3(new_n497), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n493), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  MUX2_X1   g076(.A(G102), .B(G114), .S(G2105), .Z(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2104), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n501), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(G543), .B1(new_n513), .B2(new_n512), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT72), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n521), .B1(new_n509), .B2(new_n510), .ZN(new_n522));
  OAI21_X1  g097(.A(G651), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g100(.A(KEYINPUT73), .B(G651), .C1(new_n520), .C2(new_n522), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n518), .B1(new_n525), .B2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT76), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n509), .A2(new_n510), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n513), .A2(new_n512), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT77), .B(G89), .Z(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n511), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n516), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT74), .B(G51), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n532), .A2(new_n542), .ZN(G168));
  XNOR2_X1  g118(.A(KEYINPUT78), .B(G90), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n514), .A2(new_n544), .B1(new_n516), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G651), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n514), .A2(new_n551), .B1(new_n516), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n548), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT79), .Z(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G53), .ZN(new_n566));
  OR3_X1    g141(.A1(new_n516), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n564), .B1(new_n516), .B2(new_n566), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n533), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n535), .B2(G91), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G299));
  OR2_X1    g149(.A1(new_n546), .A2(new_n549), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  NAND2_X1  g151(.A1(new_n525), .A2(new_n526), .ZN(new_n577));
  INV_X1    g152(.A(new_n518), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G303));
  NAND2_X1  g154(.A1(new_n535), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n539), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  INV_X1    g159(.A(G48), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n514), .A2(new_n584), .B1(new_n516), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n548), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n548), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT81), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n594));
  XOR2_X1   g169(.A(KEYINPUT82), .B(G47), .Z(new_n595));
  AOI22_X1  g170(.A1(new_n535), .A2(G85), .B1(new_n539), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n592), .A2(KEYINPUT81), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n599));
  NOR3_X1   g174(.A1(new_n591), .A2(new_n599), .A3(new_n548), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT83), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n597), .A2(new_n602), .ZN(G290));
  XOR2_X1   g178(.A(KEYINPUT84), .B(KEYINPUT10), .Z(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n535), .A2(G92), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n604), .B1(new_n514), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n533), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(new_n539), .B2(G54), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  MUX2_X1   g190(.A(G301), .B(new_n614), .S(new_n615), .Z(G284));
  MUX2_X1   g191(.A(G301), .B(new_n614), .S(new_n615), .Z(G321));
  NOR2_X1   g192(.A1(G299), .A2(G868), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g194(.A(new_n618), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g195(.A(new_n614), .ZN(new_n621));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G860), .ZN(G148));
  INV_X1    g198(.A(new_n556), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n614), .A2(G559), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G868), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n465), .A2(new_n467), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(new_n477), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT85), .B(G2100), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n486), .A2(G135), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  MUX2_X1   g211(.A(G99), .B(G111), .S(G2105), .Z(new_n637));
  AOI22_X1  g212(.A1(new_n488), .A2(G123), .B1(G2104), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n639), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2427), .ZN(new_n646));
  INV_X1    g221(.A(G2430), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT86), .Z(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  INV_X1    g241(.A(new_n662), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n663), .B1(new_n669), .B2(new_n660), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n661), .B2(new_n668), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n661), .A2(new_n664), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n667), .B1(new_n672), .B2(KEYINPUT17), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n666), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(new_n636), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2100), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT87), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT89), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT88), .ZN(new_n693));
  XOR2_X1   g268(.A(G1981), .B(G1986), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  NOR2_X1   g272(.A1(G6), .A2(G16), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n589), .B2(G16), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT91), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT92), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n703), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G22), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G166), .B2(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G1971), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G23), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT93), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(G288), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT33), .B(G1976), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT94), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G1971), .ZN(new_n716));
  INV_X1    g291(.A(new_n707), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n704), .A2(new_n705), .A3(new_n708), .A4(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n486), .A2(G131), .ZN(new_n724));
  MUX2_X1   g299(.A(G95), .B(G107), .S(G2105), .Z(new_n725));
  AOI22_X1  g300(.A1(new_n488), .A2(G119), .B1(G2104), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT90), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n723), .B1(new_n728), .B2(new_n722), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT35), .B(G1991), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G16), .A2(G24), .ZN(new_n732));
  INV_X1    g307(.A(G290), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(G1986), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n720), .A2(new_n721), .A3(new_n731), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT36), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G162), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2090), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n711), .A2(G20), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT23), .Z(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G299), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT31), .B(G11), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT30), .B(G28), .Z(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n711), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n711), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n749), .B1(new_n751), .B2(G1961), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n746), .B(new_n752), .C1(G1961), .C2(new_n751), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n711), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n711), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT96), .B(G1966), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G19), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n556), .B2(G16), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1341), .Z(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n760), .C1(new_n722), .C2(new_n640), .ZN(new_n761));
  NOR2_X1   g336(.A1(G4), .A2(G16), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n621), .B2(G16), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G27), .A2(G29), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G164), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2078), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(G160), .A2(G29), .ZN(new_n771));
  AND2_X1   g346(.A1(KEYINPUT24), .A2(G34), .ZN(new_n772));
  NOR2_X1   g347(.A1(KEYINPUT24), .A2(G34), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n722), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2084), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  OR4_X1    g352(.A1(new_n753), .A2(new_n761), .A3(new_n770), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n722), .A2(G26), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT28), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n488), .A2(G128), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT95), .ZN(new_n782));
  MUX2_X1   g357(.A(G104), .B(G116), .S(G2105), .Z(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(G2104), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n486), .A2(G140), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n780), .B1(new_n786), .B2(G29), .ZN(new_n787));
  INV_X1    g362(.A(G2067), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n722), .A2(G33), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n486), .A2(G139), .ZN(new_n791));
  NAND2_X1  g366(.A1(G115), .A2(G2104), .ZN(new_n792));
  INV_X1    g367(.A(G127), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n477), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n794), .A2(G2105), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n790), .B1(new_n800), .B2(new_n722), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G2072), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n486), .A2(G141), .ZN(new_n803));
  NAND3_X1  g378(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT26), .Z(new_n805));
  INV_X1    g380(.A(G105), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n629), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n488), .B2(G129), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G32), .B(new_n809), .S(G29), .Z(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT27), .B(G1996), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n802), .A2(new_n812), .ZN(new_n813));
  NOR4_X1   g388(.A1(new_n742), .A2(new_n778), .A3(new_n789), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n738), .A2(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  AOI22_X1  g391(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(new_n548), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n535), .A2(G93), .B1(G55), .B2(new_n539), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n556), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(KEYINPUT97), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n817), .A2(new_n823), .A3(new_n548), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n624), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n621), .A2(G559), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT98), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n832), .A2(new_n833), .A3(G860), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n825), .A2(G860), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(new_n800), .B(new_n809), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n499), .A2(new_n500), .ZN(new_n839));
  INV_X1    g414(.A(new_n493), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n505), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n786), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(G164), .B1(new_n784), .B2(new_n785), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n486), .A2(G142), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n488), .A2(G130), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT100), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n462), .A2(G106), .ZN(new_n851));
  NAND2_X1  g426(.A1(G118), .A2(G2105), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n464), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n848), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n727), .B(new_n631), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n846), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n846), .B1(new_n857), .B2(new_n856), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n838), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G162), .B(G160), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n640), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n856), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n845), .B2(new_n844), .ZN(new_n866));
  INV_X1    g441(.A(new_n838), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n858), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n864), .B1(new_n861), .B2(new_n868), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(G395));
  NOR2_X1   g450(.A1(new_n825), .A2(G868), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  INV_X1    g452(.A(G288), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n594), .B1(new_n593), .B2(new_n596), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n601), .A2(KEYINPUT83), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G305), .B(G166), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n597), .A2(new_n602), .A3(G288), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT104), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n881), .A2(new_n883), .A3(new_n887), .A4(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n883), .B1(new_n881), .B2(new_n884), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n877), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g467(.A(KEYINPUT105), .B(new_n890), .C1(new_n886), .C2(new_n888), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT42), .B1(new_n889), .B2(new_n891), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n827), .B(new_n626), .ZN(new_n899));
  NAND2_X1  g474(.A1(G299), .A2(new_n614), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n569), .A2(new_n609), .A3(new_n573), .A4(new_n613), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(KEYINPUT102), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(KEYINPUT102), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n900), .A2(new_n907), .A3(new_n901), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT103), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n900), .A2(new_n910), .A3(new_n907), .A4(new_n901), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n902), .A2(KEYINPUT41), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n899), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n905), .A2(new_n906), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n898), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n896), .B2(new_n897), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n876), .B1(new_n920), .B2(G868), .ZN(G331));
  NAND2_X1  g496(.A1(G331), .A2(KEYINPUT106), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n615), .B1(new_n917), .B2(new_n919), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n876), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(G295));
  OAI21_X1  g501(.A(G301), .B1(new_n532), .B2(new_n542), .ZN(new_n927));
  NAND4_X1  g502(.A1(G171), .A2(new_n531), .A3(new_n541), .A4(new_n538), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(new_n821), .B2(new_n826), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n819), .A2(new_n556), .A3(new_n820), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n825), .A2(new_n624), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n927), .A4(new_n928), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n903), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n931), .A2(new_n932), .B1(new_n927), .B2(new_n928), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n930), .A2(KEYINPUT107), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n913), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT108), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n942), .B(new_n913), .C1(new_n938), .C2(new_n939), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n935), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n889), .A2(new_n891), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT105), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n889), .A2(new_n877), .A3(new_n891), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n930), .A2(KEYINPUT107), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n936), .A2(new_n937), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n933), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n902), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n930), .A2(new_n933), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n912), .A2(new_n908), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n948), .B(new_n870), .C1(new_n894), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n894), .B2(new_n944), .ZN(new_n959));
  INV_X1    g534(.A(new_n943), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n942), .B1(new_n951), .B2(new_n913), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n934), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n892), .B2(new_n893), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT109), .B1(new_n965), .B2(KEYINPUT44), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n958), .A2(new_n967), .A3(new_n964), .A4(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n963), .A2(new_n948), .A3(new_n957), .A4(new_n870), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n959), .A2(KEYINPUT110), .A3(new_n957), .A4(new_n963), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n968), .B1(new_n956), .B2(KEYINPUT43), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n974), .B2(new_n976), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n966), .B(new_n969), .C1(new_n977), .C2(new_n978), .ZN(G397));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n501), .B2(new_n505), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n479), .A2(G2105), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n470), .A2(G40), .A3(new_n984), .A4(new_n472), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n786), .A2(G2067), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n784), .A2(new_n788), .A3(new_n785), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n809), .B(G1996), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n727), .B(new_n730), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(G290), .B(G1986), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n986), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n589), .B(G1981), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT49), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n981), .A2(new_n998), .ZN(new_n999));
  AND4_X1   g574(.A1(G40), .A2(new_n470), .A3(new_n984), .A4(new_n472), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT112), .B(new_n980), .C1(new_n501), .C2(new_n505), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(KEYINPUT49), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n997), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n878), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(G1981), .B2(G305), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n1003), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1002), .A2(G8), .A3(new_n1006), .A4(G288), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT114), .B1(new_n878), .B2(G1976), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1002), .A2(G8), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1003), .A2(new_n1010), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n1005), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n843), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n1000), .ZN(new_n1019));
  INV_X1    g594(.A(new_n983), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n716), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n999), .A2(new_n1022), .A3(new_n1001), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n985), .B1(KEYINPUT50), .B2(new_n981), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(G2090), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  NOR3_X1   g604(.A1(G166), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT113), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1028), .B1(G166), .B2(new_n1029), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1026), .A2(new_n1036), .A3(G8), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1009), .B1(new_n1017), .B2(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1015), .A2(new_n1016), .A3(new_n1005), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n843), .A2(KEYINPUT115), .A3(new_n1022), .A4(new_n980), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n985), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n999), .A2(new_n1001), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT50), .ZN(new_n1046));
  INV_X1    g621(.A(G2090), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1048), .A2(new_n1021), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1040), .B1(new_n1049), .B2(new_n1029), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n999), .B2(new_n1001), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n756), .B1(new_n1051), .B2(new_n1019), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1023), .A2(new_n776), .A3(new_n1024), .ZN(new_n1053));
  AOI211_X1 g628(.A(new_n1029), .B(G286), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1039), .A2(new_n1050), .A3(new_n1037), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT116), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT63), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1026), .A2(new_n1036), .A3(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1017), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1050), .A4(new_n1054), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n1027), .B(new_n1030), .C1(new_n1026), .C2(G8), .ZN(new_n1063));
  OR3_X1    g638(.A1(new_n1063), .A2(new_n1017), .A3(KEYINPUT117), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1037), .A2(new_n1054), .A3(KEYINPUT63), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT117), .B1(new_n1063), .B2(new_n1017), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1038), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G299), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n569), .A2(KEYINPUT118), .A3(new_n1071), .A4(new_n573), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n981), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n985), .B1(new_n1075), .B2(KEYINPUT45), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n983), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT56), .B(G2072), .Z(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1081));
  INV_X1    g656(.A(G1956), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1956), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT121), .B1(new_n1086), .B2(new_n1079), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1074), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1025), .A2(KEYINPUT119), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1023), .A2(new_n1090), .A3(new_n1024), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n764), .A3(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1002), .A2(G2067), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1092), .A2(KEYINPUT120), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT120), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1086), .A2(new_n1079), .A3(new_n1073), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n614), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1088), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT60), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1023), .A2(new_n1090), .A3(new_n1024), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1090), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1105), .A2(new_n1106), .A3(G1348), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1104), .B1(new_n1107), .B2(new_n1093), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1092), .A2(KEYINPUT120), .A3(new_n1094), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n614), .B1(new_n1110), .B2(KEYINPUT60), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1102), .B(new_n621), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1103), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1074), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n1115), .B2(new_n1098), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  INV_X1    g692(.A(G1996), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1076), .A2(new_n1118), .A3(new_n983), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1002), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n624), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1117), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1122), .B2(KEYINPUT123), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1123), .B(new_n1117), .C1(new_n1122), .C2(KEYINPUT123), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1116), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1098), .A2(new_n1114), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(new_n1088), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1101), .B1(new_n1113), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1059), .A2(new_n1050), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1134));
  OAI21_X1  g709(.A(G8), .B1(new_n1134), .B2(G286), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT51), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1134), .B2(G286), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1105), .A2(new_n1106), .A3(G1961), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1077), .A2(G2078), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1141), .A2(KEYINPUT53), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1051), .A2(new_n1019), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(KEYINPUT53), .A3(new_n768), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(G171), .B(KEYINPUT54), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n768), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n479), .B(KEYINPUT124), .Z(new_n1151));
  AOI211_X1 g726(.A(new_n1150), .B(new_n473), .C1(new_n1151), .C2(G2105), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n983), .A3(new_n1018), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1143), .A2(new_n1147), .A3(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1133), .A2(new_n1139), .A3(new_n1149), .A4(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT125), .B(new_n1068), .C1(new_n1132), .C2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1139), .B(KEYINPUT62), .Z(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(G171), .A3(new_n1133), .A4(new_n1146), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1110), .A2(KEYINPUT60), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT60), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n621), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1110), .A2(KEYINPUT60), .A3(new_n614), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1160), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g739(.A(new_n1116), .B1(new_n1126), .B2(new_n1127), .C1(new_n1129), .C2(new_n1088), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1100), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1155), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT125), .B1(new_n1168), .B2(new_n1068), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n995), .B1(new_n1159), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n986), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n728), .A2(new_n730), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1172), .A2(KEYINPUT126), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(KEYINPUT126), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n991), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1171), .B1(new_n1175), .B2(new_n988), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n986), .B1(new_n989), .B2(new_n809), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n986), .A2(new_n1118), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT46), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n993), .A2(new_n986), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n733), .A2(new_n735), .A3(new_n986), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT48), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1176), .B(new_n1182), .C1(new_n1183), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1170), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(G319), .ZN(new_n1189));
  NOR3_X1   g763(.A1(G401), .A2(new_n1189), .A3(G227), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n696), .A2(new_n1190), .ZN(new_n1191));
  NOR3_X1   g765(.A1(new_n873), .A2(new_n1191), .A3(new_n965), .ZN(G308));
  INV_X1    g766(.A(G308), .ZN(G225));
endmodule


