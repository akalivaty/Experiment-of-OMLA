

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n593), .A2(n592), .ZN(G164) );
  NOR2_X2 U554 ( .A1(n725), .A2(n724), .ZN(n738) );
  AND2_X1 U555 ( .A1(G160), .A2(G40), .ZN(n649) );
  NOR2_X4 U556 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  BUF_X4 U557 ( .A(n1006), .Z(n521) );
  NOR2_X1 U558 ( .A1(n945), .A2(n654), .ZN(n655) );
  NAND2_X2 U559 ( .A1(n649), .A2(n648), .ZN(n693) );
  NAND2_X1 U560 ( .A1(G8), .A2(n693), .ZN(n720) );
  INV_X1 U561 ( .A(G2105), .ZN(n525) );
  NOR2_X1 U562 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X2 U563 ( .A(n532), .B(KEYINPUT65), .ZN(G160) );
  XNOR2_X1 U564 ( .A(n662), .B(KEYINPUT27), .ZN(n663) );
  XNOR2_X1 U565 ( .A(n664), .B(n663), .ZN(n666) );
  INV_X1 U566 ( .A(n693), .ZN(n676) );
  INV_X1 U567 ( .A(KEYINPUT28), .ZN(n670) );
  XNOR2_X1 U568 ( .A(n684), .B(KEYINPUT30), .ZN(n685) );
  NOR2_X1 U569 ( .A1(G1966), .A2(n720), .ZN(n682) );
  INV_X1 U570 ( .A(n956), .ZN(n722) );
  NAND2_X1 U571 ( .A1(n723), .A2(n722), .ZN(n724) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n523) );
  NOR2_X1 U573 ( .A1(G651), .A2(n567), .ZN(n793) );
  NOR2_X1 U574 ( .A1(G651), .A2(G543), .ZN(n790) );
  AND2_X4 U575 ( .A1(n525), .A2(G2104), .ZN(n1005) );
  NAND2_X1 U576 ( .A1(G101), .A2(n1005), .ZN(n522) );
  XNOR2_X1 U577 ( .A(KEYINPUT23), .B(n522), .ZN(n529) );
  XNOR2_X2 U578 ( .A(n524), .B(n523), .ZN(n1006) );
  NAND2_X1 U579 ( .A1(G137), .A2(n1006), .ZN(n527) );
  NOR2_X1 U580 ( .A1(G2104), .A2(n525), .ZN(n601) );
  NAND2_X1 U581 ( .A1(G125), .A2(n601), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U583 ( .A1(n529), .A2(n528), .ZN(n531) );
  AND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n1002) );
  NAND2_X1 U585 ( .A1(n1002), .A2(G113), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n567) );
  INV_X1 U588 ( .A(G651), .ZN(n537) );
  NOR2_X1 U589 ( .A1(n567), .A2(n537), .ZN(n789) );
  NAND2_X1 U590 ( .A1(n789), .A2(G78), .ZN(n533) );
  XNOR2_X1 U591 ( .A(n533), .B(KEYINPUT66), .ZN(n535) );
  NAND2_X1 U592 ( .A1(G91), .A2(n790), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U594 ( .A(KEYINPUT67), .B(n536), .ZN(n542) );
  NOR2_X1 U595 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n538), .Z(n795) );
  NAND2_X1 U597 ( .A1(G65), .A2(n795), .ZN(n540) );
  NAND2_X1 U598 ( .A1(G53), .A2(n793), .ZN(n539) );
  AND2_X1 U599 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n542), .A2(n541), .ZN(G299) );
  NAND2_X1 U601 ( .A1(G64), .A2(n795), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G52), .A2(n793), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G77), .A2(n789), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G90), .A2(n790), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U608 ( .A1(n549), .A2(n548), .ZN(G171) );
  NAND2_X1 U609 ( .A1(G89), .A2(n790), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n550), .B(KEYINPUT74), .ZN(n551) );
  XNOR2_X1 U611 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G76), .A2(n789), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U614 ( .A(n554), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G63), .A2(n795), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G51), .A2(n793), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U618 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U620 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U621 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U622 ( .A1(G75), .A2(n789), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G88), .A2(n790), .ZN(n561) );
  NAND2_X1 U624 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U625 ( .A1(G62), .A2(n795), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G50), .A2(n793), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U628 ( .A1(n566), .A2(n565), .ZN(G166) );
  INV_X1 U629 ( .A(G166), .ZN(G303) );
  NAND2_X1 U630 ( .A1(G651), .A2(G74), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G49), .A2(n793), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G87), .A2(n567), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n795), .A2(n570), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT77), .B(n573), .Z(G288) );
  NAND2_X1 U637 ( .A1(G61), .A2(n795), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G48), .A2(n793), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n789), .A2(G73), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT2), .B(n576), .Z(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n790), .A2(G86), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(G305) );
  NAND2_X1 U645 ( .A1(G60), .A2(n795), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G47), .A2(n793), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G72), .A2(n789), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G85), .A2(n790), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  OR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(G290) );
  AND2_X1 U652 ( .A1(G138), .A2(n521), .ZN(n587) );
  XNOR2_X1 U653 ( .A(KEYINPUT81), .B(n587), .ZN(n593) );
  NAND2_X1 U654 ( .A1(n1002), .A2(G114), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G102), .A2(n1005), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G126), .A2(n601), .ZN(n588) );
  AND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U659 ( .A1(G164), .A2(G1384), .ZN(n648) );
  NAND2_X1 U660 ( .A1(G160), .A2(G40), .ZN(n594) );
  NOR2_X1 U661 ( .A1(n648), .A2(n594), .ZN(n595) );
  XNOR2_X1 U662 ( .A(KEYINPUT83), .B(n595), .ZN(n627) );
  INV_X1 U663 ( .A(n627), .ZN(n758) );
  XNOR2_X1 U664 ( .A(G2067), .B(KEYINPUT37), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT84), .ZN(n753) );
  NAND2_X1 U666 ( .A1(G104), .A2(n1005), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G140), .A2(n521), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n600) );
  XOR2_X1 U669 ( .A(KEYINPUT85), .B(KEYINPUT34), .Z(n599) );
  XNOR2_X1 U670 ( .A(n600), .B(n599), .ZN(n606) );
  BUF_X1 U671 ( .A(n601), .Z(n1001) );
  NAND2_X1 U672 ( .A1(G128), .A2(n1001), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G116), .A2(n1002), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U675 ( .A(KEYINPUT35), .B(n604), .Z(n605) );
  NOR2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U677 ( .A(KEYINPUT36), .B(n607), .ZN(n992) );
  NOR2_X1 U678 ( .A1(n753), .A2(n992), .ZN(n916) );
  NAND2_X1 U679 ( .A1(n758), .A2(n916), .ZN(n756) );
  NAND2_X1 U680 ( .A1(G95), .A2(n1005), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G131), .A2(n521), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U683 ( .A(KEYINPUT86), .B(n610), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G119), .A2(n1001), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G107), .A2(n1002), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n1012) );
  INV_X1 U688 ( .A(G1991), .ZN(n879) );
  NOR2_X1 U689 ( .A1(n1012), .A2(n879), .ZN(n626) );
  NAND2_X1 U690 ( .A1(G129), .A2(n1001), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G117), .A2(n1002), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT87), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G141), .A2(n521), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n623) );
  XOR2_X1 U696 ( .A(KEYINPUT88), .B(KEYINPUT38), .Z(n621) );
  NAND2_X1 U697 ( .A1(G105), .A2(n1005), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n624), .B(KEYINPUT89), .ZN(n745) );
  INV_X1 U701 ( .A(n745), .ZN(n1017) );
  INV_X1 U702 ( .A(G1996), .ZN(n650) );
  NOR2_X1 U703 ( .A1(n1017), .A2(n650), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n906) );
  NOR2_X1 U705 ( .A1(n906), .A2(n627), .ZN(n749) );
  INV_X1 U706 ( .A(n749), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n756), .A2(n628), .ZN(n740) );
  NAND2_X1 U708 ( .A1(G66), .A2(n795), .ZN(n630) );
  NAND2_X1 U709 ( .A1(G54), .A2(n793), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G79), .A2(n789), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G92), .A2(n790), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U715 ( .A(KEYINPUT15), .B(n635), .Z(n1023) );
  NAND2_X1 U716 ( .A1(n795), .A2(G56), .ZN(n636) );
  XNOR2_X1 U717 ( .A(KEYINPUT14), .B(n636), .ZN(n647) );
  NAND2_X1 U718 ( .A1(G43), .A2(n793), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n637), .B(KEYINPUT73), .ZN(n645) );
  NAND2_X1 U720 ( .A1(G68), .A2(n789), .ZN(n641) );
  XOR2_X1 U721 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n639) );
  NAND2_X1 U722 ( .A1(G81), .A2(n790), .ZN(n638) );
  XNOR2_X1 U723 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U725 ( .A(n642), .B(KEYINPUT13), .ZN(n643) );
  XOR2_X1 U726 ( .A(n643), .B(KEYINPUT72), .Z(n644) );
  NOR2_X1 U727 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n945) );
  NOR2_X2 U729 ( .A1(n693), .A2(n650), .ZN(n651) );
  XOR2_X1 U730 ( .A(n651), .B(KEYINPUT26), .Z(n653) );
  NAND2_X1 U731 ( .A1(n693), .A2(G1341), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n654) );
  OR2_X1 U733 ( .A1(n1023), .A2(n655), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n1023), .A2(n655), .ZN(n659) );
  NAND2_X1 U735 ( .A1(G1348), .A2(n693), .ZN(n657) );
  NAND2_X1 U736 ( .A1(n676), .A2(G2067), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n668) );
  NAND2_X1 U740 ( .A1(G2072), .A2(n676), .ZN(n664) );
  INV_X1 U741 ( .A(KEYINPUT93), .ZN(n662) );
  INV_X1 U742 ( .A(G1956), .ZN(n859) );
  NOR2_X1 U743 ( .A1(n676), .A2(n859), .ZN(n665) );
  NOR2_X1 U744 ( .A1(n666), .A2(n665), .ZN(n669) );
  INV_X1 U745 ( .A(G299), .ZN(n954) );
  NAND2_X1 U746 ( .A1(n669), .A2(n954), .ZN(n667) );
  NAND2_X1 U747 ( .A1(n668), .A2(n667), .ZN(n673) );
  NOR2_X1 U748 ( .A1(n669), .A2(n954), .ZN(n671) );
  XNOR2_X1 U749 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U750 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U751 ( .A(KEYINPUT29), .B(n674), .Z(n681) );
  NAND2_X1 U752 ( .A1(G1961), .A2(n693), .ZN(n678) );
  XNOR2_X1 U753 ( .A(G2078), .B(KEYINPUT25), .ZN(n675) );
  XNOR2_X1 U754 ( .A(n675), .B(KEYINPUT91), .ZN(n885) );
  NAND2_X1 U755 ( .A1(n676), .A2(n885), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U757 ( .A(KEYINPUT92), .B(n679), .Z(n686) );
  NAND2_X1 U758 ( .A1(G171), .A2(n686), .ZN(n680) );
  NAND2_X1 U759 ( .A1(n681), .A2(n680), .ZN(n691) );
  XOR2_X1 U760 ( .A(KEYINPUT90), .B(n682), .Z(n705) );
  INV_X1 U761 ( .A(G8), .ZN(n698) );
  NOR2_X1 U762 ( .A1(G2084), .A2(n693), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n698), .A2(n703), .ZN(n683) );
  NAND2_X1 U764 ( .A1(n705), .A2(n683), .ZN(n684) );
  NOR2_X1 U765 ( .A1(G168), .A2(n685), .ZN(n688) );
  NOR2_X1 U766 ( .A1(G171), .A2(n686), .ZN(n687) );
  NOR2_X1 U767 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U768 ( .A(KEYINPUT31), .B(n689), .Z(n690) );
  NAND2_X1 U769 ( .A1(n691), .A2(n690), .ZN(n702) );
  AND2_X1 U770 ( .A1(G286), .A2(G8), .ZN(n692) );
  NAND2_X1 U771 ( .A1(n702), .A2(n692), .ZN(n700) );
  NOR2_X1 U772 ( .A1(G1971), .A2(n720), .ZN(n695) );
  NOR2_X1 U773 ( .A1(G2090), .A2(n693), .ZN(n694) );
  NOR2_X1 U774 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U775 ( .A1(n696), .A2(G303), .ZN(n697) );
  OR2_X1 U776 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U777 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U778 ( .A(n701), .B(KEYINPUT32), .ZN(n728) );
  INV_X1 U779 ( .A(n702), .ZN(n707) );
  NAND2_X1 U780 ( .A1(G8), .A2(n703), .ZN(n704) );
  NAND2_X1 U781 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U782 ( .A1(n707), .A2(n706), .ZN(n729) );
  INV_X1 U783 ( .A(n729), .ZN(n708) );
  NAND2_X1 U784 ( .A1(G1976), .A2(G288), .ZN(n940) );
  NAND2_X1 U785 ( .A1(n708), .A2(n940), .ZN(n709) );
  NOR2_X1 U786 ( .A1(n728), .A2(n709), .ZN(n714) );
  INV_X1 U787 ( .A(n940), .ZN(n712) );
  NOR2_X1 U788 ( .A1(G1976), .A2(G288), .ZN(n943) );
  NOR2_X1 U789 ( .A1(G1971), .A2(G303), .ZN(n710) );
  NOR2_X1 U790 ( .A1(n943), .A2(n710), .ZN(n711) );
  NOR2_X1 U791 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U792 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U793 ( .A1(n715), .A2(n720), .ZN(n716) );
  XNOR2_X1 U794 ( .A(n716), .B(KEYINPUT64), .ZN(n717) );
  NOR2_X1 U795 ( .A1(KEYINPUT33), .A2(n717), .ZN(n718) );
  XNOR2_X1 U796 ( .A(n718), .B(KEYINPUT94), .ZN(n725) );
  NAND2_X1 U797 ( .A1(n943), .A2(KEYINPUT33), .ZN(n719) );
  XNOR2_X1 U798 ( .A(KEYINPUT95), .B(n719), .ZN(n721) );
  INV_X1 U799 ( .A(n720), .ZN(n733) );
  NAND2_X1 U800 ( .A1(n721), .A2(n733), .ZN(n723) );
  XNOR2_X1 U801 ( .A(G1981), .B(G305), .ZN(n956) );
  NOR2_X1 U802 ( .A1(G1981), .A2(G305), .ZN(n726) );
  XNOR2_X1 U803 ( .A(n726), .B(KEYINPUT24), .ZN(n727) );
  NAND2_X1 U804 ( .A1(n727), .A2(n733), .ZN(n736) );
  NOR2_X1 U805 ( .A1(n728), .A2(n729), .ZN(n732) );
  NAND2_X1 U806 ( .A1(G8), .A2(G166), .ZN(n730) );
  NOR2_X1 U807 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U808 ( .A1(n732), .A2(n731), .ZN(n734) );
  OR2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U811 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U812 ( .A(n741), .B(KEYINPUT96), .ZN(n744) );
  XNOR2_X1 U813 ( .A(KEYINPUT82), .B(G1986), .ZN(n742) );
  XNOR2_X1 U814 ( .A(n742), .B(G290), .ZN(n951) );
  NAND2_X1 U815 ( .A1(n951), .A2(n758), .ZN(n743) );
  NAND2_X1 U816 ( .A1(n744), .A2(n743), .ZN(n762) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n745), .ZN(n909) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n746) );
  AND2_X1 U819 ( .A1(n879), .A2(n1012), .ZN(n905) );
  NOR2_X1 U820 ( .A1(n746), .A2(n905), .ZN(n747) );
  XOR2_X1 U821 ( .A(KEYINPUT97), .B(n747), .Z(n748) );
  NOR2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U823 ( .A1(n909), .A2(n750), .ZN(n751) );
  XOR2_X1 U824 ( .A(KEYINPUT39), .B(n751), .Z(n752) );
  XNOR2_X1 U825 ( .A(n752), .B(KEYINPUT98), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n753), .A2(n992), .ZN(n918) );
  NAND2_X1 U827 ( .A1(n754), .A2(n918), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U829 ( .A(KEYINPUT99), .B(n757), .ZN(n759) );
  NAND2_X1 U830 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U831 ( .A(n760), .B(KEYINPUT100), .ZN(n761) );
  NAND2_X1 U832 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U833 ( .A(n763), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U834 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U835 ( .A(G82), .ZN(G220) );
  INV_X1 U836 ( .A(G57), .ZN(G237) );
  INV_X1 U837 ( .A(G120), .ZN(G236) );
  XOR2_X1 U838 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n766) );
  NAND2_X1 U839 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U840 ( .A(n766), .B(n765), .ZN(G223) );
  XOR2_X1 U841 ( .A(G223), .B(KEYINPUT70), .Z(n837) );
  NAND2_X1 U842 ( .A1(n837), .A2(G567), .ZN(n767) );
  XOR2_X1 U843 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  INV_X1 U844 ( .A(G860), .ZN(n772) );
  OR2_X1 U845 ( .A1(n945), .A2(n772), .ZN(G153) );
  INV_X1 U846 ( .A(G171), .ZN(G301) );
  NAND2_X1 U847 ( .A1(G868), .A2(G301), .ZN(n769) );
  OR2_X1 U848 ( .A1(n1023), .A2(G868), .ZN(n768) );
  NAND2_X1 U849 ( .A1(n769), .A2(n768), .ZN(G284) );
  INV_X1 U850 ( .A(G868), .ZN(n809) );
  NOR2_X1 U851 ( .A1(G286), .A2(n809), .ZN(n771) );
  NOR2_X1 U852 ( .A1(G868), .A2(G299), .ZN(n770) );
  NOR2_X1 U853 ( .A1(n771), .A2(n770), .ZN(G297) );
  NAND2_X1 U854 ( .A1(n772), .A2(G559), .ZN(n773) );
  NAND2_X1 U855 ( .A1(n773), .A2(n1023), .ZN(n774) );
  XNOR2_X1 U856 ( .A(n774), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U857 ( .A1(G559), .A2(n809), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n1023), .A2(n775), .ZN(n776) );
  XNOR2_X1 U859 ( .A(n776), .B(KEYINPUT75), .ZN(n778) );
  NOR2_X1 U860 ( .A1(n945), .A2(G868), .ZN(n777) );
  NOR2_X1 U861 ( .A1(n778), .A2(n777), .ZN(G282) );
  NAND2_X1 U862 ( .A1(n1001), .A2(G123), .ZN(n779) );
  XNOR2_X1 U863 ( .A(n779), .B(KEYINPUT18), .ZN(n781) );
  NAND2_X1 U864 ( .A1(G111), .A2(n1002), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U866 ( .A1(G99), .A2(n1005), .ZN(n783) );
  NAND2_X1 U867 ( .A1(G135), .A2(n521), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U869 ( .A1(n785), .A2(n784), .ZN(n996) );
  XNOR2_X1 U870 ( .A(n996), .B(G2096), .ZN(n787) );
  INV_X1 U871 ( .A(G2100), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(G156) );
  NAND2_X1 U873 ( .A1(n1023), .A2(G559), .ZN(n807) );
  XNOR2_X1 U874 ( .A(n945), .B(n807), .ZN(n788) );
  NOR2_X1 U875 ( .A1(n788), .A2(G860), .ZN(n800) );
  NAND2_X1 U876 ( .A1(G80), .A2(n789), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G93), .A2(n790), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n799) );
  NAND2_X1 U879 ( .A1(G55), .A2(n793), .ZN(n794) );
  XNOR2_X1 U880 ( .A(n794), .B(KEYINPUT76), .ZN(n797) );
  NAND2_X1 U881 ( .A1(n795), .A2(G67), .ZN(n796) );
  NAND2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n810) );
  XOR2_X1 U884 ( .A(n800), .B(n810), .Z(G145) );
  XNOR2_X1 U885 ( .A(KEYINPUT19), .B(G303), .ZN(n801) );
  XNOR2_X1 U886 ( .A(n801), .B(n945), .ZN(n804) );
  XNOR2_X1 U887 ( .A(n954), .B(G290), .ZN(n802) );
  XNOR2_X1 U888 ( .A(n802), .B(G305), .ZN(n803) );
  XNOR2_X1 U889 ( .A(n804), .B(n803), .ZN(n806) );
  XOR2_X1 U890 ( .A(G288), .B(n810), .Z(n805) );
  XNOR2_X1 U891 ( .A(n806), .B(n805), .ZN(n1022) );
  XOR2_X1 U892 ( .A(n1022), .B(n807), .Z(n808) );
  NAND2_X1 U893 ( .A1(G868), .A2(n808), .ZN(n812) );
  NAND2_X1 U894 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U895 ( .A1(n812), .A2(n811), .ZN(G295) );
  NAND2_X1 U896 ( .A1(G2078), .A2(G2084), .ZN(n813) );
  XOR2_X1 U897 ( .A(KEYINPUT20), .B(n813), .Z(n814) );
  NAND2_X1 U898 ( .A1(n814), .A2(G2090), .ZN(n815) );
  XNOR2_X1 U899 ( .A(n815), .B(KEYINPUT78), .ZN(n816) );
  XNOR2_X1 U900 ( .A(KEYINPUT21), .B(n816), .ZN(n817) );
  NAND2_X1 U901 ( .A1(G2072), .A2(n817), .ZN(G158) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U903 ( .A(KEYINPUT68), .B(G132), .Z(G219) );
  NOR2_X1 U904 ( .A1(G236), .A2(G237), .ZN(n818) );
  NAND2_X1 U905 ( .A1(G69), .A2(n818), .ZN(n819) );
  XNOR2_X1 U906 ( .A(KEYINPUT79), .B(n819), .ZN(n820) );
  NAND2_X1 U907 ( .A1(n820), .A2(G108), .ZN(n968) );
  NAND2_X1 U908 ( .A1(n968), .A2(G567), .ZN(n825) );
  NOR2_X1 U909 ( .A1(G219), .A2(G220), .ZN(n821) );
  XOR2_X1 U910 ( .A(KEYINPUT22), .B(n821), .Z(n822) );
  NOR2_X1 U911 ( .A1(G218), .A2(n822), .ZN(n823) );
  NAND2_X1 U912 ( .A1(G96), .A2(n823), .ZN(n969) );
  NAND2_X1 U913 ( .A1(n969), .A2(G2106), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n825), .A2(n824), .ZN(n970) );
  NAND2_X1 U915 ( .A1(G483), .A2(G661), .ZN(n826) );
  NOR2_X1 U916 ( .A1(n970), .A2(n826), .ZN(n842) );
  NAND2_X1 U917 ( .A1(n842), .A2(G36), .ZN(n827) );
  XNOR2_X1 U918 ( .A(KEYINPUT80), .B(n827), .ZN(G176) );
  XNOR2_X1 U919 ( .A(G1341), .B(G2454), .ZN(n828) );
  XNOR2_X1 U920 ( .A(n828), .B(G2430), .ZN(n829) );
  XNOR2_X1 U921 ( .A(n829), .B(G1348), .ZN(n835) );
  XOR2_X1 U922 ( .A(G2443), .B(G2427), .Z(n831) );
  XNOR2_X1 U923 ( .A(G2438), .B(G2446), .ZN(n830) );
  XNOR2_X1 U924 ( .A(n831), .B(n830), .ZN(n833) );
  XOR2_X1 U925 ( .A(G2451), .B(G2435), .Z(n832) );
  XNOR2_X1 U926 ( .A(n833), .B(n832), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n835), .B(n834), .ZN(n836) );
  NAND2_X1 U928 ( .A1(n836), .A2(G14), .ZN(n1028) );
  XNOR2_X1 U929 ( .A(KEYINPUT101), .B(n1028), .ZN(G401) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n837), .ZN(G217) );
  INV_X1 U931 ( .A(G661), .ZN(n839) );
  NAND2_X1 U932 ( .A1(G2), .A2(G15), .ZN(n838) );
  NOR2_X1 U933 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U934 ( .A(KEYINPUT102), .B(n840), .Z(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(G188) );
  NAND2_X1 U938 ( .A1(G100), .A2(n1005), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n843), .B(KEYINPUT106), .ZN(n850) );
  NAND2_X1 U940 ( .A1(G136), .A2(n521), .ZN(n845) );
  NAND2_X1 U941 ( .A1(G112), .A2(n1002), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n845), .A2(n844), .ZN(n848) );
  NAND2_X1 U943 ( .A1(n1001), .A2(G124), .ZN(n846) );
  XOR2_X1 U944 ( .A(KEYINPUT44), .B(n846), .Z(n847) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U947 ( .A(KEYINPUT107), .B(n851), .ZN(G162) );
  XOR2_X1 U948 ( .A(G1976), .B(G23), .Z(n853) );
  XOR2_X1 U949 ( .A(G1971), .B(G22), .Z(n852) );
  NAND2_X1 U950 ( .A1(n853), .A2(n852), .ZN(n855) );
  XNOR2_X1 U951 ( .A(G24), .B(G1986), .ZN(n854) );
  NOR2_X1 U952 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U953 ( .A(KEYINPUT58), .B(n856), .Z(n875) );
  XNOR2_X1 U954 ( .A(G1961), .B(G5), .ZN(n872) );
  XOR2_X1 U955 ( .A(KEYINPUT124), .B(G4), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1348), .B(KEYINPUT59), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n866) );
  XOR2_X1 U958 ( .A(G1341), .B(G19), .Z(n861) );
  XNOR2_X1 U959 ( .A(n859), .B(G20), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n863) );
  XNOR2_X1 U961 ( .A(G6), .B(G1981), .ZN(n862) );
  NOR2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n864), .B(KEYINPUT123), .ZN(n865) );
  NOR2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U965 ( .A(KEYINPUT60), .B(n867), .Z(n869) );
  XNOR2_X1 U966 ( .A(G1966), .B(G21), .ZN(n868) );
  NOR2_X1 U967 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U968 ( .A(KEYINPUT125), .B(n870), .ZN(n871) );
  NOR2_X1 U969 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U970 ( .A(KEYINPUT126), .B(n873), .Z(n874) );
  NOR2_X1 U971 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U972 ( .A(KEYINPUT61), .B(n876), .Z(n878) );
  XNOR2_X1 U973 ( .A(G16), .B(KEYINPUT122), .ZN(n877) );
  NOR2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n904) );
  XOR2_X1 U975 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n935) );
  XNOR2_X1 U976 ( .A(G25), .B(n879), .ZN(n880) );
  NAND2_X1 U977 ( .A1(n880), .A2(G28), .ZN(n891) );
  XOR2_X1 U978 ( .A(G2072), .B(G33), .Z(n881) );
  XNOR2_X1 U979 ( .A(KEYINPUT117), .B(n881), .ZN(n883) );
  XNOR2_X1 U980 ( .A(G26), .B(G2067), .ZN(n882) );
  NOR2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(KEYINPUT118), .B(n884), .ZN(n889) );
  XNOR2_X1 U983 ( .A(n885), .B(G27), .ZN(n887) );
  XNOR2_X1 U984 ( .A(G32), .B(G1996), .ZN(n886) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n888) );
  NAND2_X1 U986 ( .A1(n889), .A2(n888), .ZN(n890) );
  NOR2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n893) );
  XNOR2_X1 U988 ( .A(KEYINPUT53), .B(KEYINPUT119), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n898) );
  XNOR2_X1 U990 ( .A(G2084), .B(KEYINPUT54), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n894), .B(G34), .ZN(n896) );
  XNOR2_X1 U992 ( .A(G35), .B(G2090), .ZN(n895) );
  NOR2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  NAND2_X1 U994 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n935), .B(n899), .ZN(n901) );
  INV_X1 U996 ( .A(G29), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U998 ( .A1(G11), .A2(n902), .ZN(n903) );
  NOR2_X1 U999 ( .A1(n904), .A2(n903), .ZN(n939) );
  NOR2_X1 U1000 ( .A1(n905), .A2(n996), .ZN(n914) );
  XNOR2_X1 U1001 ( .A(G160), .B(G2084), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n912) );
  XOR2_X1 U1003 ( .A(G2090), .B(G162), .Z(n908) );
  NOR2_X1 U1004 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n910), .B(KEYINPUT51), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1007 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1009 ( .A(n917), .B(KEYINPUT114), .ZN(n919) );
  NAND2_X1 U1010 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1011 ( .A(KEYINPUT115), .B(n920), .Z(n933) );
  NAND2_X1 U1012 ( .A1(G103), .A2(n1005), .ZN(n922) );
  NAND2_X1 U1013 ( .A1(G139), .A2(n521), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1015 ( .A(KEYINPUT108), .B(n923), .ZN(n928) );
  NAND2_X1 U1016 ( .A1(G127), .A2(n1001), .ZN(n925) );
  NAND2_X1 U1017 ( .A1(G115), .A2(n1002), .ZN(n924) );
  NAND2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1019 ( .A(KEYINPUT47), .B(n926), .Z(n927) );
  NOR2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(n1018) );
  XOR2_X1 U1021 ( .A(G2072), .B(n1018), .Z(n930) );
  XOR2_X1 U1022 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1024 ( .A(KEYINPUT50), .B(n931), .Z(n932) );
  NOR2_X1 U1025 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1026 ( .A(KEYINPUT52), .B(n934), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1028 ( .A1(n937), .A2(G29), .ZN(n938) );
  NAND2_X1 U1029 ( .A1(n939), .A2(n938), .ZN(n966) );
  XOR2_X1 U1030 ( .A(KEYINPUT56), .B(G16), .Z(n964) );
  XNOR2_X1 U1031 ( .A(G171), .B(G1961), .ZN(n941) );
  NAND2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1033 ( .A1(n943), .A2(n942), .ZN(n953) );
  XNOR2_X1 U1034 ( .A(G1971), .B(G166), .ZN(n944) );
  XNOR2_X1 U1035 ( .A(n944), .B(KEYINPUT120), .ZN(n949) );
  XOR2_X1 U1036 ( .A(G1348), .B(n1023), .Z(n947) );
  XNOR2_X1 U1037 ( .A(n945), .B(G1341), .ZN(n946) );
  NOR2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1039 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1040 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1041 ( .A1(n953), .A2(n952), .ZN(n961) );
  XNOR2_X1 U1042 ( .A(n954), .B(G1956), .ZN(n959) );
  XOR2_X1 U1043 ( .A(G168), .B(G1966), .Z(n955) );
  NOR2_X1 U1044 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1045 ( .A(KEYINPUT57), .B(n957), .Z(n958) );
  NAND2_X1 U1046 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1047 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1048 ( .A(KEYINPUT121), .B(n962), .Z(n963) );
  NOR2_X1 U1049 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1050 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1051 ( .A(n967), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1052 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1053 ( .A(G108), .ZN(G238) );
  INV_X1 U1054 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1055 ( .A1(n969), .A2(n968), .ZN(G325) );
  INV_X1 U1056 ( .A(G325), .ZN(G261) );
  INV_X1 U1057 ( .A(n970), .ZN(G319) );
  XOR2_X1 U1058 ( .A(KEYINPUT103), .B(G2084), .Z(n972) );
  XNOR2_X1 U1059 ( .A(G2078), .B(G2067), .ZN(n971) );
  XNOR2_X1 U1060 ( .A(n972), .B(n971), .ZN(n973) );
  XOR2_X1 U1061 ( .A(n973), .B(G2678), .Z(n975) );
  XNOR2_X1 U1062 ( .A(G2072), .B(KEYINPUT42), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(n975), .B(n974), .ZN(n979) );
  XOR2_X1 U1064 ( .A(G2100), .B(G2096), .Z(n977) );
  XNOR2_X1 U1065 ( .A(G2090), .B(KEYINPUT43), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n977), .B(n976), .ZN(n978) );
  XOR2_X1 U1067 ( .A(n979), .B(n978), .Z(G227) );
  XOR2_X1 U1068 ( .A(G2474), .B(G1991), .Z(n981) );
  XNOR2_X1 U1069 ( .A(G1961), .B(G1976), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n981), .B(n980), .ZN(n982) );
  XOR2_X1 U1071 ( .A(n982), .B(G1956), .Z(n984) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G1996), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(n984), .B(n983), .ZN(n988) );
  XOR2_X1 U1074 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n986) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G1981), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(n986), .B(n985), .ZN(n987) );
  XOR2_X1 U1077 ( .A(n988), .B(n987), .Z(n990) );
  XNOR2_X1 U1078 ( .A(G1986), .B(KEYINPUT41), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(n990), .B(n989), .ZN(G229) );
  XOR2_X1 U1080 ( .A(G164), .B(G162), .Z(n991) );
  XNOR2_X1 U1081 ( .A(n992), .B(n991), .ZN(n1000) );
  XOR2_X1 U1082 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n994) );
  XNOR2_X1 U1083 ( .A(KEYINPUT110), .B(KEYINPUT48), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n994), .B(n993), .ZN(n995) );
  XOR2_X1 U1085 ( .A(n995), .B(KEYINPUT112), .Z(n998) );
  XNOR2_X1 U1086 ( .A(n996), .B(KEYINPUT111), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n998), .B(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(n1000), .B(n999), .Z(n1016) );
  NAND2_X1 U1089 ( .A1(G130), .A2(n1001), .ZN(n1004) );
  NAND2_X1 U1090 ( .A1(G118), .A2(n1002), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  NAND2_X1 U1092 ( .A1(G106), .A2(n1005), .ZN(n1008) );
  NAND2_X1 U1093 ( .A1(G142), .A2(n521), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(n1009), .B(KEYINPUT45), .Z(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(n1013), .B(n1012), .Z(n1014) );
  XNOR2_X1 U1098 ( .A(G160), .B(n1014), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(n1016), .B(n1015), .ZN(n1020) );
  XOR2_X1 U1100 ( .A(n1018), .B(n1017), .Z(n1019) );
  XNOR2_X1 U1101 ( .A(n1020), .B(n1019), .ZN(n1021) );
  NOR2_X1 U1102 ( .A1(G37), .A2(n1021), .ZN(G395) );
  XOR2_X1 U1103 ( .A(KEYINPUT113), .B(n1022), .Z(n1025) );
  XNOR2_X1 U1104 ( .A(n1023), .B(G286), .ZN(n1024) );
  XNOR2_X1 U1105 ( .A(n1025), .B(n1024), .ZN(n1026) );
  XNOR2_X1 U1106 ( .A(n1026), .B(G171), .ZN(n1027) );
  NOR2_X1 U1107 ( .A1(G37), .A2(n1027), .ZN(G397) );
  NAND2_X1 U1108 ( .A1(G319), .A2(n1028), .ZN(n1031) );
  NOR2_X1 U1109 ( .A1(G227), .A2(G229), .ZN(n1029) );
  XNOR2_X1 U1110 ( .A(KEYINPUT49), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1111 ( .A1(n1031), .A2(n1030), .ZN(n1033) );
  NOR2_X1 U1112 ( .A1(G395), .A2(G397), .ZN(n1032) );
  NAND2_X1 U1113 ( .A1(n1033), .A2(n1032), .ZN(G225) );
  INV_X1 U1114 ( .A(G225), .ZN(G308) );
  INV_X1 U1115 ( .A(G69), .ZN(G235) );
endmodule

