//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT65), .B(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G77), .A2(G244), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(G232), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G68), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G50), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  XNOR2_X1  g0044(.A(KEYINPUT8), .B(G58), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n206), .A2(G20), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  AND2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  OAI22_X1  g0055(.A1(new_n248), .A2(new_n255), .B1(new_n254), .B2(new_n246), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n201), .B1(new_n217), .B2(G58), .ZN(new_n257));
  INV_X1    g0057(.A(G159), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n257), .A2(new_n207), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G68), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT76), .B1(new_n263), .B2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT76), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(new_n266), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n207), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n262), .B1(new_n270), .B2(KEYINPUT7), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT7), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n272), .A3(new_n207), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n261), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n251), .B1(new_n274), .B2(KEYINPUT16), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT16), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n266), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(KEYINPUT77), .A3(new_n272), .A4(new_n207), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(G20), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n279), .A2(new_n282), .A3(new_n217), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n276), .B1(new_n283), .B2(new_n261), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n256), .B1(new_n275), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G1), .A3(G13), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n290), .A2(new_n286), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n288), .B1(new_n291), .B2(G232), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G226), .A2(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G223), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(G1698), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n295), .A2(new_n264), .A3(new_n267), .A4(new_n268), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT78), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G87), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT67), .B1(new_n300), .B2(new_n250), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT67), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n213), .A2(new_n302), .A3(new_n289), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n292), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n292), .C1(new_n305), .C2(new_n306), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT17), .B1(new_n285), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n256), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(G68), .A3(new_n273), .ZN(new_n316));
  INV_X1    g0116(.A(new_n261), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT16), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n249), .A2(new_n250), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n319), .A3(new_n284), .ZN(new_n320));
  AND4_X1   g0120(.A1(KEYINPUT17), .A2(new_n312), .A3(new_n314), .A4(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT80), .B1(new_n313), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT17), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n314), .ZN(new_n324));
  INV_X1    g0124(.A(new_n311), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n296), .A2(new_n298), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT78), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(new_n304), .A3(new_n299), .ZN(new_n328));
  AOI21_X1  g0128(.A(G200), .B1(new_n328), .B2(new_n292), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n323), .B1(new_n324), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT80), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n312), .A2(KEYINPUT17), .A3(new_n320), .A4(new_n314), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n307), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT79), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(new_n292), .C1(new_n305), .C2(new_n306), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n337), .B1(new_n336), .B2(new_n339), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n324), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n339), .ZN(new_n346));
  AOI21_X1  g0146(.A(G169), .B1(new_n328), .B2(new_n292), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT79), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n340), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(KEYINPUT18), .A3(new_n324), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n322), .A2(new_n334), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n247), .A2(G50), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n255), .A2(new_n352), .B1(G50), .B2(new_n254), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n207), .A2(G33), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n355), .B1(new_n356), .B2(new_n245), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n319), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT9), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n353), .B1(new_n319), .B2(new_n357), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT9), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n291), .A2(G226), .ZN(new_n364));
  INV_X1    g0164(.A(new_n288), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G1698), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n281), .A2(G222), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G77), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n281), .A2(G1698), .ZN(new_n370));
  OAI221_X1 g0170(.A(new_n368), .B1(new_n369), .B2(new_n281), .C1(new_n370), .C2(new_n294), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n371), .B2(new_n304), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n361), .B(new_n363), .C1(new_n308), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(G190), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT10), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n361), .A2(new_n363), .ZN(new_n377));
  INV_X1    g0177(.A(new_n372), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G200), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n377), .A2(new_n379), .A3(new_n380), .A4(new_n374), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT69), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n247), .A2(G77), .ZN(new_n384));
  OR3_X1    g0184(.A1(new_n255), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n383), .B1(new_n255), .B2(new_n384), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n252), .A2(new_n207), .A3(G1), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n369), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G20), .A2(G77), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n390), .B1(new_n245), .B2(new_n260), .C1(new_n356), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n319), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n387), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n288), .B1(new_n291), .B2(G244), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT68), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n281), .A2(G232), .A3(new_n367), .ZN(new_n397));
  INV_X1    g0197(.A(G107), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n397), .B1(new_n398), .B2(new_n281), .C1(new_n370), .C2(new_n219), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n304), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n308), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n291), .A2(G244), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n365), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n404), .A2(KEYINPUT68), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(KEYINPUT68), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n400), .B(new_n310), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n394), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n394), .ZN(new_n409));
  OAI21_X1  g0209(.A(G169), .B1(new_n396), .B2(new_n401), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n400), .B(G179), .C1(new_n405), .C2(new_n406), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n378), .A2(new_n338), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n372), .A2(new_n335), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n359), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n382), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n268), .A2(new_n277), .A3(G226), .A4(new_n367), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n268), .A2(new_n277), .A3(G232), .A4(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n304), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n288), .B1(new_n291), .B2(G238), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n424), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n426), .B1(KEYINPUT13), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G190), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n217), .A2(new_n207), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n260), .A2(new_n202), .B1(new_n356), .B2(new_n369), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n319), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT11), .ZN(new_n433));
  OR3_X1    g0233(.A1(new_n254), .A2(KEYINPUT12), .A3(G68), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n254), .B2(new_n217), .ZN(new_n436));
  INV_X1    g0236(.A(new_n255), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n262), .B1(new_n206), .B2(G20), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n434), .A2(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n425), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n427), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G200), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n429), .A2(new_n441), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n428), .A2(G179), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n425), .B1(new_n423), .B2(new_n424), .ZN(new_n450));
  OAI21_X1  g0250(.A(G169), .B1(new_n426), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g0251(.A(KEYINPUT74), .B(KEYINPUT14), .Z(new_n452));
  OAI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(KEYINPUT72), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT72), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(G169), .C1(new_n426), .C2(new_n450), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT73), .B1(new_n458), .B2(KEYINPUT14), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT73), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT14), .ZN(new_n461));
  AOI211_X1 g0261(.A(new_n460), .B(new_n461), .C1(new_n455), .C2(new_n457), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n454), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n448), .B1(new_n463), .B2(new_n440), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n351), .B(new_n418), .C1(new_n464), .C2(KEYINPUT75), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n440), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n447), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT75), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT81), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n322), .A2(new_n334), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n345), .A2(new_n350), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n418), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n467), .B2(new_n468), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT81), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n464), .A2(KEYINPUT75), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n206), .A2(G33), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n251), .A2(new_n254), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT85), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n481), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT85), .A2(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n480), .A2(new_n481), .B1(new_n254), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n207), .B1(new_n483), .B2(new_n484), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n263), .A2(G97), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G283), .ZN(new_n489));
  AOI21_X1  g0289(.A(G20), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n319), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(KEYINPUT20), .B(new_n319), .C1(new_n487), .C2(new_n490), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n486), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n301), .A2(new_n303), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n278), .A2(G303), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G264), .A2(G1698), .ZN(new_n498));
  INV_X1    g0298(.A(G257), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(new_n264), .A3(new_n267), .A4(new_n268), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n496), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G45), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(G1), .ZN(new_n504));
  NAND2_X1  g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(G270), .A3(new_n290), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT5), .B(G41), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G274), .A3(new_n504), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(G169), .B1(new_n502), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n495), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n509), .A2(new_n511), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n501), .A2(new_n497), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n304), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n338), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n493), .A2(new_n494), .ZN(new_n520));
  INV_X1    g0320(.A(new_n486), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n514), .A2(KEYINPUT21), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n518), .A2(G190), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n502), .A2(new_n512), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(G200), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n495), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n335), .B1(new_n515), .B2(new_n517), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT21), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT87), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(KEYINPUT87), .B(new_n530), .C1(new_n495), .C2(new_n513), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n523), .B(new_n527), .C1(new_n531), .C2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT88), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT87), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n514), .B2(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n532), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n539), .A2(KEYINPUT88), .A3(new_n523), .A4(new_n527), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT83), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT6), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G97), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n544), .A2(new_n546), .A3(G107), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n279), .A2(new_n282), .A3(G107), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n251), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n388), .A2(G97), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n480), .B2(G97), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n542), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT4), .ZN(new_n556));
  INV_X1    g0356(.A(G244), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(G1698), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n556), .B1(new_n269), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n367), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n281), .A2(G250), .A3(G1698), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n489), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n304), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n508), .A2(new_n290), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n511), .B1(new_n566), .B2(new_n499), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n335), .ZN(new_n570));
  INV_X1    g0370(.A(new_n551), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n547), .B1(new_n544), .B2(new_n543), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n572), .A2(new_n207), .B1(new_n369), .B2(new_n260), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n319), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n554), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(KEYINPUT83), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n567), .A2(KEYINPUT82), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n578), .B(new_n511), .C1(new_n566), .C2(new_n499), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n338), .A3(new_n565), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n555), .A2(new_n570), .A3(new_n576), .A4(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n552), .A2(new_n554), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n560), .A2(new_n489), .A3(new_n563), .A4(new_n562), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n567), .B1(new_n584), .B2(new_n304), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G190), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n577), .A2(new_n579), .B1(new_n584), .B2(new_n304), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n583), .B(new_n586), .C1(new_n308), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT84), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT84), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n582), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n391), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(new_n254), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT19), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n421), .B2(G20), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n264), .A2(new_n267), .A3(new_n207), .A4(new_n268), .ZN(new_n598));
  XNOR2_X1  g0398(.A(KEYINPUT86), .B(G87), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n599), .A2(G97), .A3(G107), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n421), .A2(new_n596), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(G20), .ZN(new_n602));
  OAI221_X1 g0402(.A(new_n597), .B1(new_n598), .B2(new_n262), .C1(new_n600), .C2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n595), .B1(new_n603), .B2(new_n319), .ZN(new_n604));
  INV_X1    g0404(.A(new_n480), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n594), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n263), .B1(new_n483), .B2(new_n484), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  MUX2_X1   g0409(.A(new_n219), .B(new_n557), .S(G1698), .Z(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n269), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n304), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n300), .A2(new_n250), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n504), .A2(G274), .ZN(new_n614));
  OAI21_X1  g0414(.A(G250), .B1(new_n503), .B2(G1), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n335), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n611), .B2(new_n304), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n338), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n618), .A2(G200), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(G190), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n605), .A2(G87), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n604), .A2(new_n626), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n607), .A2(new_n622), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n253), .A2(G20), .A3(new_n398), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT25), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(G107), .B2(new_n605), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n264), .A2(new_n267), .A3(new_n268), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n633));
  INV_X1    g0433(.A(G87), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G20), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT22), .B1(new_n281), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT23), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n207), .B2(G107), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n398), .A2(KEYINPUT23), .A3(G20), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n608), .A2(new_n207), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n633), .A2(KEYINPUT24), .A3(new_n637), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n319), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n485), .A2(new_n207), .A3(G33), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n640), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n636), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT24), .B1(new_n647), .B2(new_n633), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n631), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(G257), .A2(G1698), .ZN(new_n650));
  INV_X1    g0450(.A(G250), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(G1698), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n652), .A2(new_n264), .A3(new_n267), .A4(new_n268), .ZN(new_n653));
  NAND2_X1  g0453(.A1(G33), .A2(G294), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n304), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n613), .B1(new_n504), .B2(new_n510), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G264), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n310), .A2(new_n656), .A3(new_n511), .A4(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n655), .A2(new_n304), .B1(new_n657), .B2(G264), .ZN(new_n660));
  AOI21_X1  g0460(.A(G200), .B1(new_n660), .B2(new_n511), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n649), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT24), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n637), .A2(new_n641), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT22), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n598), .A2(new_n666), .A3(new_n634), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n664), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n319), .A3(new_n642), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n660), .A2(new_n511), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G169), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n660), .A2(G179), .A3(new_n511), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n669), .A2(new_n631), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT89), .B1(new_n663), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n649), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n669), .B(new_n631), .C1(new_n659), .C2(new_n661), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n628), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n478), .A2(new_n541), .A3(new_n593), .A4(new_n680), .ZN(G372));
  INV_X1    g0481(.A(new_n589), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n539), .A2(new_n523), .A3(new_n676), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n628), .A2(new_n663), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT26), .B1(new_n628), .B2(new_n582), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n574), .A2(new_n575), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n570), .A2(new_n581), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n625), .A2(new_n627), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT26), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n604), .A2(new_n606), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(new_n621), .A3(new_n619), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n689), .A2(new_n690), .A3(new_n691), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n686), .A2(new_n694), .A3(new_n693), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n685), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n478), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n346), .A2(new_n347), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n324), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n700), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n324), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n410), .A2(new_n411), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n394), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n466), .B1(new_n448), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n705), .B1(new_n708), .B2(new_n471), .ZN(new_n709));
  INV_X1    g0509(.A(new_n382), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n417), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n697), .A2(new_n712), .ZN(G369));
  NAND2_X1  g0513(.A1(new_n253), .A2(new_n207), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n714), .A2(KEYINPUT27), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(KEYINPUT27), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G213), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G343), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n495), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n541), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n539), .A2(new_n523), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n720), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G330), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n719), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n674), .A2(new_n679), .B1(new_n649), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n676), .A2(new_n719), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n719), .B(KEYINPUT91), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n673), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n722), .A2(new_n727), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n728), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n731), .A2(new_n734), .A3(new_n736), .ZN(G399));
  INV_X1    g0537(.A(new_n210), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G41), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n600), .A2(new_n481), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(G1), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n216), .B2(new_n740), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT29), .B1(new_n696), .B2(new_n733), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT26), .B1(new_n628), .B2(new_n688), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n693), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n628), .A2(new_n582), .A3(KEYINPUT26), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n589), .A2(KEYINPUT93), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT93), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n582), .A2(new_n588), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n751), .A2(new_n683), .A3(new_n684), .A4(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n727), .B1(new_n750), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n746), .B1(KEYINPUT29), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n541), .A2(new_n680), .A3(new_n593), .A4(new_n733), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n525), .A2(new_n620), .A3(G179), .A4(new_n660), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n569), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n580), .A2(new_n565), .B1(new_n511), .B2(new_n660), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n525), .A2(new_n620), .A3(G179), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n759), .A2(KEYINPUT30), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT30), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n758), .B2(new_n569), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(KEYINPUT31), .A3(new_n732), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT92), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n762), .B2(new_n764), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n760), .A2(new_n761), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n620), .A2(new_n660), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n770), .A2(new_n519), .A3(KEYINPUT30), .A4(new_n585), .ZN(new_n771));
  AND4_X1   g0571(.A1(new_n767), .A2(new_n769), .A3(new_n764), .A4(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n727), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT31), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n757), .A2(new_n766), .A3(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(G330), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n756), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n745), .B1(new_n778), .B2(G1), .ZN(G364));
  NOR2_X1   g0579(.A1(new_n252), .A2(G20), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G45), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n740), .A2(G1), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n724), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G330), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n784), .B2(new_n726), .ZN(new_n785));
  INV_X1    g0585(.A(new_n782), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT95), .Z(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n210), .A2(new_n281), .ZN(new_n792));
  XNOR2_X1  g0592(.A(G355), .B(KEYINPUT94), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n792), .A2(new_n793), .B1(G116), .B2(new_n210), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n216), .A2(new_n503), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n240), .B2(new_n503), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n738), .A2(new_n632), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n250), .B1(G20), .B2(new_n335), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n790), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT97), .Z(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT98), .Z(new_n803));
  NAND2_X1  g0603(.A1(new_n338), .A2(new_n308), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT100), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G190), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G294), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n207), .A2(new_n310), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n308), .A2(G179), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n207), .A2(G190), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n810), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n811), .A2(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n338), .A2(G200), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n816), .B1(G311), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n338), .A2(new_n308), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n809), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n281), .B1(new_n823), .B2(G326), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n813), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT33), .B(G317), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n809), .A2(new_n817), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n826), .A2(new_n827), .B1(new_n829), .B2(G322), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n808), .A2(new_n820), .A3(new_n824), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n805), .A2(new_n813), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(KEYINPUT101), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(KEYINPUT101), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n831), .B1(G329), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n811), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n599), .A2(new_n838), .B1(new_n819), .B2(G77), .ZN(new_n839));
  INV_X1    g0639(.A(new_n814), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n278), .B1(new_n840), .B2(G107), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(new_n202), .C2(new_n822), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n807), .A2(G97), .B1(G68), .B2(new_n826), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT102), .Z(new_n844));
  XOR2_X1   g0644(.A(new_n828), .B(KEYINPUT99), .Z(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n842), .B(new_n844), .C1(G58), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n835), .A2(new_n258), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT32), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n837), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n798), .A2(new_n803), .B1(new_n850), .B2(new_n800), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n786), .B1(new_n791), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n785), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G396));
  NOR2_X1   g0654(.A1(new_n799), .A2(new_n787), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n782), .B1(new_n369), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n823), .A2(G137), .B1(new_n819), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G150), .ZN(new_n858));
  INV_X1    g0658(.A(G143), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n857), .B1(new_n858), .B2(new_n825), .C1(new_n845), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n861), .A2(KEYINPUT34), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n632), .B1(new_n202), .B2(new_n811), .C1(new_n262), .C2(new_n814), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n807), .B2(G58), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(KEYINPUT34), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n836), .A2(G132), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n862), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G303), .A2(new_n823), .B1(new_n838), .B2(G107), .ZN(new_n868));
  INV_X1    g0668(.A(new_n485), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n818), .ZN(new_n870));
  INV_X1    g0670(.A(G294), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n278), .B1(new_n828), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(KEYINPUT103), .B(G283), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n825), .A2(new_n873), .B1(new_n814), .B2(new_n634), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n807), .ZN(new_n876));
  INV_X1    g0676(.A(G311), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n875), .B1(new_n546), .B2(new_n876), .C1(new_n877), .C2(new_n835), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n867), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n707), .A2(new_n727), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n409), .A2(new_n719), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n408), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n880), .B1(new_n882), .B2(new_n707), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n856), .B1(new_n879), .B2(new_n800), .C1(new_n883), .C2(new_n788), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n696), .A2(new_n733), .ZN(new_n885));
  INV_X1    g0685(.A(new_n883), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n733), .B(new_n883), .C1(new_n685), .C2(new_n695), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n776), .A2(G330), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n782), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n884), .B1(new_n892), .B2(new_n893), .ZN(G384));
  NOR2_X1   g0694(.A1(new_n780), .A2(new_n206), .ZN(new_n895));
  OAI211_X1 g0695(.A(KEYINPUT31), .B(new_n727), .C1(new_n768), .C2(new_n772), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n757), .A2(new_n775), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n478), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT104), .Z(new_n899));
  NOR2_X1   g0699(.A1(new_n441), .A2(new_n719), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n456), .B1(new_n445), .B2(G169), .ZN(new_n902));
  INV_X1    g0702(.A(new_n457), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT14), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n460), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n458), .A2(KEYINPUT73), .A3(KEYINPUT14), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n453), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n447), .B(new_n901), .C1(new_n907), .C2(new_n441), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n463), .A2(new_n900), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n910), .A2(new_n897), .A3(new_n883), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n285), .A2(new_n312), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n318), .A2(new_n319), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n274), .A2(KEYINPUT16), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n314), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n698), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n718), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n912), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT37), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n324), .A2(new_n718), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n343), .A2(new_n920), .A3(new_n912), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(KEYINPUT38), .B(new_n923), .C1(new_n351), .C2(new_n917), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n313), .A2(new_n321), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n921), .B1(new_n704), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n912), .A2(new_n920), .A3(new_n921), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n912), .A2(new_n699), .A3(new_n921), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n928), .A2(new_n343), .B1(new_n929), .B2(KEYINPUT37), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n925), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n911), .A2(KEYINPUT40), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n917), .B1(new_n471), .B2(new_n472), .ZN(new_n934));
  INV_X1    g0734(.A(new_n923), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n925), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n924), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n911), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n933), .B1(new_n938), .B2(KEYINPUT40), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n899), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n899), .A2(new_n939), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(G330), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n466), .A2(new_n727), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n924), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n332), .B1(new_n331), .B2(new_n333), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT18), .B1(new_n349), .B2(new_n324), .ZN(new_n948));
  AOI221_X4 g0748(.A(new_n344), .B1(new_n314), .B2(new_n320), .C1(new_n348), .C2(new_n340), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n946), .A2(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n917), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT38), .B1(new_n952), .B2(new_n923), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT39), .B1(new_n945), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT39), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n924), .A2(new_n931), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n944), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n880), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n888), .A2(new_n958), .B1(new_n908), .B2(new_n909), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n937), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n705), .A2(new_n717), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n957), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n711), .B1(new_n478), .B2(new_n756), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n895), .B1(new_n942), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n942), .B2(new_n965), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n369), .B(new_n216), .C1(new_n217), .C2(G58), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n262), .A2(G50), .ZN(new_n969));
  OAI211_X1 g0769(.A(G1), .B(new_n252), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n215), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n971), .B(G116), .C1(KEYINPUT35), .C2(new_n549), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(KEYINPUT35), .B2(new_n549), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT36), .Z(new_n974));
  NAND3_X1  g0774(.A1(new_n967), .A2(new_n970), .A3(new_n974), .ZN(G367));
  AOI22_X1  g0775(.A1(new_n797), .A2(new_n235), .B1(new_n738), .B2(new_n594), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n802), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n786), .B1(new_n977), .B2(KEYINPUT107), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(KEYINPUT107), .B2(new_n977), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n719), .B1(new_n604), .B2(new_n626), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n690), .B2(new_n693), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n693), .A2(new_n980), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G150), .A2(new_n829), .B1(new_n840), .B2(G77), .ZN(new_n984));
  INV_X1    g0784(.A(G58), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n984), .B1(new_n985), .B2(new_n811), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n281), .B1(new_n818), .B2(new_n202), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n822), .A2(new_n859), .B1(new_n825), .B2(new_n258), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n807), .A2(G68), .ZN(new_n990));
  INV_X1    g0790(.A(G137), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n989), .B(new_n990), .C1(new_n991), .C2(new_n835), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT108), .Z(new_n993));
  NAND3_X1  g0793(.A1(new_n838), .A2(KEYINPUT46), .A3(G116), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n546), .B2(new_n814), .C1(new_n871), .C2(new_n825), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT46), .B1(new_n838), .B2(new_n485), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n822), .A2(new_n877), .B1(new_n818), .B2(new_n873), .ZN(new_n997));
  OR3_X1    g0797(.A1(new_n996), .A2(new_n997), .A3(new_n632), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n995), .B(new_n998), .C1(G303), .C2(new_n846), .ZN(new_n999));
  INV_X1    g0799(.A(G317), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n999), .B1(new_n398), .B2(new_n876), .C1(new_n1000), .C2(new_n835), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT47), .B1(new_n993), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n993), .A2(KEYINPUT47), .A3(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n799), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n979), .B1(new_n790), .B2(new_n983), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n751), .B(new_n753), .C1(new_n583), .C2(new_n733), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n732), .A2(new_n570), .A3(new_n581), .A4(new_n687), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n731), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(KEYINPUT105), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1008), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(new_n730), .A3(new_n735), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n582), .B1(new_n1008), .B2(new_n676), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1016), .A2(KEYINPUT42), .B1(new_n733), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT42), .B2(new_n1016), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1011), .A2(KEYINPUT105), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1013), .A2(new_n1014), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1014), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1020), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n1023), .B2(new_n1012), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n781), .A2(G1), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n736), .A2(new_n734), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n1008), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1028), .B(new_n1029), .Z(new_n1030));
  NOR2_X1   g0830(.A1(new_n1027), .A2(new_n1008), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT45), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n726), .A3(new_n730), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n731), .A3(new_n1032), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n730), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n724), .B2(new_n725), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n731), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n722), .B2(new_n727), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n731), .A2(new_n735), .A3(new_n1038), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n778), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n739), .B(KEYINPUT41), .Z(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1026), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1005), .B1(new_n1025), .B2(new_n1046), .ZN(G387));
  OAI21_X1  g0847(.A(new_n269), .B1(new_n869), .B2(new_n814), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n823), .A2(G322), .B1(new_n819), .B2(G303), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n877), .B2(new_n825), .C1(new_n845), .C2(new_n1000), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT48), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT48), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n873), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n807), .A2(new_n1054), .B1(G294), .B2(new_n838), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(KEYINPUT109), .B(KEYINPUT49), .Z(new_n1057));
  XNOR2_X1  g0857(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1048), .B(new_n1058), .C1(G326), .C2(new_n836), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n807), .A2(new_n594), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G159), .A2(new_n823), .B1(new_n838), .B2(G77), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G50), .A2(new_n829), .B1(new_n826), .B2(new_n246), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n262), .A2(new_n818), .B1(new_n814), .B2(new_n546), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(new_n269), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n836), .B2(G150), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n799), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n803), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n232), .A2(G45), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n246), .A2(new_n202), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT50), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n742), .B(new_n503), .C1(new_n262), .C2(new_n369), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1069), .B(new_n797), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(G107), .B2(new_n210), .C1(new_n742), .C2(new_n792), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n782), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1067), .B(new_n1075), .C1(new_n730), .C2(new_n790), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1026), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n778), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n739), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1078), .A2(new_n778), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1076), .B1(new_n1042), .B2(new_n1077), .C1(new_n1080), .C2(new_n1081), .ZN(G393));
  INV_X1    g0882(.A(new_n1079), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1036), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n740), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1035), .B1(new_n1034), .B2(KEYINPUT110), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(KEYINPUT110), .B2(new_n1034), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1087), .B2(new_n1083), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1015), .A2(new_n790), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n836), .A2(G322), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n807), .A2(new_n485), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n278), .B1(new_n814), .B2(new_n398), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n825), .A2(new_n812), .B1(new_n818), .B2(new_n871), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(new_n838), .C2(new_n1054), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n822), .A2(new_n1000), .B1(new_n828), .B2(new_n877), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1090), .A2(new_n1091), .A3(new_n1094), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n836), .A2(G143), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n807), .A2(G77), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n822), .A2(new_n858), .B1(new_n828), .B2(new_n258), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT51), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n218), .A2(new_n811), .B1(new_n814), .B2(new_n634), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n825), .A2(new_n202), .B1(new_n818), .B2(new_n245), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1103), .A2(new_n1104), .A3(new_n269), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .A4(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n800), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n797), .A2(new_n243), .B1(G97), .B2(new_n738), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n782), .B(new_n1107), .C1(new_n802), .C2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1087), .A2(new_n1026), .B1(new_n1089), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT112), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1088), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n739), .B1(new_n1079), .B2(new_n1036), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1034), .A2(KEYINPUT110), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1034), .A2(KEYINPUT110), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n1035), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1113), .B1(new_n1116), .B2(new_n1079), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1089), .A2(new_n1109), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1116), .B2(new_n1077), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT112), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1112), .A2(new_n1120), .ZN(G390));
  NAND4_X1  g0921(.A1(new_n910), .A2(new_n897), .A3(G330), .A4(new_n883), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n955), .B1(new_n936), .B2(new_n924), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n888), .A2(new_n958), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n943), .B1(new_n1125), .B2(new_n910), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n924), .A2(new_n931), .A3(new_n955), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n882), .A2(new_n707), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n880), .B1(new_n755), .B2(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n908), .A2(new_n909), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n932), .B(new_n944), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1123), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT113), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n777), .A2(new_n1135), .A3(new_n883), .A4(new_n910), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n910), .A2(new_n776), .A3(G330), .A4(new_n883), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT113), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n888), .A2(new_n958), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n944), .B1(new_n1140), .B2(new_n1131), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n954), .A2(new_n1141), .A3(new_n956), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1139), .A2(new_n1142), .A3(new_n1132), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1134), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1026), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n788), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n954), .A2(new_n1146), .A3(new_n956), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n855), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n786), .B1(new_n246), .B2(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n836), .A2(G125), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT53), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n838), .B2(G150), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n278), .B(new_n1152), .C1(new_n819), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n807), .A2(G159), .ZN(new_n1156));
  INV_X1    g0956(.A(G128), .ZN(new_n1157));
  INV_X1    g0957(.A(G132), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n822), .A2(new_n1157), .B1(new_n828), .B2(new_n1158), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n825), .A2(new_n991), .B1(new_n814), .B2(new_n202), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n838), .A2(new_n1151), .A3(G150), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1155), .A2(new_n1156), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n835), .A2(new_n871), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n634), .A2(new_n811), .B1(new_n825), .B2(new_n398), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G283), .B2(new_n823), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n281), .B1(new_n840), .B2(G68), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G116), .A2(new_n829), .B1(new_n819), .B2(G97), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1100), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1150), .A2(new_n1163), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1149), .B1(new_n1170), .B2(new_n799), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1147), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1145), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT114), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n465), .A2(new_n469), .A3(KEYINPUT81), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n475), .B1(new_n474), .B2(new_n476), .ZN(new_n1177));
  OAI211_X1 g0977(.A(G330), .B(new_n897), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n897), .A2(G330), .A3(new_n883), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n1131), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n1130), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1131), .B1(new_n890), .B2(new_n886), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1140), .B1(new_n1183), .B2(new_n1122), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n964), .B(new_n1178), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1134), .A2(new_n1143), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1175), .B(new_n739), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1181), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1184), .B1(new_n1139), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n478), .A2(new_n756), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1178), .A2(new_n1190), .A3(new_n712), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1187), .B1(new_n1144), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1144), .A2(new_n1192), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1175), .B1(new_n1194), .B2(new_n739), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1174), .B1(new_n1193), .B2(new_n1195), .ZN(G378));
  OAI21_X1  g0996(.A(new_n943), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n937), .A2(new_n959), .B1(new_n705), .B2(new_n717), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n382), .A2(new_n417), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n362), .A2(new_n717), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  XOR2_X1   g1001(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1202));
  XOR2_X1   g1002(.A(new_n1201), .B(new_n1202), .Z(new_n1203));
  AND3_X1   g1003(.A1(new_n1197), .A2(new_n1198), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT40), .B1(new_n911), .B2(new_n937), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n932), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n910), .A2(new_n897), .A3(KEYINPUT40), .A4(new_n883), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1205), .A2(new_n1208), .A3(new_n725), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1203), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1204), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(G330), .B(new_n933), .C1(new_n938), .C2(KEYINPUT40), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1203), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n957), .B2(new_n962), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1197), .A2(new_n1198), .A3(new_n1203), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1212), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1026), .B1(new_n1211), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1203), .A2(new_n1146), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n786), .B1(G50), .B2(new_n1148), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n369), .A2(new_n811), .B1(new_n828), .B2(new_n398), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n825), .A2(new_n546), .B1(new_n818), .B2(new_n391), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n822), .A2(new_n481), .B1(new_n814), .B2(new_n985), .ZN(new_n1222));
  INV_X1    g1022(.A(G41), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n269), .A2(new_n1223), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n990), .C1(new_n835), .C2(new_n815), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT58), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G33), .A2(G41), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT115), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G50), .B(new_n1229), .C1(new_n1223), .C2(new_n269), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT116), .Z(new_n1231));
  AOI22_X1  g1031(.A1(G132), .A2(new_n826), .B1(new_n838), .B2(new_n1154), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1157), .B2(new_n828), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n823), .A2(G125), .B1(new_n819), .B2(G137), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n858), .C2(new_n876), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1229), .B1(new_n258), .B2(new_n814), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n836), .B2(G124), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1227), .B(new_n1231), .C1(new_n1237), .C2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1219), .B1(new_n1242), .B2(new_n799), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1218), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1217), .A2(KEYINPUT117), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT117), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1209), .B1(new_n1204), .B2(new_n1210), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1214), .A2(new_n1212), .A3(new_n1215), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1077), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1244), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1246), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1245), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT118), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1191), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n964), .A2(KEYINPUT118), .A3(new_n1178), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1144), .A2(new_n1192), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT57), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n964), .A2(KEYINPUT118), .A3(new_n1178), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT118), .B1(new_n964), .B2(new_n1178), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1185), .A2(new_n1186), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT57), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1258), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1252), .B1(new_n1265), .B2(new_n739), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(G375));
  OAI22_X1  g1067(.A1(new_n835), .A2(new_n812), .B1(new_n546), .B2(new_n811), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(KEYINPUT120), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n822), .A2(new_n871), .B1(new_n828), .B2(new_n815), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n281), .B(new_n1270), .C1(G77), .C2(new_n840), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n485), .A2(new_n826), .B1(new_n819), .B2(G107), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT119), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1272), .A2(KEYINPUT119), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1271), .A2(new_n1060), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(G159), .A2(new_n838), .B1(new_n840), .B2(G58), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1277), .B1(new_n1158), .B2(new_n822), .C1(new_n825), .C2(new_n1153), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n269), .B(new_n1278), .C1(G137), .C2(new_n846), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n807), .A2(G50), .B1(G150), .B2(new_n819), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT121), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1279), .B(new_n1281), .C1(new_n1157), .C2(new_n835), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1276), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT122), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n799), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1283), .A2(KEYINPUT122), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n786), .B1(G68), .B2(new_n1148), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n787), .B2(new_n1131), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1189), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(new_n1026), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1185), .A2(new_n1045), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1290), .B1(new_n1291), .B2(new_n1292), .ZN(G381));
  INV_X1    g1093(.A(new_n1046), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1112), .A2(new_n1120), .A3(new_n1295), .A4(new_n1005), .ZN(new_n1296));
  OR2_X1    g1096(.A1(G393), .A2(G396), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(new_n1296), .A2(G384), .A3(G381), .A4(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(G375), .A2(G378), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(G407));
  INV_X1    g1100(.A(G343), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(G213), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(KEYINPUT123), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(G407), .A2(G213), .A3(new_n1304), .ZN(G409));
  AOI21_X1  g1105(.A(new_n1111), .B1(new_n1088), .B2(new_n1110), .ZN(new_n1306));
  NOR3_X1   g1106(.A1(new_n1117), .A2(new_n1119), .A3(KEYINPUT112), .ZN(new_n1307));
  OAI21_X1  g1107(.A(G387), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1296), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(G393), .B(new_n853), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1310), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1308), .A2(new_n1296), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT125), .B1(new_n1217), .B2(new_n1244), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1256), .A2(new_n1257), .A3(new_n1044), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1217), .A2(KEYINPUT125), .A3(new_n1244), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G378), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT124), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1266), .B2(G378), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1262), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n739), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1245), .A2(new_n1251), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1325), .A2(new_n1326), .A3(G378), .A4(new_n1321), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1320), .B1(new_n1322), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1303), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT60), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1292), .A2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1292), .A2(new_n1332), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n739), .B(new_n1185), .C1(new_n1333), .C2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1290), .ZN(new_n1336));
  INV_X1    g1136(.A(G384), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1335), .A2(G384), .A3(new_n1290), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .A4(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1303), .A2(G2897), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1340), .A2(new_n1343), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1338), .A2(G2897), .A3(new_n1303), .A4(new_n1339), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1325), .A2(new_n1326), .A3(G378), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(KEYINPUT124), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1319), .B1(new_n1348), .B2(new_n1327), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1346), .B1(new_n1349), .B2(new_n1303), .ZN(new_n1350));
  XOR2_X1   g1150(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1351));
  NAND3_X1  g1151(.A1(new_n1342), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1349), .A2(new_n1303), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1330), .B1(new_n1353), .B2(new_n1341), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1314), .B1(new_n1352), .B2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT126), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1329), .A2(new_n1356), .A3(new_n1331), .ZN(new_n1357));
  OAI21_X1  g1157(.A(KEYINPUT126), .B1(new_n1349), .B2(new_n1303), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1357), .A2(new_n1358), .A3(new_n1346), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1329), .A2(new_n1331), .A3(new_n1341), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT63), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1353), .A2(KEYINPUT63), .A3(new_n1341), .ZN(new_n1363));
  AND3_X1   g1163(.A1(new_n1308), .A2(new_n1296), .A3(new_n1312), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1312), .B1(new_n1308), .B2(new_n1296), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1364), .A2(new_n1365), .A3(KEYINPUT61), .ZN(new_n1366));
  NAND4_X1  g1166(.A1(new_n1359), .A2(new_n1362), .A3(new_n1363), .A4(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1355), .A2(new_n1367), .ZN(G405));
  OAI21_X1  g1168(.A(new_n1340), .B1(new_n1364), .B2(new_n1365), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1311), .A2(new_n1313), .A3(new_n1341), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  INV_X1    g1171(.A(G378), .ZN(new_n1372));
  AOI22_X1  g1172(.A1(new_n1348), .A2(new_n1327), .B1(G375), .B2(new_n1372), .ZN(new_n1373));
  XNOR2_X1  g1173(.A(new_n1371), .B(new_n1373), .ZN(G402));
endmodule


