//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  XNOR2_X1  g002(.A(G125), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT74), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT74), .A3(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(KEYINPUT16), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n192), .B2(G140), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n188), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT67), .A2(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT67), .A2(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G119), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(G119), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n202), .A2(new_n205), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n204), .B1(new_n201), .B2(G119), .ZN(new_n211));
  XOR2_X1   g025(.A(KEYINPUT24), .B(G110), .Z(new_n212));
  OAI22_X1  g026(.A1(new_n210), .A2(G110), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n189), .A2(new_n188), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n198), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n210), .A2(G110), .B1(new_n211), .B2(new_n212), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n194), .A2(new_n188), .A3(new_n196), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(new_n197), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G137), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n220), .B(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n215), .A2(new_n218), .A3(new_n223), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n187), .B1(new_n227), .B2(G902), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n225), .A2(KEYINPUT25), .A3(new_n229), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G217), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(G234), .B2(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(G902), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n227), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(KEYINPUT75), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT75), .ZN(new_n240));
  INV_X1    g054(.A(new_n233), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n228), .B2(new_n230), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n240), .B1(new_n242), .B2(new_n237), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G119), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT68), .A2(G116), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT68), .A2(G116), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n246), .B1(new_n249), .B2(G119), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT2), .B(G113), .Z(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OR2_X1    g066(.A1(KEYINPUT68), .A2(G116), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT68), .A2(G116), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(G119), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n246), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n250), .A2(KEYINPUT69), .A3(new_n251), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n252), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT11), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(G137), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT11), .A3(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(G137), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G131), .ZN(new_n270));
  INV_X1    g084(.A(G131), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n265), .A2(new_n267), .A3(new_n271), .A4(new_n268), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(KEYINPUT66), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT0), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(new_n203), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT64), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(KEYINPUT0), .B2(G128), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n203), .A3(KEYINPUT64), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n280));
  INV_X1    g094(.A(G143), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(G146), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n188), .A2(KEYINPUT65), .A3(G143), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G143), .B(G146), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n279), .A2(new_n285), .B1(new_n275), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n269), .A2(new_n288), .A3(G131), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n273), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n268), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n264), .A2(G137), .ZN(new_n292));
  OAI21_X1  g106(.A(G131), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n293), .A2(new_n272), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n203), .A2(KEYINPUT1), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n286), .A2(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n297));
  OR2_X1    g111(.A1(KEYINPUT67), .A2(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(KEYINPUT67), .A2(G128), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n188), .A2(G143), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(KEYINPUT1), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n296), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n294), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n290), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n262), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT72), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(KEYINPUT70), .B(new_n296), .C1(new_n297), .C2(new_n301), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n294), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n261), .A3(new_n290), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT71), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n310), .A2(new_n313), .A3(new_n261), .A4(new_n290), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n262), .A2(new_n304), .A3(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n306), .A2(new_n312), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT28), .ZN(new_n318));
  INV_X1    g132(.A(new_n311), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT28), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G237), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n221), .A3(G210), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT27), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G101), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n310), .A2(KEYINPUT30), .A3(new_n290), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT30), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n304), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n331), .A3(new_n262), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n332), .A2(new_n312), .A3(new_n314), .A4(new_n327), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT31), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n312), .A2(new_n314), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n336), .A2(KEYINPUT31), .A3(new_n327), .A4(new_n332), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n322), .A2(new_n328), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(G472), .A2(G902), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT32), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n335), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n333), .A2(new_n334), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n320), .B1(new_n317), .B2(KEYINPUT28), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n342), .A2(new_n343), .B1(new_n344), .B2(new_n327), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n339), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n336), .A2(new_n328), .A3(new_n332), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n344), .B2(new_n328), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n310), .A2(new_n290), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n262), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n312), .A2(new_n354), .A3(new_n314), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT28), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n328), .A2(new_n351), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n321), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n229), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n352), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G472), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n244), .B1(new_n348), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G210), .B1(G237), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(G101), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(new_n367), .B2(G107), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n369));
  INV_X1    g183(.A(G107), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G104), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(G107), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n366), .A2(new_n368), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n372), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n367), .A2(G107), .ZN(new_n375));
  OAI21_X1  g189(.A(G101), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G113), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT5), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n246), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n255), .A2(new_n256), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(new_n380), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT69), .B1(new_n250), .B2(new_n251), .ZN(new_n384));
  AND4_X1   g198(.A1(KEYINPUT69), .A2(new_n251), .A3(new_n255), .A4(new_n256), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n378), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n368), .A2(new_n371), .A3(new_n372), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G101), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n387), .B1(new_n389), .B2(new_n373), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT4), .B1(new_n388), .B2(G101), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n386), .B1(new_n261), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G122), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n386), .B(new_n394), .C1(new_n261), .C2(new_n392), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(KEYINPUT6), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n393), .A2(new_n399), .A3(new_n395), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n287), .A2(G125), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n302), .A2(new_n192), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT82), .B(G224), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n221), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n398), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(KEYINPUT7), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n409), .A2(KEYINPUT83), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(KEYINPUT83), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n403), .A2(KEYINPUT7), .A3(new_n405), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n394), .B(KEYINPUT8), .ZN(new_n414));
  INV_X1    g228(.A(new_n386), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n260), .A2(new_n259), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n378), .B1(new_n416), .B2(new_n383), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n414), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n397), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n229), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n365), .B1(new_n407), .B2(new_n420), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n413), .A2(new_n419), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n398), .A2(new_n400), .A3(new_n406), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n229), .A4(new_n364), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G214), .B1(G237), .B2(G902), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n373), .A2(KEYINPUT10), .A3(new_n376), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n308), .A2(new_n309), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n287), .B1(new_n390), .B2(new_n391), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n273), .A2(new_n289), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n300), .A2(KEYINPUT1), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n286), .B1(G128), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n286), .A2(new_n295), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n373), .B(new_n376), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT10), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n430), .A2(new_n431), .A3(new_n432), .A4(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  INV_X1    g254(.A(G227), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G953), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n440), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n439), .A2(KEYINPUT80), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT80), .B1(new_n439), .B2(new_n444), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n298), .A2(new_n299), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n433), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n285), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n377), .A2(new_n449), .A3(new_n296), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n450), .A2(new_n436), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT79), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n273), .A2(new_n452), .A3(new_n289), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT12), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n436), .ZN(new_n455));
  INV_X1    g269(.A(new_n432), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n452), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n445), .A2(new_n446), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n430), .A2(new_n431), .A3(new_n438), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n456), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n444), .B1(new_n462), .B2(new_n439), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n428), .B(new_n229), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(G469), .A2(G902), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n454), .A2(new_n439), .A3(new_n458), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n443), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n462), .A2(new_n439), .A3(new_n444), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(G469), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT9), .B(G234), .ZN(new_n471));
  OAI21_X1  g285(.A(G221), .B1(new_n471), .B2(G902), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT76), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n473), .B(KEYINPUT77), .Z(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT81), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n470), .A2(KEYINPUT81), .A3(new_n475), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n427), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n471), .A2(new_n232), .A3(G953), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n281), .A2(G128), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT88), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n201), .B2(G143), .ZN(new_n485));
  NOR4_X1   g299(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT90), .A4(new_n281), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT89), .B(KEYINPUT13), .Z(new_n488));
  NAND3_X1  g302(.A1(new_n298), .A2(G143), .A3(new_n299), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT90), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n298), .A2(new_n484), .A3(G143), .A4(new_n299), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n487), .B1(new_n492), .B2(new_n264), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n491), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n494), .A2(G134), .A3(new_n483), .A4(new_n488), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G122), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n247), .A2(new_n248), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n245), .A2(G122), .ZN(new_n499));
  OAI21_X1  g313(.A(G107), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n253), .A2(G122), .A3(new_n254), .ZN(new_n501));
  INV_X1    g315(.A(new_n499), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n370), .A3(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n500), .A2(KEYINPUT87), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT87), .B1(new_n500), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n496), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT91), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n496), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n501), .B1(KEYINPUT14), .B2(new_n499), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n512), .A2(KEYINPUT92), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n512), .B(KEYINPUT92), .C1(KEYINPUT14), .C2(new_n501), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(G107), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n487), .A2(new_n264), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n494), .A2(G134), .A3(new_n483), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n515), .A2(new_n503), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n481), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n496), .A2(new_n509), .A3(new_n506), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n509), .B1(new_n496), .B2(new_n506), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n518), .B(new_n481), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n229), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT93), .ZN(new_n525));
  INV_X1    g339(.A(G478), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n532));
  INV_X1    g346(.A(new_n481), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n522), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n229), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n525), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(G113), .B(G122), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(new_n367), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n323), .A2(new_n221), .A3(G214), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n281), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n323), .A2(new_n221), .A3(G143), .A4(G214), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT85), .B1(new_n545), .B2(new_n271), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT85), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n547), .A3(G131), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n271), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT84), .B1(new_n191), .B2(new_n193), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n191), .A2(KEYINPUT84), .A3(new_n193), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(KEYINPUT19), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT19), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n189), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n198), .B(new_n550), .C1(new_n557), .C2(G146), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n552), .A2(G146), .A3(new_n553), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n214), .ZN(new_n560));
  NAND2_X1  g374(.A1(KEYINPUT18), .A2(G131), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n544), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n540), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n546), .A2(new_n548), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT86), .B1(new_n565), .B2(KEYINPUT17), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT86), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n568));
  AOI211_X1 g382(.A(new_n567), .B(new_n568), .C1(new_n546), .C2(new_n548), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n217), .A2(new_n197), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n546), .A2(new_n568), .A3(new_n548), .A4(new_n549), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n570), .A2(new_n573), .B1(new_n560), .B2(new_n562), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n564), .B1(new_n574), .B2(new_n540), .ZN(new_n575));
  NOR2_X1   g389(.A1(G475), .A2(G902), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT20), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n566), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n565), .A2(KEYINPUT86), .A3(KEYINPUT17), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n573), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n540), .A3(new_n563), .ZN(new_n582));
  INV_X1    g396(.A(new_n564), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT20), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n576), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n581), .A2(new_n540), .A3(new_n563), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n540), .B1(new_n581), .B2(new_n563), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n229), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n578), .A2(new_n586), .B1(new_n589), .B2(G475), .ZN(new_n590));
  INV_X1    g404(.A(G952), .ZN(new_n591));
  AOI211_X1 g405(.A(G953), .B(new_n591), .C1(G234), .C2(G237), .ZN(new_n592));
  AOI211_X1 g406(.A(new_n229), .B(new_n221), .C1(G234), .C2(G237), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT21), .B(G898), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n524), .A2(new_n531), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n538), .A2(new_n590), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n363), .A2(new_n480), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n366), .ZN(G3));
  NAND2_X1  g416(.A1(new_n578), .A2(new_n586), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n589), .A2(G475), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n427), .A2(new_n595), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n607));
  INV_X1    g421(.A(new_n518), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n508), .B2(new_n510), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n607), .B1(new_n609), .B2(new_n481), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n535), .A2(KEYINPUT33), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n534), .B(new_n522), .C1(new_n607), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n526), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n525), .A2(new_n526), .A3(new_n537), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n616), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n611), .B2(new_n613), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n615), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n605), .B(new_n606), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n345), .A2(new_n229), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n624), .A2(G472), .B1(new_n345), .B2(new_n339), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n239), .A2(new_n243), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n470), .A2(KEYINPUT81), .A3(new_n475), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT81), .B1(new_n470), .B2(new_n475), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NAND2_X1  g446(.A1(new_n538), .A2(new_n598), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n606), .A2(new_n633), .A3(new_n590), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n625), .A2(new_n626), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n478), .A2(new_n479), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n219), .A2(KEYINPUT97), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n215), .A2(new_n218), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(KEYINPUT36), .B2(new_n224), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n641), .A2(new_n646), .A3(new_n643), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n645), .A2(new_n235), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n640), .B1(new_n649), .B2(new_n242), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n234), .A2(KEYINPUT98), .A3(new_n648), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n480), .A2(new_n600), .A3(new_n625), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT37), .B(G110), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT99), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n654), .B(new_n656), .ZN(G12));
  INV_X1    g471(.A(new_n426), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n421), .B2(new_n424), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n659), .B1(new_n627), .B2(new_n628), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n341), .A2(new_n347), .B1(new_n361), .B2(G472), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n592), .B1(new_n593), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n633), .A2(new_n663), .A3(new_n590), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n633), .A2(new_n590), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT100), .B1(new_n668), .B2(new_n665), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n662), .A2(new_n653), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  NAND2_X1  g485(.A1(new_n355), .A2(new_n328), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n333), .ZN(new_n673));
  AOI21_X1  g487(.A(G902), .B1(new_n673), .B2(KEYINPUT101), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(KEYINPUT101), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G472), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n348), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n425), .B(KEYINPUT38), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n633), .A2(new_n605), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n649), .A2(new_n242), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n426), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n678), .A2(new_n679), .A3(new_n680), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n665), .B(KEYINPUT39), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n636), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT102), .B(G143), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G45));
  OAI211_X1 g504(.A(new_n605), .B(new_n666), .C1(new_n619), .C2(new_n622), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT103), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n614), .A2(new_n616), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT96), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n617), .A3(new_n618), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n605), .A4(new_n666), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n692), .A2(new_n697), .A3(new_n653), .A4(new_n662), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  AOI21_X1  g513(.A(new_n536), .B1(new_n535), .B2(new_n229), .ZN(new_n700));
  AOI211_X1 g514(.A(KEYINPUT93), .B(G902), .C1(new_n534), .C2(new_n522), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n526), .A2(new_n702), .B1(new_n621), .B2(new_n615), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n590), .B1(new_n703), .B2(new_n694), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n446), .A2(new_n459), .ZN(new_n705));
  INV_X1    g519(.A(new_n445), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n463), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(G469), .B1(new_n707), .B2(G902), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n464), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n473), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n704), .A2(new_n363), .A3(new_n606), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND3_X1  g530(.A1(new_n634), .A2(new_n363), .A3(new_n713), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  INV_X1    g532(.A(new_n473), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n711), .A2(new_n719), .A3(new_n659), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n599), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n338), .A2(KEYINPUT32), .A3(new_n340), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n346), .B1(new_n345), .B2(new_n339), .ZN(new_n723));
  INV_X1    g537(.A(G472), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n359), .B1(new_n350), .B2(new_n351), .ZN(new_n725));
  OAI22_X1  g539(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n721), .A2(new_n726), .A3(new_n653), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  AND4_X1   g542(.A1(new_n596), .A2(new_n708), .A3(new_n464), .A4(new_n719), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n605), .A2(new_n633), .A3(new_n659), .A4(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n724), .B1(new_n345), .B2(new_n229), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n356), .A2(new_n321), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n328), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n337), .A2(new_n335), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n340), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n242), .A2(new_n237), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n730), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  NOR3_X1   g554(.A1(new_n731), .A2(new_n681), .A3(new_n735), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n720), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n692), .A2(new_n697), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n692), .A2(new_n746), .A3(new_n697), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n465), .B(KEYINPUT104), .Z(new_n748));
  NAND3_X1  g562(.A1(new_n464), .A2(new_n469), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n719), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(KEYINPUT105), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n749), .B2(new_n719), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n421), .A2(new_n426), .A3(new_n424), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n363), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n726), .A2(new_n737), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n751), .A2(new_n754), .A3(new_n755), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n692), .A2(new_n697), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n747), .A2(new_n757), .B1(new_n760), .B2(KEYINPUT42), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n757), .A2(new_n763), .A3(new_n667), .A4(new_n669), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n669), .A2(new_n759), .A3(new_n363), .A4(new_n667), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT106), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  NAND2_X1  g582(.A1(new_n695), .A2(new_n590), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n625), .A2(new_n681), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n755), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n774), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n467), .A2(new_n468), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(KEYINPUT45), .ZN(new_n779));
  OAI21_X1  g593(.A(G469), .B1(new_n778), .B2(KEYINPUT45), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n782), .B2(new_n748), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n710), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n748), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n786), .A2(new_n719), .A3(new_n684), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n719), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT47), .Z(new_n791));
  NOR3_X1   g605(.A1(new_n726), .A2(new_n626), .A3(new_n755), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n692), .A2(new_n697), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT107), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NAND2_X1  g612(.A1(new_n712), .A2(KEYINPUT49), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n474), .A2(new_n658), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n799), .A2(new_n679), .A3(new_n737), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n712), .A2(KEYINPUT49), .ZN(new_n802));
  OR4_X1    g616(.A1(new_n677), .A2(new_n801), .A3(new_n769), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n680), .A2(new_n427), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n681), .A2(new_n666), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT112), .ZN(new_n807));
  INV_X1    g621(.A(new_n750), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n805), .A2(new_n807), .A3(new_n677), .A4(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n698), .A2(new_n744), .A3(new_n670), .A4(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(KEYINPUT52), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(KEYINPUT52), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n804), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n744), .A2(new_n670), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n698), .A4(new_n809), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n810), .A2(KEYINPUT52), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(KEYINPUT113), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n752), .A2(new_n756), .A3(new_n741), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n692), .A2(new_n820), .A3(new_n697), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT111), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n692), .A2(new_n820), .A3(new_n697), .A4(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n822), .A2(new_n824), .B1(new_n764), .B2(new_n766), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT108), .B1(new_n601), .B2(new_n630), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n363), .A2(new_n480), .A3(new_n600), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT108), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n827), .B(new_n828), .C1(new_n623), .C2(new_n629), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n637), .A2(new_n654), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n826), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n714), .A2(new_n717), .A3(new_n727), .A4(new_n739), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n636), .A2(new_n726), .A3(new_n653), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n426), .A2(new_n421), .A3(new_n424), .A4(new_n666), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n538), .A3(new_n590), .A4(new_n598), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT109), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n597), .B1(new_n702), .B2(new_n531), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(KEYINPUT109), .A3(new_n590), .A4(new_n834), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n833), .A2(KEYINPUT110), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT110), .B1(new_n833), .B2(new_n840), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n832), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n825), .A2(new_n831), .A3(new_n843), .A4(new_n761), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n819), .A2(KEYINPUT114), .A3(KEYINPUT53), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n847), .B(new_n844), .C1(new_n813), .C2(new_n818), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n816), .A2(new_n817), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n846), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n712), .A2(new_n473), .A3(new_n755), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n770), .A2(new_n592), .A3(new_n771), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n742), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n626), .A2(new_n592), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n678), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n861), .A2(new_n605), .A3(new_n695), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n713), .A2(new_n658), .A3(new_n679), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT117), .Z(new_n864));
  NAND4_X1  g678(.A1(new_n770), .A2(new_n592), .A3(new_n738), .A4(new_n771), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT50), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n866), .B1(new_n864), .B2(new_n865), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n858), .B(new_n862), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n865), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n474), .B1(new_n711), .B2(KEYINPUT115), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(KEYINPUT115), .B2(new_n711), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n870), .B(new_n776), .C1(new_n791), .C2(new_n872), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n869), .B(new_n873), .C1(KEYINPUT116), .C2(KEYINPUT51), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n858), .A2(new_n862), .ZN(new_n875));
  INV_X1    g689(.A(new_n868), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n873), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  OAI211_X1 g693(.A(KEYINPUT116), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n758), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n857), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT48), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n591), .B(G953), .C1(new_n860), .C2(new_n704), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n720), .B2(new_n865), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n874), .A2(new_n881), .A3(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n845), .A2(KEYINPUT53), .A3(new_n816), .A4(new_n817), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n844), .B1(new_n813), .B2(new_n818), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(KEYINPUT53), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n855), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(G952), .A2(G953), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n803), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(KEYINPUT118), .B(new_n803), .C1(new_n893), .C2(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(G75));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  INV_X1    g714(.A(new_n853), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(G902), .ZN(new_n902));
  INV_X1    g716(.A(G210), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n398), .A2(new_n400), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(new_n406), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(KEYINPUT56), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n221), .A2(G952), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n904), .B2(new_n909), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n910), .A2(new_n913), .ZN(G51));
  NOR2_X1   g728(.A1(new_n902), .A2(new_n782), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n846), .B(KEYINPUT54), .C1(new_n848), .C2(new_n852), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n855), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n748), .B(KEYINPUT57), .Z(new_n918));
  AOI21_X1  g732(.A(new_n707), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n919), .B2(KEYINPUT120), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n921));
  INV_X1    g735(.A(new_n918), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n855), .B2(new_n916), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n923), .B2(new_n707), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n911), .B1(new_n920), .B2(new_n924), .ZN(G54));
  AND4_X1   g739(.A1(KEYINPUT58), .A2(new_n901), .A3(G475), .A4(G902), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n912), .B1(new_n926), .B2(new_n584), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n584), .B2(new_n926), .ZN(G60));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n855), .B2(new_n892), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n912), .B1(new_n931), .B2(new_n614), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n611), .B2(new_n613), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n917), .A2(KEYINPUT121), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n917), .A2(new_n933), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n932), .B1(new_n934), .B2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n853), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n227), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n645), .A2(new_n647), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n942), .B(new_n912), .C1(new_n943), .C2(new_n941), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n911), .B1(new_n941), .B2(new_n227), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n947), .B(KEYINPUT61), .C1(new_n943), .C2(new_n941), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n594), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n221), .B1(new_n950), .B2(new_n404), .ZN(new_n951));
  INV_X1    g765(.A(new_n832), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n831), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n953), .B2(new_n221), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n905), .B1(G898), .B2(new_n221), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT122), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  XOR2_X1   g771(.A(new_n557), .B(KEYINPUT123), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n329), .A2(new_n331), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n814), .A2(new_n698), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n688), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT62), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n838), .A2(new_n605), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n363), .B(new_n776), .C1(new_n704), .C2(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n797), .B(new_n788), .C1(new_n685), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(G953), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n221), .A2(G900), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n787), .A2(new_n805), .A3(new_n758), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT126), .Z(new_n971));
  AND3_X1   g785(.A1(new_n971), .A2(new_n761), .A3(new_n767), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT125), .B1(new_n788), .B2(new_n961), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n788), .A2(KEYINPUT125), .A3(new_n961), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n972), .B(new_n797), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n969), .B1(new_n975), .B2(new_n221), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n968), .B1(new_n976), .B2(new_n960), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n441), .B2(new_n664), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT124), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n977), .B(new_n979), .ZN(G72));
  NAND2_X1  g794(.A1(new_n336), .A2(new_n332), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n327), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n967), .A2(new_n831), .A3(new_n952), .ZN(new_n983));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n982), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n987), .B2(new_n986), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n985), .B1(new_n975), .B2(new_n953), .ZN(new_n990));
  INV_X1    g804(.A(new_n349), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n911), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n891), .A2(new_n349), .A3(new_n982), .A4(new_n985), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n989), .A2(new_n992), .A3(new_n993), .ZN(G57));
endmodule


