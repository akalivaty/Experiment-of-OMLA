//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT92), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(new_n205), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G43gat), .B(G50gat), .Z(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n212), .A2(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT91), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT91), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT14), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n219), .A2(KEYINPUT14), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n214), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n212), .A2(new_n213), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n223), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n225), .A2(new_n214), .A3(new_n220), .A4(new_n221), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n226), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n209), .B(G8gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n229), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n202), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G169gat), .B(G197gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT12), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n211), .A2(new_n227), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n235), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n233), .B(KEYINPUT13), .Z(new_n248));
  AOI22_X1  g047(.A1(new_n236), .A2(new_n237), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n232), .A2(new_n235), .A3(KEYINPUT18), .A4(new_n233), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n249), .B(new_n250), .C1(new_n238), .C2(new_n244), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT94), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT94), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(G211gat), .B(G218gat), .Z(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n260));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT22), .ZN(new_n262));
  INV_X1    g061(.A(G211gat), .ZN(new_n263));
  INV_X1    g062(.A(G218gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n260), .B(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G226gat), .ZN(new_n268));
  INV_X1    g067(.A(G233gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT26), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G183gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT27), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT27), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G183gat), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT66), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(KEYINPUT66), .A3(KEYINPUT28), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n279), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n273), .A2(KEYINPUT24), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI211_X1 g096(.A(KEYINPUT65), .B(new_n291), .C1(new_n292), .C2(new_n294), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n271), .A2(KEYINPUT23), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n297), .A2(new_n298), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n292), .A2(new_n294), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT64), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n299), .A2(new_n302), .A3(new_n301), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT25), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n290), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n270), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n270), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n310), .B(KEYINPUT25), .C1(new_n296), .C2(new_n295), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n302), .A3(new_n301), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n308), .A2(new_n306), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(new_n305), .ZN(new_n319));
  OAI22_X1  g118(.A1(new_n316), .A2(new_n298), .B1(new_n319), .B2(KEYINPUT25), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n315), .B1(new_n320), .B2(new_n290), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n267), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n312), .A2(new_n270), .ZN(new_n323));
  INV_X1    g122(.A(new_n267), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT29), .B1(new_n320), .B2(new_n290), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n270), .ZN(new_n326));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT71), .ZN(new_n328));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n322), .A2(KEYINPUT30), .A3(new_n326), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT72), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n322), .A2(new_n330), .A3(new_n326), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n322), .A2(new_n326), .ZN(new_n337));
  INV_X1    g136(.A(new_n330), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342));
  INV_X1    g141(.A(G155gat), .ZN(new_n343));
  INV_X1    g142(.A(G162gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  INV_X1    g145(.A(G148gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(G141gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n345), .A2(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G141gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G148gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(G141gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT73), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n351), .A2(G148gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n342), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G155gat), .B(G162gat), .Z(new_n357));
  AOI22_X1  g156(.A1(new_n350), .A2(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359));
  AND2_X1   g158(.A1(G113gat), .A2(G120gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(G113gat), .A2(G120gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(G127gat), .A2(G134gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(G127gat), .A2(G134gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT67), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n359), .B(new_n362), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G113gat), .ZN(new_n368));
  INV_X1    g167(.A(G120gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G113gat), .A2(G120gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n359), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n366), .A3(new_n371), .ZN(new_n373));
  XNOR2_X1  g172(.A(G127gat), .B(G134gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n358), .A2(new_n376), .A3(KEYINPUT75), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT75), .B1(new_n358), .B2(new_n376), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT74), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n356), .A2(new_n357), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n345), .A2(new_n346), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n348), .A2(new_n349), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n354), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n384), .B1(new_n389), .B2(KEYINPUT3), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n358), .A2(KEYINPUT74), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n376), .B1(new_n389), .B2(KEYINPUT3), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n383), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n358), .A2(new_n376), .A3(KEYINPUT4), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n367), .A2(new_n375), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(new_n389), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n358), .A2(new_n376), .A3(KEYINPUT75), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n389), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n398), .B1(new_n404), .B2(new_n383), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT76), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(new_n406), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n397), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT4), .B1(new_n377), .B2(new_n378), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n380), .B1(new_n400), .B2(new_n389), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n395), .A2(new_n398), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT0), .ZN(new_n415));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT77), .B1(new_n413), .B2(new_n418), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT77), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n409), .A2(new_n423), .A3(new_n417), .A4(new_n412), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n419), .A2(new_n420), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n341), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT89), .ZN(new_n428));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429));
  INV_X1    g228(.A(G50gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G22gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n393), .A2(new_n313), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n324), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n393), .A2(KEYINPUT80), .A3(new_n313), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n391), .B1(new_n267), .B2(KEYINPUT29), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n389), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(G228gat), .A3(G233gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n433), .A2(new_n267), .ZN(new_n443));
  INV_X1    g242(.A(new_n266), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n444), .A2(new_n259), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n313), .B1(new_n444), .B2(new_n259), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n391), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n389), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n443), .A2(new_n448), .B1(G228gat), .B2(G233gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n432), .B1(new_n442), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n440), .B1(new_n436), .B2(new_n435), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n452), .A2(G22gat), .A3(new_n449), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n431), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n442), .A2(new_n450), .A3(new_n432), .ZN(new_n455));
  OAI21_X1  g254(.A(G22gat), .B1(new_n452), .B2(new_n449), .ZN(new_n456));
  INV_X1    g255(.A(new_n431), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n454), .A2(new_n460), .A3(new_n458), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT34), .ZN(new_n465));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(KEYINPUT69), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n312), .A2(new_n376), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n320), .A2(new_n400), .A3(new_n290), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n468), .B1(new_n471), .B2(new_n466), .ZN(new_n472));
  INV_X1    g271(.A(new_n466), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n473), .B(new_n467), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n473), .A3(new_n470), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT33), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G43gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT68), .ZN(new_n480));
  INV_X1    g279(.A(G71gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G99gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n476), .A2(KEYINPUT32), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n478), .B(new_n484), .C1(new_n472), .C2(new_n474), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n486), .B2(new_n489), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n428), .B1(new_n464), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n462), .A2(new_n493), .A3(KEYINPUT89), .A4(new_n463), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n427), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n464), .A2(new_n494), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n417), .B1(new_n409), .B2(new_n412), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n502));
  INV_X1    g301(.A(new_n420), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n501), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n422), .A2(new_n424), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n501), .A2(new_n503), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT81), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n333), .B2(new_n340), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n336), .A2(new_n339), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n513), .B(KEYINPUT81), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n519));
  NAND3_X1  g318(.A1(new_n510), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI22_X1  g319(.A1(new_n497), .A2(new_n498), .B1(new_n500), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT40), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT74), .B1(new_n358), .B2(new_n391), .ZN(new_n523));
  AND4_X1   g322(.A1(KEYINPUT74), .A2(new_n385), .A3(new_n388), .A4(new_n391), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n394), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n410), .A2(new_n525), .A3(new_n411), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n526), .A2(KEYINPUT82), .A3(new_n383), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT82), .B1(new_n526), .B2(new_n383), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n379), .A2(new_n382), .A3(new_n403), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT39), .B1(new_n530), .B2(KEYINPUT84), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(KEYINPUT84), .B2(new_n530), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n522), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT39), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n527), .B2(new_n528), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT83), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n535), .A2(new_n536), .A3(new_n417), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n535), .B2(new_n417), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n539), .A2(new_n512), .A3(new_n516), .A4(new_n419), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n526), .A2(new_n383), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT82), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n526), .A2(KEYINPUT82), .A3(new_n383), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT39), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT83), .B1(new_n545), .B2(new_n418), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n535), .A2(new_n536), .A3(new_n417), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n532), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT40), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT85), .B1(new_n540), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n537), .B2(new_n538), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n522), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT85), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n501), .B1(new_n548), .B2(new_n533), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n517), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n464), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n337), .A2(KEYINPUT37), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT38), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n330), .B1(new_n337), .B2(KEYINPUT37), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n334), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n560), .A2(KEYINPUT87), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(KEYINPUT87), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n558), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n562), .B1(new_n565), .B2(KEYINPUT38), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(new_n506), .A3(new_n509), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n551), .A2(new_n556), .A3(new_n557), .A4(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n492), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n569), .A2(KEYINPUT36), .A3(new_n490), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT36), .B1(new_n569), .B2(new_n490), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n572), .B1(new_n427), .B2(new_n464), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n258), .B1(new_n521), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n425), .A2(new_n426), .ZN(new_n576));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n577), .A2(KEYINPUT96), .ZN(new_n578));
  NOR2_X1   g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n577), .A2(KEYINPUT96), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n581), .B1(new_n579), .B2(KEYINPUT95), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n586));
  OAI221_X1 g385(.A(new_n585), .B1(KEYINPUT95), .B2(new_n581), .C1(new_n577), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G127gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n211), .B1(new_n589), .B2(new_n588), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n343), .ZN(new_n598));
  XOR2_X1   g397(.A(G183gat), .B(G211gat), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n600), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT41), .ZN(new_n606));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  OAI22_X1  g406(.A1(new_n605), .A2(KEYINPUT99), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n609));
  INV_X1    g408(.A(G85gat), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT8), .A2(new_n615), .B1(new_n610), .B2(new_n611), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G99gat), .B(G106gat), .Z(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n608), .B1(new_n622), .B2(new_n229), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n228), .A2(new_n231), .A3(new_n621), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n624), .A2(KEYINPUT98), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(KEYINPUT98), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n605), .A2(KEYINPUT99), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT100), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n631), .B(new_n623), .C1(new_n625), .C2(new_n626), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n607), .A2(new_n606), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n630), .A2(new_n636), .A3(new_n632), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n603), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n619), .A2(new_n587), .A3(new_n584), .A4(new_n620), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(KEYINPUT10), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT101), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n621), .A2(new_n588), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n646), .A3(new_n642), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT102), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(new_n642), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G120gat), .B(G148gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n654), .A2(new_n656), .A3(new_n660), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n641), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT103), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n575), .A2(new_n576), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g468(.A1(new_n575), .A2(new_n517), .A3(new_n667), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  AND2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n670), .A2(new_n210), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT42), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(KEYINPUT42), .B2(new_n672), .ZN(G1325gat));
  AND2_X1   g474(.A1(new_n575), .A2(new_n667), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n572), .ZN(new_n678));
  OAI21_X1  g477(.A(G15gat), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n494), .A2(G15gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n677), .B2(new_n680), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n464), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(new_n603), .ZN(new_n687));
  INV_X1    g486(.A(new_n664), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n575), .A2(new_n640), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n215), .A3(new_n576), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT45), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n521), .A2(new_n574), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n640), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT44), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n568), .A2(KEYINPUT106), .A3(new_n573), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT106), .B1(new_n568), .B2(new_n573), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n521), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699));
  INV_X1    g498(.A(new_n640), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n699), .B1(new_n698), .B2(new_n701), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n695), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n576), .ZN(new_n706));
  INV_X1    g505(.A(new_n689), .ZN(new_n707));
  INV_X1    g506(.A(new_n254), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n705), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n692), .B1(new_n711), .B2(new_n215), .ZN(G1328gat));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n705), .A2(new_n518), .A3(new_n710), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n216), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n690), .A2(new_n216), .A3(new_n517), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n713), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n717), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n719), .B(KEYINPUT108), .C1(new_n216), .C2(new_n714), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(G1329gat));
  NAND3_X1  g520(.A1(new_n704), .A2(new_n572), .A3(new_n709), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G43gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n494), .A2(G43gat), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n690), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(KEYINPUT47), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n722), .A2(new_n728), .A3(G43gat), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n722), .B2(G43gat), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n729), .A2(new_n730), .A3(new_n725), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(G1330gat));
  NAND2_X1  g532(.A1(new_n464), .A2(new_n430), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT111), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n690), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n705), .A2(new_n557), .A3(new_n710), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(new_n430), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT48), .B(new_n736), .C1(new_n737), .C2(new_n430), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1331gat));
  NAND4_X1  g541(.A1(new_n698), .A2(new_n708), .A3(new_n641), .A4(new_n688), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n576), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n518), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n743), .B2(new_n678), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n493), .A2(new_n481), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n743), .B2(new_n753), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g554(.A1(new_n744), .A2(new_n464), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g556(.A1(new_n687), .A2(new_n254), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n688), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT112), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n705), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n706), .ZN(new_n762));
  INV_X1    g561(.A(new_n698), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n758), .A2(new_n640), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n576), .A2(new_n610), .A3(new_n688), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n762), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n705), .A2(new_n518), .A3(new_n760), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n611), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n517), .A2(new_n611), .A3(new_n688), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT52), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  OAI221_X1 g575(.A(new_n776), .B1(new_n768), .B2(new_n773), .C1(new_n771), .C2(new_n611), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n761), .B2(new_n678), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n688), .A2(new_n483), .A3(new_n493), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n768), .B2(new_n780), .ZN(G1338gat));
  NOR2_X1   g580(.A1(new_n664), .A2(G106gat), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n464), .B(new_n782), .C1(new_n766), .C2(new_n767), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n705), .A2(new_n557), .A3(new_n760), .ZN(new_n784));
  INV_X1    g583(.A(G106gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  OAI221_X1 g589(.A(new_n783), .B1(new_n788), .B2(new_n787), .C1(new_n784), .C2(new_n785), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1339gat));
  NAND4_X1  g591(.A1(new_n645), .A2(new_n649), .A3(new_n652), .A4(new_n647), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n650), .A2(new_n795), .A3(new_n653), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n794), .A2(KEYINPUT55), .A3(new_n661), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n663), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n663), .A3(KEYINPUT114), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  INV_X1    g601(.A(new_n794), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n796), .A2(new_n661), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n800), .A2(new_n254), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n249), .A2(new_n244), .A3(new_n250), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n247), .A2(new_n248), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n233), .B1(new_n232), .B2(new_n235), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n243), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n688), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n640), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n800), .A2(new_n801), .A3(new_n805), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n640), .A2(new_n811), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n603), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n641), .A2(new_n708), .A3(new_n664), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n500), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n706), .A2(new_n517), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n821), .A2(new_n368), .A3(new_n258), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n818), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n820), .ZN(new_n824));
  INV_X1    g623(.A(new_n495), .ZN(new_n825));
  INV_X1    g624(.A(new_n496), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n254), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n822), .B1(new_n831), .B2(new_n368), .ZN(G1340gat));
  NOR3_X1   g631(.A1(new_n821), .A2(new_n369), .A3(new_n664), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n688), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(new_n369), .ZN(G1341gat));
  OAI21_X1  g634(.A(G127gat), .B1(new_n821), .B2(new_n603), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n687), .A2(new_n593), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n829), .B2(new_n837), .ZN(G1342gat));
  NOR3_X1   g637(.A1(new_n829), .A2(G134gat), .A3(new_n700), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n821), .B2(new_n700), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n557), .A2(new_n572), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n824), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n258), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n351), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(KEYINPUT58), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n823), .A2(new_n464), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  INV_X1    g653(.A(new_n804), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT55), .B1(new_n855), .B2(new_n794), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n854), .B1(new_n798), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n805), .A2(KEYINPUT115), .A3(new_n663), .A4(new_n797), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n256), .A2(new_n857), .A3(new_n257), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n640), .B1(new_n859), .B2(new_n812), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n603), .B1(new_n860), .B2(new_n816), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n818), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n557), .A2(new_n852), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n853), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n862), .B2(new_n864), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n706), .A2(new_n517), .A3(new_n572), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n254), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n351), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n850), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G141gat), .B1(new_n870), .B2(new_n258), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n849), .B2(new_n848), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n873), .B2(new_n877), .ZN(G1344gat));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n861), .B1(new_n666), .B2(new_n847), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n852), .A3(new_n464), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n881), .A2(new_n688), .A3(new_n869), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n879), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n688), .B(new_n869), .C1(new_n866), .C2(new_n867), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n347), .A2(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n885), .A2(KEYINPUT118), .A3(new_n886), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n846), .A2(new_n347), .A3(new_n688), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n885), .A2(KEYINPUT118), .A3(new_n886), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT118), .B1(new_n885), .B2(new_n886), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n895), .B(new_n892), .C1(new_n898), .C2(new_n884), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n894), .A2(new_n899), .ZN(G1345gat));
  AOI21_X1  g699(.A(G155gat), .B1(new_n846), .B2(new_n687), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n687), .A2(G155gat), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT120), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n871), .B2(new_n903), .ZN(G1346gat));
  NAND3_X1  g703(.A1(new_n846), .A2(new_n344), .A3(new_n640), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n870), .B2(new_n700), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G162gat), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n870), .A2(new_n906), .A3(new_n700), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n576), .A2(new_n518), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n819), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n275), .A3(new_n258), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n576), .B1(new_n817), .B2(new_n818), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n517), .A3(new_n828), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT122), .Z(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n254), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n913), .B1(new_n917), .B2(new_n275), .ZN(G1348gat));
  NOR3_X1   g717(.A1(new_n912), .A2(new_n276), .A3(new_n664), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n688), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n276), .ZN(G1349gat));
  OAI21_X1  g721(.A(G183gat), .B1(new_n912), .B2(new_n603), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n687), .A2(new_n281), .A3(new_n283), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n915), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n926));
  NAND2_X1  g725(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n916), .A2(new_n284), .A3(new_n640), .ZN(new_n929));
  OAI21_X1  g728(.A(G190gat), .B1(new_n912), .B2(new_n700), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(KEYINPUT125), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(KEYINPUT61), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n929), .B(new_n933), .C1(KEYINPUT61), .C2(new_n932), .ZN(G1351gat));
  NAND2_X1  g733(.A1(new_n845), .A2(new_n517), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT126), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n936), .A2(new_n914), .ZN(new_n937));
  AOI21_X1  g736(.A(G197gat), .B1(new_n937), .B2(new_n254), .ZN(new_n938));
  AND4_X1   g737(.A1(new_n678), .A2(new_n881), .A3(new_n882), .A4(new_n911), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n847), .A2(G197gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(G1352gat));
  INV_X1    g740(.A(G204gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n937), .A2(new_n942), .A3(new_n688), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT62), .Z(new_n944));
  AND2_X1   g743(.A1(new_n939), .A2(new_n688), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n942), .ZN(G1353gat));
  NAND3_X1  g745(.A1(new_n937), .A2(new_n263), .A3(new_n687), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n939), .A2(new_n687), .ZN(new_n948));
  AND4_X1   g747(.A1(KEYINPUT127), .A2(new_n948), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n948), .A2(new_n951), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n947), .B1(new_n949), .B2(new_n952), .ZN(G1354gat));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n264), .A3(new_n640), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n939), .A2(new_n640), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n264), .ZN(G1355gat));
endmodule


