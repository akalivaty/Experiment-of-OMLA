//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1205, new_n1206, new_n1207,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT65), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  NAND3_X1  g0006(.A1(new_n201), .A2(KEYINPUT65), .A3(new_n202), .ZN(new_n207));
  AND3_X1   g0007(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(G353));
  NOR2_X1   g0008(.A1(G97), .A2(G107), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G87), .ZN(G355));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n213), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  INV_X1    g0029(.A(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G107), .ZN(new_n231));
  INV_X1    g0031(.A(G264), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n229), .B1(new_n206), .B2(new_n230), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n215), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n218), .B1(new_n221), .B2(new_n222), .C1(KEYINPUT1), .C2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(KEYINPUT1), .B2(new_n234), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n252), .A2(new_n213), .A3(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n219), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n212), .A2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G77), .A3(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n252), .A2(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(G77), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n263), .A2(new_n264), .B1(G20), .B2(G77), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n213), .A2(G33), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT15), .B(G87), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n261), .B1(new_n268), .B2(new_n255), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n276), .A2(G238), .B1(G107), .B2(new_n274), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1698), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G232), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n271), .B1(new_n284), .B2(KEYINPUT67), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT67), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n277), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(new_n271), .A3(G274), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n271), .A2(new_n289), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n291), .B1(new_n230), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n269), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n293), .B1(new_n285), .B2(new_n287), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n298), .A2(KEYINPUT68), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT68), .B1(new_n298), .B2(new_n299), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n298), .A2(G190), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n303), .B(new_n269), .C1(new_n304), .C2(new_n298), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT69), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n213), .B1(new_n205), .B2(new_n207), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n264), .A2(G150), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n262), .B2(new_n266), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n255), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G50), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n212), .B2(G20), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n256), .A2(new_n313), .B1(new_n312), .B2(new_n253), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G226), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n291), .B1(new_n316), .B2(new_n292), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n276), .A2(G223), .B1(G77), .B2(new_n274), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n282), .A2(G222), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n271), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n299), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n315), .B(new_n323), .C1(G169), .C2(new_n322), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(G190), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n304), .B2(new_n322), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT9), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(new_n315), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n311), .A2(KEYINPUT9), .A3(new_n314), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT70), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(KEYINPUT10), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n324), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G232), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n291), .B1(new_n335), .B2(new_n292), .ZN(new_n336));
  INV_X1    g0136(.A(G223), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(G1698), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n272), .B2(new_n273), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT75), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n280), .A2(new_n281), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT75), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(new_n338), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(G226), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT74), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n345), .A2(new_n346), .B1(G33), .B2(G87), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n341), .A2(KEYINPUT74), .A3(G226), .A4(G1698), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n336), .B1(new_n349), .B2(new_n321), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n296), .ZN(new_n351));
  AOI211_X1 g0151(.A(new_n299), .B(new_n336), .C1(new_n349), .C2(new_n321), .ZN(new_n352));
  INV_X1    g0152(.A(G58), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(new_n224), .ZN(new_n354));
  OAI21_X1  g0154(.A(G20), .B1(new_n354), .B2(new_n202), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n264), .A2(G159), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(KEYINPUT16), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n274), .B2(new_n213), .ZN(new_n359));
  NOR4_X1   g0159(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT7), .A4(G20), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT73), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n274), .A2(new_n213), .ZN(new_n362));
  NOR2_X1   g0162(.A1(KEYINPUT73), .A2(KEYINPUT7), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n224), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n357), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT7), .B1(new_n341), .B2(G20), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n274), .A2(new_n358), .A3(new_n213), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(G68), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n355), .A2(new_n356), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT16), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n255), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n365), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n262), .B1(new_n212), .B2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n256), .B1(new_n262), .B2(new_n253), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n351), .A2(new_n352), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n349), .A2(new_n321), .ZN(new_n379));
  INV_X1    g0179(.A(new_n336), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(G179), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n296), .B2(new_n350), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n368), .A2(new_n369), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n357), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n366), .B2(new_n367), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n362), .A2(new_n363), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G68), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n386), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n385), .A2(new_n391), .A3(new_n255), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n374), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n382), .A2(new_n393), .A3(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT76), .ZN(new_n396));
  AOI21_X1  g0196(.A(G200), .B1(new_n379), .B2(new_n380), .ZN(new_n397));
  AOI211_X1 g0197(.A(G190), .B(new_n336), .C1(new_n349), .C2(new_n321), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n396), .B1(new_n399), .B2(new_n393), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n379), .A2(new_n401), .A3(new_n380), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(G200), .B2(new_n350), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n361), .A2(new_n364), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n371), .B1(new_n404), .B2(new_n386), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n375), .B1(new_n405), .B2(new_n385), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n378), .A2(new_n394), .B1(new_n400), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n256), .A2(G68), .A3(new_n257), .ZN(new_n411));
  XOR2_X1   g0211(.A(new_n411), .B(KEYINPUT72), .Z(new_n412));
  AOI22_X1  g0212(.A1(new_n264), .A2(G50), .B1(G20), .B2(new_n224), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n206), .B2(new_n266), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n414), .A2(new_n255), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n253), .A2(new_n224), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT12), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n412), .A2(new_n416), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n291), .B1(new_n225), .B2(new_n292), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G97), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n335), .A2(G1698), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(G226), .B2(G1698), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n424), .B1(new_n426), .B2(new_n274), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n321), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n422), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n423), .B1(new_n422), .B2(new_n428), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G169), .B1(new_n429), .B2(new_n430), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n431), .A2(new_n299), .B1(new_n432), .B2(KEYINPUT14), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n420), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n431), .A2(new_n401), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n420), .ZN(new_n437));
  OAI21_X1  g0237(.A(G200), .B1(new_n429), .B2(new_n430), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT71), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n410), .A2(new_n435), .A3(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n307), .A2(new_n334), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G41), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n212), .B(G45), .C1(new_n444), .C2(KEYINPUT5), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT5), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G41), .ZN(new_n447));
  OAI211_X1 g0247(.A(G257), .B(new_n271), .C1(new_n445), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n282), .A2(G244), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n276), .A2(G250), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n452), .A2(new_n453), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n449), .B1(new_n456), .B2(new_n321), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT79), .B1(new_n446), .B2(G41), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(new_n444), .A3(KEYINPUT5), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n446), .A2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n458), .A2(new_n460), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n271), .A2(G274), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n457), .A2(G179), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n466), .ZN(new_n468));
  AOI211_X1 g0268(.A(new_n449), .B(new_n468), .C1(new_n456), .C2(new_n321), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n469), .B2(new_n296), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n366), .A2(G107), .A3(new_n367), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT77), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n231), .A2(KEYINPUT6), .A3(G97), .ZN(new_n474));
  INV_X1    g0274(.A(G97), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n231), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n209), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n477), .B2(KEYINPUT6), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n264), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n471), .A2(new_n472), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n255), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n260), .A2(G97), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n212), .A2(G33), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n371), .A2(new_n260), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n483), .B1(new_n486), .B2(G97), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n470), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(KEYINPUT78), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT78), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n482), .A2(new_n491), .A3(new_n487), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n457), .A2(new_n466), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n304), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n469), .A2(new_n401), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n489), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G116), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT80), .B1(new_n485), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT80), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n256), .A2(new_n501), .A3(G116), .A4(new_n484), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n455), .B(new_n213), .C1(G33), .C2(new_n475), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(G20), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n255), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n504), .A2(KEYINPUT20), .A3(new_n255), .A4(new_n505), .ZN(new_n509));
  INV_X1    g0309(.A(new_n505), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n508), .A2(new_n509), .B1(new_n259), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n503), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n341), .A2(G264), .A3(G1698), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n341), .A2(G257), .A3(new_n275), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n274), .A2(G303), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n321), .ZN(new_n517));
  OAI211_X1 g0317(.A(G270), .B(new_n271), .C1(new_n445), .C2(new_n447), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n466), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n512), .A2(new_n519), .A3(G169), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(G200), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n466), .A2(new_n518), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G190), .A3(new_n517), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n523), .A2(new_n526), .A3(new_n503), .A4(new_n511), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n512), .A2(G179), .A3(new_n517), .A4(new_n525), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n512), .A2(new_n519), .A3(KEYINPUT21), .A4(G169), .ZN(new_n529));
  AND4_X1   g0329(.A1(new_n522), .A2(new_n527), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT25), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n260), .B2(G107), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n231), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n486), .A2(G107), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT82), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT81), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n213), .A3(G87), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n274), .B2(new_n538), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n226), .A2(KEYINPUT81), .A3(G20), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n341), .A2(KEYINPUT22), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(G20), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n213), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n231), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n539), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT24), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n539), .A2(new_n541), .A3(new_n547), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n535), .B1(new_n552), .B2(new_n255), .ZN(new_n553));
  AOI211_X1 g0353(.A(KEYINPUT82), .B(new_n371), .C1(new_n549), .C2(new_n551), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n534), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n271), .B1(new_n445), .B2(new_n447), .ZN(new_n556));
  OAI22_X1  g0356(.A1(new_n556), .A2(new_n232), .B1(new_n464), .B2(new_n465), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G257), .B(G1698), .C1(new_n272), .C2(new_n273), .ZN(new_n559));
  OAI211_X1 g0359(.A(G250), .B(new_n275), .C1(new_n272), .C2(new_n273), .ZN(new_n560));
  INV_X1    g0360(.A(G294), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n559), .B(new_n560), .C1(new_n279), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n321), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n296), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n555), .B(new_n565), .C1(G179), .C2(new_n564), .ZN(new_n566));
  OR3_X1    g0366(.A1(new_n462), .A2(G1), .A3(G274), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n227), .B1(new_n462), .B2(G1), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n271), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n282), .A2(G238), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n341), .A2(G244), .A3(G1698), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n572), .A3(new_n542), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n570), .B1(new_n573), .B2(new_n321), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G200), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(G190), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n341), .A2(new_n213), .A3(G68), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n213), .B1(new_n424), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(G87), .B2(new_n210), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n266), .B2(new_n475), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(new_n255), .B1(new_n267), .B2(new_n253), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n486), .A2(G87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n267), .B2(new_n485), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n574), .A2(new_n299), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n574), .A2(G169), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n578), .A2(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n282), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n271), .B1(new_n594), .B2(new_n559), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n595), .A2(new_n401), .A3(new_n557), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n304), .B1(new_n558), .B2(new_n563), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n598), .B(new_n534), .C1(new_n553), .C2(new_n554), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n530), .A2(new_n566), .A3(new_n593), .A4(new_n599), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n443), .A2(new_n498), .A3(new_n600), .ZN(G372));
  OAI211_X1 g0401(.A(new_n440), .B(new_n297), .C1(new_n301), .C2(new_n300), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(new_n435), .B1(new_n409), .B2(new_n400), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT84), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n382), .A2(new_n393), .A3(KEYINPUT18), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT18), .B1(new_n382), .B2(new_n393), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n378), .A2(KEYINPUT84), .A3(new_n394), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n603), .A2(new_n609), .B1(new_n332), .B2(new_n333), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n324), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n590), .A2(new_n591), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n585), .A2(new_n614), .A3(new_n586), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n585), .B2(new_n586), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n576), .B(new_n577), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n599), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n522), .A2(new_n528), .A3(new_n529), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n566), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n494), .A2(G169), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(new_n467), .B1(new_n482), .B2(new_n487), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n482), .A2(new_n491), .A3(new_n487), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n491), .B1(new_n482), .B2(new_n487), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n496), .B1(G200), .B2(new_n469), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n613), .B1(new_n621), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n593), .A2(new_n623), .A3(KEYINPUT26), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n470), .B1(new_n624), .B2(new_n625), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n618), .B1(new_n591), .B2(new_n590), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n630), .B1(new_n633), .B2(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n612), .B1(new_n443), .B2(new_n636), .ZN(G369));
  NAND2_X1  g0437(.A1(new_n259), .A2(new_n213), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n512), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT85), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n522), .A2(new_n528), .A3(new_n529), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n620), .A2(new_n527), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n645), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n649), .A2(KEYINPUT86), .A3(G330), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT86), .B1(new_n649), .B2(G330), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n566), .A2(new_n599), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n555), .A2(new_n643), .ZN(new_n656));
  INV_X1    g0456(.A(new_n643), .ZN(new_n657));
  OAI22_X1  g0457(.A1(new_n655), .A2(new_n656), .B1(new_n566), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n566), .A2(new_n643), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n646), .A2(new_n657), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n659), .A2(new_n660), .A3(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n216), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n210), .A2(G87), .A3(G116), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G1), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n222), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n635), .A2(new_n657), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(KEYINPUT29), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n489), .A2(new_n592), .A3(KEYINPUT26), .ZN(new_n674));
  INV_X1    g0474(.A(new_n578), .ZN(new_n675));
  INV_X1    g0475(.A(new_n617), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n615), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n613), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(new_n493), .A3(new_n470), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n674), .B1(KEYINPUT26), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n643), .B1(new_n629), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT87), .B1(new_n519), .B2(new_n299), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n575), .A2(new_n564), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT87), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n525), .A2(new_n687), .A3(G179), .A4(new_n517), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n685), .A2(new_n686), .A3(new_n688), .A4(new_n457), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n564), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n457), .A2(new_n692), .A3(new_n574), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT30), .A3(new_n688), .A4(new_n685), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n692), .A2(new_n574), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(new_n494), .A3(new_n299), .A4(new_n519), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n691), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n643), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n600), .A2(new_n498), .A3(new_n643), .ZN(new_n703));
  OAI21_X1  g0503(.A(G330), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n684), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n671), .B1(new_n706), .B2(G1), .ZN(G364));
  NOR2_X1   g0507(.A1(new_n649), .A2(G330), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT88), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n252), .A2(G20), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n212), .B1(new_n710), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n666), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(new_n652), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT89), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n216), .A2(new_n341), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(KEYINPUT90), .B2(G355), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(KEYINPUT90), .B2(G355), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(G116), .B2(new_n216), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n247), .A2(G45), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n665), .A2(new_n341), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n222), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n462), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n720), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(G13), .A2(G33), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n219), .B1(G20), .B2(new_n296), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n713), .B1(new_n726), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n213), .A2(new_n401), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n299), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n213), .A2(G190), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n735), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(G58), .A2(new_n737), .B1(new_n740), .B2(G77), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n741), .A2(KEYINPUT91), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n738), .A2(new_n299), .A3(G200), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n734), .A2(new_n299), .A3(G200), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n341), .B1(new_n743), .B2(new_n231), .C1(new_n226), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(KEYINPUT91), .B2(new_n741), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT32), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n738), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n748), .B1(new_n751), .B2(G159), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n213), .B1(new_n749), .B2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n475), .ZN(new_n754));
  INV_X1    g0554(.A(G159), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n750), .A2(KEYINPUT32), .A3(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT92), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n401), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n759), .A2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n757), .B1(new_n312), .B2(new_n761), .C1(new_n224), .C2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n743), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n765), .A2(G283), .B1(new_n751), .B2(G329), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT93), .ZN(new_n767));
  INV_X1    g0567(.A(G303), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n744), .A2(new_n768), .B1(new_n736), .B2(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n341), .B(new_n770), .C1(G311), .C2(new_n740), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n767), .B(new_n771), .C1(new_n561), .C2(new_n753), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n760), .A2(G326), .ZN(new_n773));
  XOR2_X1   g0573(.A(KEYINPUT33), .B(G317), .Z(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n763), .B2(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n747), .A2(new_n764), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n733), .B1(new_n776), .B2(new_n730), .ZN(new_n777));
  INV_X1    g0577(.A(new_n729), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n649), .B2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT94), .Z(new_n780));
  NAND2_X1  g0580(.A1(new_n716), .A2(new_n780), .ZN(G396));
  NOR2_X1   g0581(.A1(new_n269), .A2(new_n657), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n302), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n302), .A2(new_n305), .A3(new_n783), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT97), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n672), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT98), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT98), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n643), .B1(new_n629), .B2(new_n634), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n786), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n713), .B1(new_n793), .B2(new_n704), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n704), .B2(new_n793), .ZN(new_n795));
  INV_X1    g0595(.A(new_n730), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n728), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n713), .B1(G77), .B2(new_n797), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n744), .A2(new_n231), .B1(new_n743), .B2(new_n226), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n739), .A2(new_n499), .B1(new_n750), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n274), .B1(new_n736), .B2(new_n561), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n799), .A2(new_n801), .A3(new_n802), .A4(new_n754), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n804), .B2(new_n763), .C1(new_n768), .C2(new_n761), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT95), .B(G143), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n737), .A2(new_n806), .B1(new_n740), .B2(G159), .ZN(new_n807));
  INV_X1    g0607(.A(G150), .ZN(new_n808));
  INV_X1    g0608(.A(G137), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n763), .B2(new_n808), .C1(new_n809), .C2(new_n761), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n744), .A2(new_n312), .B1(new_n750), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n743), .A2(new_n224), .ZN(new_n815));
  NOR3_X1   g0615(.A1(new_n814), .A2(new_n274), .A3(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n812), .B(new_n816), .C1(new_n353), .C2(new_n753), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n810), .A2(new_n811), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n805), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT96), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n796), .B1(new_n819), .B2(new_n820), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n798), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n786), .B2(new_n728), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n795), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  AND2_X1   g0626(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n827), .A2(new_n828), .A3(new_n221), .A4(new_n499), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT36), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n201), .A2(G68), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n724), .B(G77), .C1(new_n353), .C2(new_n224), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n212), .B(G13), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n710), .A2(new_n212), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT40), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n378), .A2(new_n394), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n400), .A2(new_n409), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n391), .A2(new_n255), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT16), .B1(new_n404), .B2(new_n369), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n374), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n641), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n392), .B(new_n374), .C1(new_n397), .C2(new_n398), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT37), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n843), .B1(new_n372), .B2(new_n375), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n376), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n381), .B(new_n641), .C1(new_n296), .C2(new_n350), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n851), .A2(new_n842), .B1(new_n403), .B2(new_n406), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT38), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n853), .B(KEYINPUT38), .C1(new_n410), .C2(new_n844), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT102), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n702), .B2(new_n703), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n648), .A2(new_n592), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n861), .A2(new_n628), .A3(new_n654), .A4(new_n657), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n862), .A2(KEYINPUT102), .A3(new_n700), .A4(new_n701), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n440), .A2(new_n435), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(new_n420), .A3(new_n643), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n420), .A2(new_n643), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n440), .A2(new_n435), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n860), .A2(new_n786), .A3(new_n863), .A4(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n836), .B1(new_n858), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n855), .A2(KEYINPUT99), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT99), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n846), .A2(new_n872), .A3(KEYINPUT38), .A4(new_n853), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n607), .A2(new_n608), .A3(new_n838), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n641), .B1(new_n392), .B2(new_n374), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n847), .A2(new_n849), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n350), .A2(new_n296), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n406), .B1(new_n879), .B2(new_n381), .ZN(new_n880));
  NOR4_X1   g0680(.A1(new_n878), .A2(new_n880), .A3(new_n604), .A4(new_n848), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n876), .B1(new_n406), .B2(new_n403), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n847), .A2(new_n604), .A3(new_n849), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n376), .A2(new_n882), .B1(new_n883), .B2(KEYINPUT37), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n874), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT40), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n870), .B(G330), .C1(new_n869), .C2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n860), .A2(G330), .A3(new_n863), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n443), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT103), .Z(new_n896));
  OR2_X1    g0696(.A1(new_n890), .A2(new_n869), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n870), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n442), .A2(new_n860), .A3(new_n863), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n435), .A2(new_n643), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT100), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n874), .A2(new_n902), .A3(new_n903), .A4(new_n888), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n871), .A2(new_n873), .A3(new_n903), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n877), .B2(new_n885), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT100), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n901), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n302), .A2(new_n643), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n791), .B2(new_n786), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n857), .A3(new_n868), .ZN(new_n915));
  INV_X1    g0715(.A(new_n609), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n915), .B1(new_n916), .B2(new_n843), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n442), .B1(new_n673), .B2(new_n683), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT101), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT101), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n922), .B(new_n442), .C1(new_n673), .C2(new_n683), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n612), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n918), .B(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n835), .B1(new_n900), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT104), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n927), .A2(new_n928), .B1(new_n926), .B2(new_n900), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n834), .B1(new_n929), .B2(new_n930), .ZN(G367));
  NOR2_X1   g0731(.A1(new_n677), .A2(new_n657), .ZN(new_n932));
  MUX2_X1   g0732(.A(new_n678), .B(new_n613), .S(new_n932), .Z(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n628), .B1(new_n626), .B2(new_n657), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n493), .A2(new_n470), .A3(new_n643), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(new_n663), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT42), .Z(new_n939));
  OAI21_X1  g0739(.A(new_n489), .B1(new_n937), .B2(new_n566), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n940), .A2(new_n657), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n934), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT43), .B1(new_n933), .B2(KEYINPUT105), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(KEYINPUT105), .B2(new_n933), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT106), .Z(new_n945));
  AND2_X1   g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n942), .A2(new_n945), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n659), .A2(new_n937), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n666), .B(KEYINPUT41), .Z(new_n951));
  INV_X1    g0751(.A(new_n659), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n663), .A2(new_n660), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n937), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n937), .A2(new_n954), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT44), .Z(new_n958));
  NAND3_X1  g0758(.A1(new_n953), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n663), .B1(new_n658), .B2(new_n662), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(new_n652), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n705), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n951), .B1(new_n966), .B2(new_n706), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n950), .B1(new_n967), .B2(new_n712), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n731), .B1(new_n216), .B2(new_n267), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n722), .B2(new_n243), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n714), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n744), .A2(new_n499), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(KEYINPUT46), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n341), .B(new_n973), .C1(G283), .C2(new_n740), .ZN(new_n974));
  INV_X1    g0774(.A(G317), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n743), .A2(new_n475), .B1(new_n750), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G303), .B2(new_n737), .ZN(new_n977));
  INV_X1    g0777(.A(new_n753), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n972), .A2(KEYINPUT46), .B1(G107), .B2(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G294), .A2(new_n762), .B1(new_n760), .B2(G311), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n974), .A2(new_n977), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n744), .A2(new_n353), .B1(new_n750), .B2(new_n809), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n341), .B1(new_n753), .B2(new_n224), .C1(new_n808), .C2(new_n736), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(G77), .C2(new_n765), .ZN(new_n984));
  INV_X1    g0784(.A(new_n201), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n762), .A2(G159), .B1(new_n985), .B2(new_n740), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n760), .A2(new_n806), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n981), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT47), .Z(new_n992));
  OAI221_X1 g0792(.A(new_n971), .B1(new_n778), .B2(new_n933), .C1(new_n992), .C2(new_n796), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n968), .A2(new_n993), .ZN(G387));
  INV_X1    g0794(.A(new_n965), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n705), .A2(new_n964), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n995), .A2(new_n666), .A3(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n668), .B(new_n462), .C1(new_n224), .C2(new_n206), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT109), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(KEYINPUT50), .B1(new_n262), .B2(G50), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n262), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n998), .A2(new_n999), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n722), .B1(new_n1003), .B2(new_n1004), .C1(new_n240), .C2(new_n462), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(G107), .B2(new_n216), .C1(new_n668), .C2(new_n717), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n714), .B1(new_n1006), .B2(new_n731), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G317), .A2(new_n737), .B1(new_n740), .B2(G303), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n763), .B2(new_n800), .C1(new_n769), .C2(new_n761), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT48), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n744), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1013), .A2(G294), .B1(new_n978), .B2(G283), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT110), .Z(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n743), .A2(new_n499), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n341), .B(new_n1019), .C1(G326), .C2(new_n751), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n744), .A2(new_n206), .B1(new_n739), .B2(new_n224), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n736), .A2(new_n312), .B1(new_n750), .B2(new_n808), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n341), .B1(new_n743), .B2(new_n475), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n753), .A2(new_n267), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n755), .B2(new_n761), .C1(new_n262), .C2(new_n763), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1007), .B1(new_n658), .B2(new_n778), .C1(new_n1028), .C2(new_n796), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n997), .B(new_n1029), .C1(new_n711), .C2(new_n964), .ZN(G393));
  INV_X1    g0830(.A(new_n962), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n995), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n667), .B1(new_n962), .B2(new_n965), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n937), .A2(new_n729), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G294), .A2(new_n740), .B1(new_n978), .B2(G116), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n763), .B2(new_n768), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT112), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n760), .A2(G317), .B1(G311), .B2(new_n737), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT52), .Z(new_n1040));
  OAI22_X1  g0840(.A1(new_n744), .A2(new_n804), .B1(new_n750), .B2(new_n769), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n341), .B(new_n1041), .C1(G107), .C2(new_n765), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n760), .A2(G150), .B1(G159), .B2(new_n737), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT51), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1013), .A2(G68), .B1(new_n751), .B2(new_n806), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT111), .Z(new_n1047));
  NOR2_X1   g0847(.A1(new_n753), .A2(new_n206), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n341), .B1(new_n743), .B2(new_n226), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n263), .C2(new_n740), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1047), .B(new_n1050), .C1(new_n201), .C2(new_n763), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1043), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n730), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n731), .B1(new_n475), .B2(new_n216), .C1(new_n723), .C2(new_n250), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1035), .A2(new_n713), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1034), .B(new_n1055), .C1(new_n711), .C2(new_n1031), .ZN(G390));
  INV_X1    g0856(.A(KEYINPUT115), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n868), .A2(new_n786), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n892), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n868), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n901), .B1(new_n913), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1061), .A2(new_n904), .A3(new_n909), .A4(new_n905), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n912), .B1(new_n681), .B2(new_n786), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n889), .B(new_n901), .C1(new_n1060), .C2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g0864(.A(KEYINPUT113), .B(new_n1059), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT113), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1059), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n704), .B1(new_n785), .B2(new_n784), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n868), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1062), .A2(new_n1064), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1065), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n611), .B(new_n893), .C1(new_n920), .C2(new_n923), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1070), .A2(new_n868), .B1(new_n892), .B2(new_n1058), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n914), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT114), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n787), .B1(new_n892), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n860), .A2(KEYINPUT114), .A3(new_n863), .A4(G330), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n868), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1071), .A2(new_n1063), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1076), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1074), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1057), .B1(new_n1073), .B2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1074), .A2(new_n1082), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1072), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1059), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n1066), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1085), .B(KEYINPUT115), .C1(new_n1088), .C2(new_n1065), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n667), .B1(new_n1073), .B2(new_n1083), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1073), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n906), .A2(new_n727), .A3(new_n909), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n713), .B1(new_n263), .B2(new_n797), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n743), .A2(new_n224), .B1(new_n739), .B2(new_n475), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n274), .B1(new_n744), .B2(new_n226), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n736), .A2(new_n499), .B1(new_n750), .B2(new_n561), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1048), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n231), .B2(new_n763), .C1(new_n804), .C2(new_n761), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n744), .A2(new_n808), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1102));
  OAI22_X1  g0902(.A1(new_n1101), .A2(new_n1102), .B1(new_n755), .B2(new_n753), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1104));
  INV_X1    g0904(.A(G125), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n201), .A2(new_n743), .B1(new_n750), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n274), .B(new_n1106), .C1(G132), .C2(new_n737), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT54), .B(G143), .Z(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT116), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n740), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1104), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(G128), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1112), .A2(new_n761), .B1(new_n763), .B2(new_n809), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1100), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1095), .B1(new_n1114), .B2(new_n730), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1093), .A2(new_n712), .B1(new_n1094), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1092), .A2(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(KEYINPUT57), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1074), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n334), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n315), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n641), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n334), .A2(new_n315), .A3(new_n843), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n891), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n897), .A2(new_n1128), .A3(G330), .A4(new_n870), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n918), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1130), .B(new_n1131), .C1(new_n910), .C2(new_n917), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(KEYINPUT119), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT119), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1136), .A3(new_n918), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1118), .B1(new_n1120), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT120), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(KEYINPUT120), .B(new_n1118), .C1(new_n1120), .C2(new_n1138), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1120), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(new_n1118), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n667), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1141), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1135), .A2(new_n712), .A3(new_n1137), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n713), .B1(new_n985), .B2(new_n797), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n279), .B(new_n444), .C1(new_n743), .C2(new_n755), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n753), .A2(new_n808), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n736), .A2(new_n1112), .B1(new_n739), .B2(new_n809), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(new_n1109), .C2(new_n1013), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n1105), .B2(new_n761), .C1(new_n813), .C2(new_n763), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1154), .A2(KEYINPUT59), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1150), .B(new_n1155), .C1(G124), .C2(new_n751), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(KEYINPUT59), .B2(new_n1154), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n341), .A2(G41), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G50), .B(new_n1158), .C1(new_n279), .C2(new_n444), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT118), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G107), .A2(new_n737), .B1(new_n751), .B2(G283), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n353), .B2(new_n743), .C1(new_n267), .C2(new_n739), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n761), .A2(new_n499), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n763), .A2(new_n475), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1158), .B1(new_n224), .B2(new_n753), .C1(new_n206), .C2(new_n744), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1160), .B1(new_n1166), .B2(KEYINPUT58), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1157), .B(new_n1167), .C1(KEYINPUT58), .C2(new_n1166), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1149), .B1(new_n1168), .B2(new_n730), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1129), .B2(new_n728), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1148), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1147), .A2(new_n1171), .ZN(G375));
  NAND3_X1  g0972(.A1(new_n1082), .A2(KEYINPUT121), .A3(new_n712), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n713), .B1(G68), .B2(new_n797), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n868), .A2(new_n728), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n744), .A2(new_n475), .B1(new_n736), .B2(new_n804), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n739), .A2(new_n231), .B1(new_n750), .B2(new_n768), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n274), .B1(new_n743), .B2(new_n206), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .A4(new_n1025), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n499), .B2(new_n763), .C1(new_n561), .C2(new_n761), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1109), .A2(new_n762), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n760), .A2(G132), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n744), .A2(new_n755), .B1(new_n739), .B2(new_n808), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n736), .A2(new_n809), .B1(new_n750), .B2(new_n1112), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n341), .B1(new_n743), .B2(new_n353), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G50), .B2(new_n978), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1182), .A2(new_n1183), .A3(new_n1186), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1181), .A2(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1190), .A2(KEYINPUT122), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n796), .B1(new_n1190), .B2(KEYINPUT122), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1175), .B(new_n1176), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT121), .B1(new_n1082), .B2(new_n712), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1174), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1074), .A2(new_n1082), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n951), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(new_n1197), .A3(new_n1083), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1195), .A2(new_n1198), .ZN(G381));
  OR2_X1    g0999(.A1(G393), .A2(G396), .ZN(new_n1200));
  OR4_X1    g1000(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(G378), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1147), .A2(new_n1202), .A3(new_n1171), .ZN(new_n1203));
  OR3_X1    g1003(.A1(new_n1201), .A2(new_n1203), .A3(G381), .ZN(G407));
  NAND2_X1  g1004(.A1(new_n642), .A2(G213), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT123), .Z(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G407), .B(G213), .C1(new_n1203), .C2(new_n1207), .ZN(G409));
  NAND2_X1  g1008(.A1(new_n1083), .A2(KEYINPUT60), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n666), .B1(new_n1209), .B2(new_n1196), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1196), .B2(new_n1209), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1195), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(new_n825), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1147), .A2(G378), .A3(new_n1171), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1170), .B1(new_n1144), .B2(new_n711), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1120), .A2(new_n1138), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1217), .B2(new_n1197), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT124), .B1(new_n1218), .B2(G378), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT124), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1120), .A2(new_n951), .A3(new_n1138), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1202), .B(new_n1220), .C1(new_n1221), .C2(new_n1216), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1207), .B(new_n1214), .C1(new_n1215), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT62), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1207), .B1(new_n1215), .B2(new_n1223), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1213), .B(G384), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1206), .A2(G2897), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1227), .B(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT61), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1147), .A2(G378), .A3(new_n1171), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(new_n1219), .A3(new_n1222), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT62), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1207), .A4(new_n1214), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1225), .A2(new_n1230), .A3(new_n1231), .A4(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1055), .B1(new_n1031), .B2(new_n711), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G387), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(G390), .A2(new_n968), .A3(new_n993), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(G393), .B(G396), .Z(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1239), .A2(new_n1242), .A3(new_n1240), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT125), .Z(new_n1247));
  NAND2_X1  g1047(.A1(new_n1236), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT63), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1246), .B1(new_n1224), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(new_n1249), .C2(new_n1224), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1252), .ZN(G405));
  INV_X1    g1053(.A(KEYINPUT126), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT127), .B1(new_n1214), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT127), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1227), .A2(KEYINPUT126), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(new_n1246), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G375), .A2(new_n1202), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n1232), .C1(KEYINPUT126), .C2(new_n1227), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(new_n1259), .B(new_n1261), .ZN(G402));
endmodule


