//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006;
  AND2_X1   g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT41), .ZN(new_n203));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G190gat), .B(G218gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT96), .ZN(new_n208));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209));
  INV_X1    g008(.A(G85gat), .ZN(new_n210));
  INV_X1    g009(.A(G92gat), .ZN(new_n211));
  AOI22_X1  g010(.A1(KEYINPUT8), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(new_n210), .B2(new_n211), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G99gat), .B(G106gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT95), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G43gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G50gat), .ZN(new_n228));
  INV_X1    g027(.A(G50gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G43gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT15), .ZN(new_n231));
  NAND2_X1  g030(.A1(G29gat), .A2(G36gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n226), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(KEYINPUT87), .A2(G50gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT87), .A2(G50gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(new_n227), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n230), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT15), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT88), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT15), .B1(new_n237), .B2(new_n230), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT88), .B1(new_n243), .B2(new_n233), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n246), .B(new_n232), .C1(new_n226), .C2(KEYINPUT86), .ZN(new_n247));
  INV_X1    g046(.A(new_n231), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n220), .A2(new_n250), .B1(KEYINPUT41), .B2(new_n202), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT17), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n218), .B(KEYINPUT95), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n242), .A2(new_n244), .B1(new_n248), .B2(new_n247), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT17), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n208), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT96), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(new_n206), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n251), .A2(new_n257), .A3(KEYINPUT96), .A4(new_n207), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT94), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n205), .B1(new_n262), .B2(KEYINPUT97), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(KEYINPUT97), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT97), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n265), .A3(new_n261), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n263), .B1(new_n267), .B2(new_n205), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G155gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n269), .B(KEYINPUT93), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G15gat), .B(G22gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT16), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(G1gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(G1gat), .B2(new_n272), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n275), .B(G8gat), .Z(new_n276));
  INV_X1    g075(.A(KEYINPUT21), .ZN(new_n277));
  XNOR2_X1  g076(.A(G57gat), .B(G64gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G71gat), .B(G78gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(G71gat), .A2(G78gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G71gat), .A2(G78gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT91), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n278), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT92), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT9), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n278), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n279), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G231gat), .A2(G233gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n294), .B(G183gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n297), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n271), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n293), .A2(new_n277), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(G211gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n304), .B(new_n306), .Z(new_n307));
  NAND3_X1  g106(.A1(new_n299), .A2(new_n301), .A3(new_n271), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n307), .ZN(new_n310));
  INV_X1    g109(.A(new_n308), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(new_n302), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n268), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n315));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(new_n210), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT0), .B(G57gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT76), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT2), .ZN(new_n324));
  OR2_X1    g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G155gat), .B(G162gat), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n327), .A2(KEYINPUT75), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n328), .B1(new_n327), .B2(KEYINPUT75), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n322), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G141gat), .B(G148gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n333), .B1(G155gat), .B2(G162gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT75), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n328), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n327), .A2(KEYINPUT75), .A3(new_n328), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(KEYINPUT3), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(KEYINPUT1), .ZN(new_n343));
  XNOR2_X1  g142(.A(G127gat), .B(G134gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n346));
  INV_X1    g145(.A(G113gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(G120gat), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G113gat), .ZN(new_n350));
  OAI211_X1 g149(.A(KEYINPUT66), .B(new_n346), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n341), .B(new_n344), .C1(new_n342), .C2(KEYINPUT1), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n321), .B1(new_n340), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n354), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n356), .A2(KEYINPUT76), .A3(new_n339), .A4(new_n331), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n337), .A2(new_n338), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT4), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n352), .A2(new_n353), .B1(new_n337), .B2(new_n338), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n366), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n354), .A2(new_n359), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(new_n362), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(KEYINPUT77), .B(new_n368), .C1(new_n369), .C2(new_n362), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n367), .A2(new_n374), .A3(KEYINPUT5), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n368), .B1(new_n355), .B2(new_n357), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT5), .ZN(new_n377));
  OR3_X1    g176(.A1(new_n360), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n361), .A2(KEYINPUT78), .A3(new_n364), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n320), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT6), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n375), .A2(new_n380), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n319), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n375), .A2(new_n320), .A3(new_n380), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n384), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT38), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT73), .B(G64gat), .Z(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT74), .B(G92gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G8gat), .B(G36gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G183gat), .A2(G190gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT64), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT24), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n295), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n401), .B1(new_n399), .B2(new_n400), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(G169gat), .B2(G176gat), .ZN(new_n411));
  INV_X1    g210(.A(G169gat), .ZN(new_n412));
  INV_X1    g211(.A(G176gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT23), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n409), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT25), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT26), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT26), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(G169gat), .B2(G176gat), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n417), .B(new_n399), .C1(new_n419), .C2(new_n408), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n403), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(KEYINPUT65), .A3(KEYINPUT28), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT27), .B(G183gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n427));
  OR2_X1    g226(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n426), .A2(new_n403), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n415), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n404), .A2(KEYINPUT24), .A3(new_n399), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n399), .A2(KEYINPUT24), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT25), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(G226gat), .A2(G233gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n437), .B(KEYINPUT71), .Z(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(G211gat), .ZN(new_n443));
  INV_X1    g242(.A(G218gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(G211gat), .A2(G218gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n444), .A2(KEYINPUT69), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT69), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G218gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n451), .A3(G211gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT22), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G197gat), .B(G204gat), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n448), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n448), .B1(new_n454), .B2(new_n455), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT70), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n447), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n440), .A2(new_n442), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n430), .A2(new_n435), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT25), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n405), .A2(new_n406), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(new_n431), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n441), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n438), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT72), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n442), .A2(KEYINPUT72), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n439), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n464), .B1(new_n475), .B2(new_n463), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n392), .B(new_n398), .C1(new_n476), .C2(KEYINPUT37), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n442), .A2(KEYINPUT72), .ZN(new_n478));
  AOI211_X1 g277(.A(new_n472), .B(new_n438), .C1(new_n436), .C2(new_n441), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n478), .A2(new_n479), .A3(new_n440), .ZN(new_n480));
  INV_X1    g279(.A(new_n463), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n463), .B1(new_n440), .B2(new_n442), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n482), .A2(KEYINPUT37), .A3(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT82), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n464), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(new_n398), .C1(new_n480), .C2(new_n481), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n398), .A2(KEYINPUT37), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n482), .A2(KEYINPUT37), .A3(new_n483), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n392), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n487), .A2(new_n488), .B1(new_n476), .B2(KEYINPUT37), .ZN(new_n494));
  OAI22_X1  g293(.A1(new_n494), .A2(new_n392), .B1(new_n476), .B2(new_n398), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n391), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G228gat), .A2(G233gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n448), .A2(new_n454), .A3(new_n455), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n461), .B1(new_n460), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n457), .A2(KEYINPUT70), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n441), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n359), .B1(new_n502), .B2(new_n322), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(new_n359), .B2(new_n322), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n463), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n498), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G78gat), .B(G106gat), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n359), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT29), .B1(new_n460), .B2(new_n499), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT80), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n322), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI211_X1 g311(.A(KEYINPUT80), .B(KEYINPUT29), .C1(new_n460), .C2(new_n499), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n463), .A2(new_n504), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n497), .A3(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n506), .A2(new_n508), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n508), .B1(new_n506), .B2(new_n516), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(G22gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G50gat), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n517), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n514), .A2(new_n497), .A3(new_n515), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT29), .B1(new_n458), .B2(new_n462), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n509), .B1(new_n525), .B2(KEYINPUT3), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n497), .B1(new_n526), .B2(new_n515), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n507), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n506), .A2(new_n508), .A3(new_n516), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n521), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT40), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT39), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n369), .A2(new_n362), .A3(new_n368), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n358), .A2(new_n378), .A3(new_n379), .ZN(new_n535));
  AOI211_X1 g334(.A(new_n533), .B(new_n534), .C1(new_n535), .C2(new_n368), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n533), .A3(new_n368), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n320), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n532), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n534), .B1(new_n535), .B2(new_n368), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT39), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n541), .A2(KEYINPUT40), .A3(new_n320), .A4(new_n537), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n542), .A3(new_n386), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n476), .B2(new_n398), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n486), .B1(new_n480), .B2(new_n481), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(KEYINPUT30), .A3(new_n397), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n545), .A2(new_n547), .A3(new_n487), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n531), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n315), .B1(new_n496), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n522), .B1(new_n517), .B2(new_n518), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n528), .A2(new_n521), .A3(new_n529), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT81), .ZN(new_n554));
  INV_X1    g353(.A(new_n388), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n555), .A2(new_n381), .A3(KEYINPUT6), .ZN(new_n556));
  INV_X1    g355(.A(new_n382), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n548), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n436), .A2(KEYINPUT67), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT67), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n416), .A2(new_n430), .A3(new_n560), .A4(new_n435), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n356), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G227gat), .A2(G233gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n436), .A2(KEYINPUT67), .A3(new_n354), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT33), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G15gat), .B(G43gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G71gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G99gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n562), .A2(new_n565), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n563), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT34), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n576), .B1(new_n563), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n563), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n573), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n566), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT32), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n571), .B1(new_n566), .B2(new_n567), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n580), .B1(new_n574), .B2(new_n563), .ZN(new_n587));
  AOI211_X1 g386(.A(new_n564), .B(new_n578), .C1(new_n562), .C2(new_n565), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n582), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n585), .B1(new_n582), .B2(new_n589), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n592), .B1(new_n590), .B2(new_n591), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n554), .A2(new_n558), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n539), .A2(new_n542), .A3(new_n386), .ZN(new_n597));
  INV_X1    g396(.A(new_n548), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n553), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n476), .A2(new_n398), .ZN(new_n600));
  INV_X1    g399(.A(new_n494), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(KEYINPUT38), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n602), .A2(new_n389), .A3(new_n384), .A4(new_n390), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n599), .B(KEYINPUT84), .C1(new_n603), .C2(new_n493), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n550), .A2(new_n596), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n582), .A2(new_n589), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n566), .A2(KEYINPUT32), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n582), .A2(new_n585), .A3(new_n589), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n608), .A2(new_n552), .A3(new_n551), .A4(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT35), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n548), .A4(new_n391), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT85), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n614), .B(KEYINPUT35), .C1(new_n558), .C2(new_n610), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n590), .A2(new_n591), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n389), .A2(new_n382), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n531), .A4(new_n548), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n614), .B1(new_n619), .B2(KEYINPUT35), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n613), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n314), .B1(new_n605), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n288), .A2(KEYINPUT98), .A3(new_n292), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT98), .B1(new_n288), .B2(new_n292), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n218), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  INV_X1    g430(.A(new_n218), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n293), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n630), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n293), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n627), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n626), .B1(new_n630), .B2(new_n634), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n625), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n635), .A2(new_n637), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n639), .B1(new_n642), .B2(new_n626), .ZN(new_n643));
  INV_X1    g442(.A(new_n625), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR4_X1   g444(.A1(new_n638), .A2(KEYINPUT99), .A3(new_n639), .A4(new_n625), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g448(.A(KEYINPUT100), .B(new_n640), .C1(new_n645), .C2(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT89), .B1(new_n276), .B2(new_n255), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n275), .B(G8gat), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT89), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n250), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n250), .B2(new_n653), .ZN(new_n657));
  NAND2_X1  g456(.A1(G229gat), .A2(G233gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT13), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n253), .A2(new_n256), .A3(new_n276), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n656), .A2(new_n661), .A3(new_n658), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT90), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n656), .A2(new_n661), .A3(new_n658), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n660), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G113gat), .B(G141gat), .ZN(new_n669));
  INV_X1    g468(.A(G197gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT11), .B(G169gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT12), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n660), .A2(new_n665), .A3(new_n667), .A4(new_n674), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n651), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n622), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n618), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT101), .B(G1gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1324gat));
  INV_X1    g482(.A(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n598), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G8gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT103), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n685), .A2(KEYINPUT102), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(KEYINPUT42), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT16), .B(G8gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR4_X1   g491(.A1(new_n688), .A2(KEYINPUT42), .A3(new_n685), .A4(new_n690), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n687), .B1(new_n692), .B2(new_n693), .ZN(G1325gat));
  INV_X1    g493(.A(G15gat), .ZN(new_n695));
  INV_X1    g494(.A(new_n595), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT104), .B1(new_n696), .B2(new_n593), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n594), .A2(new_n698), .A3(new_n595), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n680), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n617), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n695), .B2(new_n702), .ZN(G1326gat));
  INV_X1    g502(.A(new_n554), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n680), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT105), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n605), .A2(new_n621), .ZN(new_n710));
  INV_X1    g509(.A(new_n263), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n260), .A2(new_n265), .A3(new_n261), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(KEYINPUT97), .B2(new_n262), .ZN(new_n713));
  INV_X1    g512(.A(new_n205), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n709), .B1(new_n710), .B2(new_n715), .ZN(new_n716));
  AOI211_X1 g515(.A(KEYINPUT44), .B(new_n268), .C1(new_n605), .C2(new_n621), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n313), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n679), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n618), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G29gat), .ZN(new_n725));
  AOI211_X1 g524(.A(new_n268), .B(new_n720), .C1(new_n605), .C2(new_n621), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(new_n222), .A3(new_n723), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(KEYINPUT106), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(KEYINPUT106), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(KEYINPUT45), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n725), .A2(new_n730), .A3(new_n733), .ZN(G1328gat));
  NAND3_X1  g533(.A1(new_n726), .A2(new_n223), .A3(new_n598), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT46), .Z(new_n736));
  NAND2_X1  g535(.A1(new_n722), .A2(new_n598), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(new_n223), .ZN(G1329gat));
  NOR2_X1   g538(.A1(new_n696), .A2(new_n593), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n718), .A2(new_n740), .A3(new_n721), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n268), .B1(new_n605), .B2(new_n621), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n743), .A2(new_n227), .A3(new_n617), .A4(new_n721), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n726), .A2(KEYINPUT107), .A3(new_n227), .A4(new_n617), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n742), .A2(KEYINPUT47), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750));
  INV_X1    g549(.A(new_n700), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n721), .C1(new_n716), .C2(new_n717), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G43gat), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n748), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI211_X1 g555(.A(KEYINPUT108), .B(KEYINPUT47), .C1(new_n753), .C2(new_n748), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n749), .B1(new_n756), .B2(new_n757), .ZN(G1330gat));
  OAI211_X1 g557(.A(new_n553), .B(new_n721), .C1(new_n716), .C2(new_n717), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n235), .A3(new_n236), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n235), .A2(new_n236), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n726), .A2(new_n761), .A3(new_n554), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(KEYINPUT48), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT109), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n554), .B(new_n721), .C1(new_n716), .C2(new_n717), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n762), .B1(new_n766), .B2(new_n761), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n760), .A2(new_n762), .A3(new_n770), .A4(KEYINPUT48), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n764), .A2(new_n769), .A3(new_n771), .ZN(G1331gat));
  NAND3_X1  g571(.A1(new_n622), .A2(new_n678), .A3(new_n651), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n723), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g575(.A1(new_n773), .A2(new_n548), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  AND2_X1   g577(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n777), .B2(new_n778), .ZN(G1333gat));
  INV_X1    g580(.A(new_n617), .ZN(new_n782));
  OR3_X1    g581(.A1(new_n773), .A2(KEYINPUT111), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(G71gat), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT111), .B1(new_n773), .B2(new_n782), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n622), .A2(G71gat), .A3(new_n678), .A4(new_n651), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n787), .A2(KEYINPUT110), .A3(new_n700), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT110), .B1(new_n787), .B2(new_n700), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT50), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n786), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n774), .A2(new_n554), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g596(.A1(new_n676), .A2(new_n677), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n313), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT112), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n651), .B(new_n800), .C1(new_n716), .C2(new_n717), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n801), .A2(new_n210), .A3(new_n618), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n743), .A2(new_n800), .ZN(new_n803));
  AND2_X1   g602(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n804));
  NOR2_X1   g603(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n804), .B1(new_n743), .B2(new_n800), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n651), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n723), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n802), .B1(new_n812), .B2(new_n210), .ZN(G1336gat));
  OAI21_X1  g612(.A(G92gat), .B1(new_n801), .B2(new_n548), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n548), .A2(G92gat), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n651), .B(new_n816), .C1(new_n807), .C2(new_n808), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n801), .A2(new_n548), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n803), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT51), .B1(new_n803), .B2(KEYINPUT114), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n651), .A2(new_n816), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n819), .A2(G92gat), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n824), .B2(new_n815), .ZN(G1337gat));
  INV_X1    g624(.A(G99gat), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n826), .A3(new_n617), .ZN(new_n827));
  OAI21_X1  g626(.A(G99gat), .B1(new_n801), .B2(new_n700), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1338gat));
  OAI21_X1  g628(.A(G106gat), .B1(new_n801), .B2(new_n531), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n810), .A2(G106gat), .A3(new_n531), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n830), .B(new_n831), .C1(new_n809), .C2(new_n833), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n801), .A2(new_n704), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n835), .A2(G106gat), .B1(new_n822), .B2(new_n832), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(G1339gat));
  NOR2_X1   g637(.A1(new_n657), .A2(new_n659), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n658), .B1(new_n656), .B2(new_n661), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n673), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n677), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n649), .B2(new_n650), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n642), .A2(new_n626), .ZN(new_n844));
  INV_X1    g643(.A(new_n639), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n644), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT99), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n643), .A2(new_n641), .A3(new_n644), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT54), .B1(new_n642), .B2(new_n626), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n638), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n625), .B1(new_n844), .B2(KEYINPUT54), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n644), .B1(new_n638), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n856), .B(KEYINPUT55), .C1(new_n638), .C2(new_n851), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n849), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n678), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n268), .B1(new_n843), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n842), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n849), .A2(new_n854), .A3(new_n857), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n715), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n313), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n314), .A2(new_n798), .A3(new_n651), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n723), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(new_n610), .A3(new_n598), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n347), .A3(new_n798), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT100), .B1(new_n849), .B2(new_n640), .ZN(new_n869));
  INV_X1    g668(.A(new_n650), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n861), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n862), .A2(new_n798), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n715), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n268), .A2(new_n842), .A3(new_n858), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n719), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n865), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n598), .A2(new_n618), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n554), .A2(new_n782), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G113gat), .B1(new_n880), .B2(new_n678), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n868), .A2(new_n881), .ZN(G1340gat));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n349), .A3(new_n651), .ZN(new_n883));
  OAI21_X1  g682(.A(G120gat), .B1(new_n880), .B2(new_n810), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1341gat));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n313), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(KEYINPUT116), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(KEYINPUT116), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(G127gat), .ZN(new_n889));
  INV_X1    g688(.A(new_n880), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n313), .A2(G127gat), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(G1342gat));
  NOR3_X1   g691(.A1(new_n866), .A2(G134gat), .A3(new_n610), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n268), .A2(new_n598), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT56), .ZN(new_n896));
  OAI21_X1  g695(.A(G134gat), .B1(new_n880), .B2(new_n268), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(KEYINPUT56), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(G1343gat));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n900));
  OAI211_X1 g699(.A(KEYINPUT57), .B(new_n554), .C1(new_n864), .C2(new_n865), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n531), .B1(new_n875), .B2(new_n876), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(KEYINPUT57), .ZN(new_n903));
  INV_X1    g702(.A(new_n740), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n878), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n903), .A2(new_n798), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G141gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n697), .A2(new_n699), .A3(new_n553), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n697), .A2(new_n699), .A3(KEYINPUT117), .A4(new_n553), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n678), .A2(G141gat), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n866), .A2(new_n913), .A3(new_n598), .A4(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n900), .B1(new_n918), .B2(KEYINPUT58), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n916), .B1(new_n907), .B2(G141gat), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT58), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n920), .A2(KEYINPUT118), .A3(new_n921), .ZN(new_n922));
  AND4_X1   g721(.A1(KEYINPUT119), .A2(new_n908), .A3(new_n921), .A4(new_n917), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT119), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  OAI22_X1  g723(.A1(new_n919), .A2(new_n922), .B1(new_n923), .B2(new_n924), .ZN(G1344gat));
  NOR3_X1   g724(.A1(new_n866), .A2(new_n913), .A3(new_n598), .ZN(new_n926));
  INV_X1    g725(.A(G148gat), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n927), .A3(new_n651), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT57), .ZN(new_n930));
  OR3_X1    g729(.A1(new_n268), .A2(KEYINPUT120), .A3(new_n858), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT120), .B1(new_n268), .B2(new_n858), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n861), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n313), .B1(new_n933), .B2(new_n860), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n930), .B(new_n554), .C1(new_n934), .C2(new_n865), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n860), .A2(new_n863), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n865), .B1(new_n936), .B2(new_n719), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT57), .B1(new_n937), .B2(new_n531), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n935), .A2(new_n651), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n906), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n929), .B1(new_n940), .B2(G148gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n930), .B1(new_n937), .B2(new_n531), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n905), .B1(new_n942), .B2(new_n901), .ZN(new_n943));
  AOI211_X1 g742(.A(KEYINPUT59), .B(new_n927), .C1(new_n943), .C2(new_n651), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n928), .B1(new_n941), .B2(new_n944), .ZN(G1345gat));
  INV_X1    g744(.A(G155gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n926), .A2(new_n946), .A3(new_n313), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n943), .A2(new_n313), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n946), .ZN(G1346gat));
  NAND2_X1  g748(.A1(new_n943), .A2(new_n715), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(KEYINPUT121), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(KEYINPUT121), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(G162gat), .A3(new_n952), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n866), .A2(new_n913), .A3(G162gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n894), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1347gat));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n957), .B1(new_n937), .B2(new_n723), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n877), .A2(KEYINPUT122), .A3(new_n618), .ZN(new_n959));
  AOI211_X1 g758(.A(new_n610), .B(new_n548), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n412), .A3(new_n798), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n598), .A2(new_n618), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT123), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n877), .A2(new_n879), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(G169gat), .B1(new_n964), .B2(new_n678), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n961), .A2(new_n965), .ZN(G1348gat));
  NOR3_X1   g765(.A1(new_n964), .A2(new_n413), .A3(new_n810), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n960), .A2(new_n651), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n413), .ZN(G1349gat));
  NAND2_X1  g768(.A1(new_n958), .A2(new_n959), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n313), .A2(new_n426), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n970), .A2(new_n611), .A3(new_n598), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n973));
  OAI21_X1  g772(.A(G183gat), .B1(new_n964), .B2(new_n719), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n976));
  XOR2_X1   g775(.A(new_n975), .B(new_n976), .Z(G1350gat));
  OAI21_X1  g776(.A(G190gat), .B1(new_n964), .B2(new_n268), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT61), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n960), .A2(new_n403), .A3(new_n715), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1351gat));
  AOI211_X1 g780(.A(new_n548), .B(new_n909), .C1(new_n958), .C2(new_n959), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n982), .A2(new_n670), .A3(new_n798), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n700), .A2(new_n963), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n935), .A2(new_n938), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(G197gat), .B1(new_n985), .B2(new_n678), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n983), .A2(new_n986), .ZN(G1352gat));
  XOR2_X1   g786(.A(KEYINPUT125), .B(G204gat), .Z(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n982), .A2(new_n651), .A3(new_n989), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n939), .A2(new_n984), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(new_n988), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n990), .A2(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(G1353gat));
  NAND3_X1  g794(.A1(new_n982), .A2(new_n443), .A3(new_n313), .ZN(new_n996));
  OAI21_X1  g795(.A(G211gat), .B1(new_n985), .B2(new_n719), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT63), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n996), .B1(new_n999), .B2(new_n1000), .ZN(G1354gat));
  AOI21_X1  g800(.A(G218gat), .B1(new_n982), .B2(new_n715), .ZN(new_n1002));
  OR2_X1    g801(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n268), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n449), .A2(new_n451), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1355gat));
endmodule


