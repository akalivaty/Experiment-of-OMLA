//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G20), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR3_X1   g0012(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT0), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n207), .A2(new_n210), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G68), .A2(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n221), .B(new_n222), .C1(new_n202), .C2(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n220), .B(new_n224), .C1(G97), .C2(G257), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(G1), .B2(G20), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n216), .B(new_n228), .C1(new_n215), .C2(new_n214), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  OR2_X1    g0044(.A1(KEYINPUT3), .A2(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G222), .ZN(new_n249));
  INV_X1    g0049(.A(G223), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n247), .B(new_n249), .C1(new_n250), .C2(new_n248), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n251), .B(new_n252), .C1(G77), .C2(new_n247), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT66), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT66), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G33), .A3(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n257), .A3(new_n209), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G226), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n253), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G169), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n212), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT67), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT67), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(new_n212), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n203), .A2(G20), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n275), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n208), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G13), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G1), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G20), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G50), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n284), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(new_n211), .A3(G20), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n288), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n292), .B1(new_n211), .B2(G20), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G50), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n285), .A2(new_n290), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n267), .B(new_n298), .C1(G179), .C2(new_n265), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT69), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(KEYINPUT3), .A2(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT3), .A2(G33), .ZN(new_n303));
  OAI211_X1 g0103(.A(G232), .B(new_n248), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT70), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n247), .A2(new_n306), .A3(G232), .A4(new_n248), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n302), .A2(new_n303), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G107), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n247), .A2(G238), .A3(G1698), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n305), .A2(new_n307), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n263), .B1(new_n311), .B2(new_n252), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n260), .A2(G244), .ZN(new_n313));
  AOI21_X1  g0113(.A(G169), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n296), .A2(G77), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT15), .B(G87), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n278), .A2(new_n273), .B1(new_n316), .B2(new_n268), .ZN(new_n317));
  INV_X1    g0117(.A(G77), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n212), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n284), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n288), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n318), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n315), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n312), .A2(new_n313), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT71), .B1(new_n325), .B2(G179), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT71), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n312), .A2(new_n327), .A3(new_n328), .A4(new_n313), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n314), .B(new_n324), .C1(new_n326), .C2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n301), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n247), .A2(G232), .A3(G1698), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n247), .A2(G226), .A3(new_n248), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G97), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n263), .B1(new_n335), .B2(new_n252), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n260), .A2(G238), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(KEYINPUT13), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n336), .B2(new_n337), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT14), .B1(new_n342), .B2(new_n266), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n338), .B(KEYINPUT13), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(G169), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n343), .B(new_n346), .C1(new_n328), .C2(new_n344), .ZN(new_n347));
  INV_X1    g0147(.A(G68), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n272), .A2(G77), .B1(G20), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n277), .A2(G50), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n291), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n287), .A2(G20), .A3(new_n348), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT12), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n296), .A2(G68), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n352), .A2(new_n354), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  XOR2_X1   g0157(.A(new_n357), .B(KEYINPUT75), .Z(new_n358));
  NAND2_X1  g0158(.A1(new_n347), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(G200), .B1(new_n339), .B2(new_n341), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT74), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(KEYINPUT74), .B(G200), .C1(new_n339), .C2(new_n341), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n357), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n342), .A2(G190), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n325), .A2(G200), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n312), .A2(G190), .A3(new_n313), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n324), .A3(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n331), .A2(new_n359), .A3(new_n366), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n282), .A2(new_n284), .B1(new_n296), .B2(G50), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT9), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(new_n290), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n265), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n265), .A2(G200), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n373), .B1(new_n372), .B2(new_n290), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n280), .B1(new_n272), .B2(new_n274), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n291), .B1(new_n384), .B2(new_n276), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n294), .A2(new_n202), .A3(new_n295), .ZN(new_n386));
  NOR4_X1   g0186(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT9), .A4(new_n289), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n377), .B(KEYINPUT72), .C1(new_n383), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n379), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT72), .B1(new_n375), .B2(new_n377), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT10), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT73), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT73), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n393), .B(KEYINPUT10), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n382), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n288), .A2(new_n273), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n296), .B2(new_n273), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n245), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n246), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT76), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n308), .A2(new_n400), .A3(KEYINPUT7), .A4(new_n212), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n245), .A2(new_n212), .A3(new_n246), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G68), .ZN(new_n406));
  INV_X1    g0206(.A(G58), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(new_n348), .ZN(new_n408));
  OAI21_X1  g0208(.A(G20), .B1(new_n408), .B2(new_n201), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n277), .A2(G159), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT16), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT7), .B1(new_n308), .B2(new_n212), .ZN(new_n414));
  INV_X1    g0214(.A(new_n398), .ZN(new_n415));
  OAI21_X1  g0215(.A(G68), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(KEYINPUT16), .A3(new_n412), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n284), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n397), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT77), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n411), .B1(new_n405), .B2(G68), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n284), .B(new_n417), .C1(new_n421), .C2(KEYINPUT16), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT77), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n397), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n250), .A2(new_n248), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n223), .A2(G1698), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n426), .B(new_n427), .C1(new_n302), .C2(new_n303), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT78), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT78), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n428), .A2(new_n432), .A3(new_n429), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n252), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n260), .A2(G232), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n264), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G169), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n434), .A2(G179), .A3(new_n435), .A4(new_n264), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n425), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT18), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n436), .A2(G200), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n434), .A2(G190), .A3(new_n435), .A4(new_n264), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n442), .A2(new_n422), .A3(new_n443), .A4(new_n397), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT17), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n425), .A2(new_n446), .A3(new_n439), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n370), .A2(new_n395), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n405), .A2(G107), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n451));
  INV_X1    g0251(.A(G97), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(G107), .ZN(new_n453));
  XNOR2_X1  g0253(.A(G97), .B(G107), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(G20), .C1(new_n454), .C2(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n277), .A2(G77), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n450), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT80), .B1(new_n457), .B2(new_n284), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(KEYINPUT80), .A3(new_n284), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G1), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n258), .A2(new_n466), .A3(G257), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G250), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n245), .B2(new_n246), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT4), .ZN(new_n471));
  OAI21_X1  g0271(.A(G1698), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(G244), .B1(new_n302), .B2(new_n303), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(new_n471), .B1(G33), .B2(G283), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n247), .A2(KEYINPUT4), .A3(G244), .A4(new_n248), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n468), .B1(new_n476), .B2(new_n252), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT81), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n463), .B(G274), .C1(new_n465), .C2(new_n464), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g0281(.A(G190), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n288), .A2(G97), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n211), .A2(G33), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n291), .A2(new_n288), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n483), .B1(new_n486), .B2(G97), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n476), .A2(new_n252), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n479), .A3(new_n467), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G200), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n461), .A2(new_n482), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n457), .A2(KEYINPUT80), .A3(new_n284), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n487), .B1(new_n492), .B2(new_n458), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(KEYINPUT81), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(new_n266), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n477), .A2(new_n328), .A3(new_n479), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n212), .B(G87), .C1(new_n302), .C2(new_n303), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n247), .A2(new_n502), .A3(new_n212), .A4(G87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n505));
  INV_X1    g0305(.A(G107), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n507), .B(KEYINPUT23), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AND4_X1   g0309(.A1(new_n499), .A2(new_n504), .A3(new_n505), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n501), .B2(new_n503), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n499), .B1(new_n511), .B2(new_n505), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n284), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n507), .A2(G1), .A3(new_n286), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n485), .A2(new_n506), .B1(new_n515), .B2(KEYINPUT25), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n258), .A2(new_n466), .A3(G264), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G294), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n247), .B1(G257), .B2(new_n248), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G250), .A2(G1698), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n519), .B1(new_n523), .B2(new_n252), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n479), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G190), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(G200), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n515), .A2(KEYINPUT25), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n518), .A2(new_n527), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n491), .A2(new_n498), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n258), .A2(new_n466), .A3(G270), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n248), .A2(G257), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G264), .A2(G1698), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(new_n302), .C2(new_n303), .ZN(new_n535));
  INV_X1    g0335(.A(G303), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n245), .A2(new_n536), .A3(new_n246), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n252), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n532), .A2(new_n538), .A3(new_n479), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n532), .A2(new_n538), .A3(KEYINPUT83), .A4(new_n479), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(new_n376), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n321), .A2(new_n218), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n291), .A2(new_n288), .A3(G116), .A4(new_n484), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n283), .A2(new_n208), .B1(G20), .B2(new_n218), .ZN(new_n547));
  AOI21_X1  g0347(.A(G20), .B1(G33), .B2(G283), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G33), .B2(new_n452), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n547), .A2(new_n549), .A3(KEYINPUT20), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT20), .B1(new_n547), .B2(new_n549), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n545), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n541), .A2(new_n542), .ZN(new_n554));
  INV_X1    g0354(.A(G200), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n544), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g0357(.A(new_n557), .B(KEYINPUT84), .Z(new_n558));
  NAND3_X1  g0358(.A1(new_n247), .A2(new_n212), .A3(G68), .ZN(new_n559));
  XOR2_X1   g0359(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n560));
  NOR2_X1   g0360(.A1(new_n268), .A2(new_n452), .ZN(new_n561));
  INV_X1    g0361(.A(new_n334), .ZN(new_n562));
  AOI21_X1  g0362(.A(G20), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NOR3_X1   g0363(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n564));
  OAI221_X1 g0364(.A(new_n559), .B1(new_n560), .B2(new_n561), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n284), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n321), .A2(new_n316), .ZN(new_n567));
  INV_X1    g0367(.A(new_n316), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n486), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n247), .A2(G238), .A3(new_n248), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G116), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n248), .C2(new_n473), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n252), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n463), .A2(G274), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n258), .B(G250), .C1(G1), .C2(new_n462), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n266), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n574), .A2(new_n328), .A3(new_n575), .A4(new_n576), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n570), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n541), .A2(G169), .A3(new_n552), .A4(new_n542), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT21), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n539), .A2(new_n328), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(new_n553), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n513), .A2(new_n529), .A3(new_n517), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n525), .A2(new_n266), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n526), .A2(new_n328), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n577), .A2(G200), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n565), .A2(new_n284), .B1(new_n321), .B2(new_n316), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n574), .A2(G190), .A3(new_n575), .A4(new_n576), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n486), .A2(G87), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  AND4_X1   g0396(.A1(new_n580), .A2(new_n587), .A3(new_n591), .A4(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n449), .A2(new_n531), .A3(new_n558), .A4(new_n597), .ZN(G372));
  NAND2_X1  g0398(.A1(new_n392), .A2(new_n394), .ZN(new_n599));
  INV_X1    g0399(.A(new_n382), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT88), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT88), .ZN(new_n602));
  AOI211_X1 g0402(.A(new_n602), .B(new_n382), .C1(new_n392), .C2(new_n394), .ZN(new_n603));
  OR2_X1    g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n439), .A2(new_n419), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT87), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT87), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n439), .A2(new_n419), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n446), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(KEYINPUT18), .A3(new_n608), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n366), .A2(new_n330), .B1(new_n358), .B2(new_n347), .ZN(new_n613));
  INV_X1    g0413(.A(new_n445), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n301), .B1(new_n604), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n596), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n587), .A2(new_n591), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(new_n491), .A3(new_n498), .A4(new_n530), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n496), .A2(new_n497), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT86), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n496), .A2(KEYINPUT86), .A3(new_n497), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n493), .A4(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n617), .B1(new_n619), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT26), .B1(new_n498), .B2(new_n617), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n580), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n449), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n616), .A2(new_n629), .ZN(G369));
  NOR2_X1   g0430(.A1(new_n286), .A2(G20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n211), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n552), .ZN(new_n638));
  OR3_X1    g0438(.A1(new_n587), .A2(KEYINPUT89), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n558), .A2(new_n638), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT89), .B1(new_n640), .B2(new_n587), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n587), .A2(new_n638), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G330), .ZN(new_n644));
  INV_X1    g0444(.A(new_n591), .ZN(new_n645));
  INV_X1    g0445(.A(new_n637), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n588), .A2(new_n637), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n645), .B1(new_n530), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n644), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n648), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n587), .A2(new_n637), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n647), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n651), .A2(new_n655), .ZN(G399));
  INV_X1    g0456(.A(new_n213), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G41), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n564), .A2(new_n218), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(G1), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n206), .B2(new_n659), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT28), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n531), .A2(new_n558), .A3(new_n597), .A4(new_n646), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n494), .A2(new_n495), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n577), .A2(new_n585), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n524), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT30), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n666), .A2(KEYINPUT30), .A3(new_n524), .A4(new_n667), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n543), .A2(new_n328), .A3(new_n577), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT90), .Z(new_n673));
  NAND2_X1  g0473(.A1(new_n489), .A2(new_n525), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n670), .B(new_n671), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n637), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n665), .A2(new_n676), .A3(KEYINPUT31), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT31), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n678), .A3(new_n637), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n646), .B1(new_n626), .B2(new_n628), .ZN(new_n682));
  XOR2_X1   g0482(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n622), .A2(new_n493), .A3(new_n596), .A4(new_n624), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT26), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n580), .ZN(new_n688));
  INV_X1    g0488(.A(new_n498), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n623), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n617), .B1(new_n619), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n646), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n684), .B1(new_n685), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n681), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n664), .B1(new_n694), .B2(G1), .ZN(G364));
  AOI21_X1  g0495(.A(new_n208), .B1(G20), .B2(new_n266), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n555), .A2(G179), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n212), .A2(G190), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(G179), .A2(G200), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(G283), .A2(new_n700), .B1(new_n703), .B2(G329), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n212), .A2(new_n376), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n328), .A2(new_n555), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G326), .ZN(new_n709));
  INV_X1    g0509(.A(G311), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n328), .A2(G200), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n698), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n704), .B(new_n709), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n705), .A2(new_n697), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n247), .B1(new_n715), .B2(G303), .ZN(new_n716));
  INV_X1    g0516(.A(G294), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n212), .B1(new_n701), .B2(G190), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n706), .A2(new_n698), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT33), .B(G317), .Z(new_n720));
  OAI221_X1 g0520(.A(new_n716), .B1(new_n717), .B2(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n705), .A2(new_n711), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI211_X1 g0523(.A(new_n713), .B(new_n721), .C1(G322), .C2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n712), .ZN(new_n725));
  AOI22_X1  g0525(.A1(G50), .A2(new_n708), .B1(new_n725), .B2(G77), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n715), .A2(G87), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n726), .B(new_n727), .C1(new_n506), .C2(new_n699), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n719), .A2(new_n348), .B1(new_n718), .B2(new_n452), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT93), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n722), .A2(new_n407), .ZN(new_n731));
  INV_X1    g0531(.A(G159), .ZN(new_n732));
  OR3_X1    g0532(.A1(new_n702), .A2(KEYINPUT32), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT32), .B1(new_n702), .B2(new_n732), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n247), .A3(new_n734), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n728), .A2(new_n730), .A3(new_n731), .A4(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n696), .B1(new_n724), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n631), .A2(G45), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n659), .A2(G1), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n207), .A2(G45), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n657), .A2(new_n247), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n741), .B(new_n742), .C1(new_n462), .C2(new_n240), .ZN(new_n743));
  INV_X1    g0543(.A(G355), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n247), .A2(new_n213), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT92), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n743), .B1(G116), .B2(new_n213), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n696), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n737), .A2(new_n740), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT94), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n750), .B(KEYINPUT95), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n643), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n754), .B2(new_n753), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT96), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n740), .B1(new_n643), .B2(G330), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G330), .B2(new_n643), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n761), .ZN(G396));
  NAND2_X1  g0562(.A1(new_n619), .A2(new_n625), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n596), .ZN(new_n764));
  INV_X1    g0564(.A(new_n628), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n637), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n326), .A2(new_n329), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n325), .A2(new_n266), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n767), .A2(new_n768), .A3(new_n323), .A4(new_n646), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT99), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n324), .B1(new_n326), .B2(new_n329), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n323), .A2(new_n637), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n772), .A2(new_n768), .B1(new_n369), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n368), .A2(new_n324), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n555), .B1(new_n312), .B2(new_n313), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n772), .B2(new_n768), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n771), .A2(new_n774), .B1(new_n778), .B2(new_n770), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT100), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n777), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n769), .B(new_n770), .C1(new_n330), .C2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(KEYINPUT99), .B1(new_n330), .B2(new_n777), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n783), .A2(KEYINPUT100), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n766), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n785), .ZN(new_n788));
  AOI21_X1  g0588(.A(KEYINPUT100), .B1(new_n783), .B2(new_n784), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n682), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n681), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(KEYINPUT101), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n792), .A2(new_n681), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(KEYINPUT101), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n739), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT102), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n786), .A2(new_n749), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n719), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G143), .A2(new_n723), .B1(new_n802), .B2(G150), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n803), .B1(new_n804), .B2(new_n707), .C1(new_n732), .C2(new_n712), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT34), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n308), .B1(new_n703), .B2(G132), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n807), .A2(KEYINPUT98), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(KEYINPUT98), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n700), .A2(G68), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n407), .B2(new_n718), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n806), .B(new_n812), .C1(new_n202), .C2(new_n714), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n714), .A2(new_n506), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n308), .B1(new_n712), .B2(new_n218), .C1(new_n815), .C2(new_n719), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n700), .A2(G87), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n710), .B2(new_n702), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n816), .B(new_n818), .C1(G303), .C2(new_n708), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n722), .A2(new_n717), .B1(new_n718), .B2(new_n452), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(KEYINPUT97), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n820), .A2(KEYINPUT97), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n813), .B1(new_n814), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n696), .A2(new_n748), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n824), .A2(new_n696), .B1(new_n318), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n739), .B1(new_n801), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n798), .A2(new_n799), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n799), .B1(new_n798), .B2(new_n828), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(G384));
  INV_X1    g0631(.A(KEYINPUT108), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT16), .B1(new_n416), .B2(new_n412), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n397), .B1(new_n418), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n635), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n439), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n444), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT37), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT103), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n837), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n444), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n425), .B2(new_n439), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT104), .B1(new_n425), .B2(new_n835), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT104), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n847), .B(new_n635), .C1(new_n420), .C2(new_n424), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n845), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT105), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(KEYINPUT105), .B(new_n845), .C1(new_n846), .C2(new_n848), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n842), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n448), .A2(new_n835), .A3(new_n834), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n846), .A2(new_n848), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n444), .A2(KEYINPUT106), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n444), .A2(KEYINPUT106), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(new_n606), .A3(new_n608), .A4(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n852), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n422), .A2(new_n423), .A3(new_n397), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n423), .B1(new_n422), .B2(new_n397), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n835), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n847), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n425), .A2(KEYINPUT104), .A3(new_n835), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT105), .B1(new_n868), .B2(new_n845), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n861), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n610), .A2(new_n445), .A3(new_n611), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n857), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n832), .B1(new_n856), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n858), .A2(new_n608), .A3(new_n606), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n868), .A2(new_n875), .A3(new_n859), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n851), .A2(new_n852), .B1(new_n876), .B2(KEYINPUT37), .ZN(new_n877));
  INV_X1    g0677(.A(new_n872), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n854), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n840), .A2(new_n841), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n862), .B2(new_n869), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n448), .A2(new_n835), .A3(new_n834), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(KEYINPUT108), .A3(new_n883), .ZN(new_n884));
  AOI221_X4 g0684(.A(new_n357), .B1(G190), .B2(new_n342), .C1(new_n362), .C2(new_n363), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n358), .B(new_n637), .C1(new_n885), .C2(new_n347), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n358), .A2(new_n637), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n359), .A2(new_n366), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n677), .A2(new_n786), .A3(new_n889), .A4(new_n679), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n874), .A2(new_n884), .A3(new_n892), .ZN(new_n893));
  AND4_X1   g0693(.A1(new_n677), .A2(new_n786), .A3(new_n889), .A4(new_n679), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n881), .B2(new_n882), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n894), .B1(new_n856), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n891), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n680), .A2(new_n449), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n898), .B(new_n899), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n684), .B(new_n449), .C1(new_n685), .C2(new_n692), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n616), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT107), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n901), .B(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n856), .B2(new_n873), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n359), .A2(new_n637), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n854), .B1(new_n853), .B2(new_n855), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n883), .A3(KEYINPUT39), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n612), .A2(new_n835), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n769), .B1(new_n790), .B2(new_n682), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n889), .C1(new_n856), .C2(new_n895), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n905), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n211), .B2(new_n631), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n453), .B1(new_n454), .B2(new_n451), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT35), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n210), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(G116), .C1(new_n919), .C2(new_n918), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT36), .ZN(new_n922));
  OAI21_X1  g0722(.A(G77), .B1(new_n407), .B2(new_n348), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n923), .A2(new_n206), .B1(G50), .B2(new_n348), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n286), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n917), .A2(new_n922), .A3(new_n925), .ZN(G367));
  NAND4_X1  g0726(.A1(new_n622), .A2(new_n493), .A3(new_n624), .A4(new_n637), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT111), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n493), .A2(new_n637), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n491), .A2(new_n498), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n651), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n654), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT42), .Z(new_n935));
  AOI21_X1  g0735(.A(new_n689), .B1(new_n931), .B2(new_n645), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n637), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT110), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n646), .B1(new_n593), .B2(new_n595), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT109), .ZN(new_n940));
  INV_X1    g0740(.A(new_n580), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n940), .A2(new_n941), .A3(new_n617), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n938), .B2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n932), .B1(new_n937), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n937), .A2(new_n932), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n951), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n953), .A2(new_n948), .B1(KEYINPUT43), .B2(new_n946), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n658), .B(KEYINPUT41), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n931), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n655), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT44), .ZN(new_n959));
  INV_X1    g0759(.A(new_n655), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n960), .A2(KEYINPUT45), .A3(new_n931), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT45), .B1(new_n960), .B2(new_n931), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n959), .A2(new_n651), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n651), .B1(new_n959), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n652), .A2(new_n653), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n933), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n644), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n643), .B(G330), .C1(new_n933), .C2(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n964), .A2(new_n694), .A3(new_n965), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n956), .B1(new_n971), .B2(new_n694), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n738), .A2(G1), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n952), .B(new_n954), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n742), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n751), .B1(new_n213), .B2(new_n316), .C1(new_n236), .C2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n718), .A2(new_n506), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n308), .B1(new_n699), .B2(new_n452), .C1(new_n717), .C2(new_n719), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(G283), .C2(new_n725), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT112), .B1(new_n714), .B2(new_n218), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT46), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT46), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G311), .A2(new_n708), .B1(new_n723), .B2(G303), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(G317), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n979), .B(new_n984), .C1(new_n985), .C2(new_n702), .ZN(new_n986));
  INV_X1    g0786(.A(G143), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n707), .A2(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n719), .A2(new_n732), .B1(new_n702), .B2(new_n804), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G50), .B2(new_n725), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n247), .B1(new_n722), .B2(new_n279), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G77), .B2(new_n700), .ZN(new_n992));
  INV_X1    g0792(.A(new_n718), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(G68), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n715), .A2(G58), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n992), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n986), .B1(new_n988), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT47), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n739), .B1(new_n998), .B2(new_n696), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n976), .B(new_n999), .C1(new_n946), .C2(new_n756), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n974), .A2(new_n1000), .ZN(G387));
  AOI21_X1  g0801(.A(new_n659), .B1(new_n970), .B2(new_n694), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT115), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(KEYINPUT115), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n1004), .C1(new_n694), .C2(new_n970), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n970), .A2(new_n973), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n696), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n708), .A2(G322), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n802), .A2(G311), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n723), .A2(G317), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n725), .A2(G303), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n1014));
  AOI22_X1  g0814(.A1(new_n1013), .A2(new_n1014), .B1(G283), .B2(new_n993), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n717), .B2(new_n714), .C1(new_n1014), .C2(new_n1013), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n703), .A2(G326), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n247), .B1(new_n700), .B2(G116), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n718), .A2(new_n316), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n247), .B1(new_n699), .B2(new_n452), .C1(new_n202), .C2(new_n722), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(G68), .C2(new_n725), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n715), .A2(G77), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n273), .B2(new_n719), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT113), .B1(new_n707), .B2(new_n732), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n707), .A2(KEYINPUT113), .A3(new_n732), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1025), .B(new_n1030), .C1(new_n279), .C2(new_n702), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1007), .B1(new_n1022), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n742), .B1(new_n233), .B2(new_n462), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n661), .B2(new_n746), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n348), .A2(new_n318), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n274), .A2(new_n202), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n660), .B1(new_n1036), .B2(KEYINPUT50), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n462), .C1(KEYINPUT50), .C2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1034), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(G107), .B2(new_n213), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1032), .B1(new_n751), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n740), .C1(new_n652), .C2(new_n756), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1005), .A2(new_n1006), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT116), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1005), .A2(KEYINPUT116), .A3(new_n1006), .A4(new_n1042), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(G393));
  OAI221_X1 g0847(.A(new_n751), .B1(new_n452), .B2(new_n213), .C1(new_n243), .C2(new_n975), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n712), .A2(new_n273), .B1(new_n702), .B2(new_n987), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G50), .B2(new_n802), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n348), .B2(new_n714), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n718), .A2(new_n318), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n707), .A2(new_n279), .B1(new_n722), .B2(new_n732), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1053), .A2(new_n247), .A3(new_n817), .A4(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n308), .B1(new_n699), .B2(new_n506), .C1(new_n815), .C2(new_n714), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G322), .B2(new_n703), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT117), .Z(new_n1059));
  OAI22_X1  g0859(.A1(new_n707), .A2(new_n985), .B1(new_n722), .B2(new_n710), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n802), .A2(G303), .B1(new_n993), .B2(G116), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n712), .A2(new_n717), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1056), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n739), .B1(new_n1065), .B2(new_n696), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n750), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1048), .B(new_n1066), .C1(new_n931), .C2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n964), .A2(new_n965), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n973), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n970), .A2(new_n694), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n659), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1071), .B1(new_n971), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G390));
  AOI21_X1  g0875(.A(new_n908), .B1(new_n913), .B2(new_n889), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n910), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT39), .B1(new_n879), .B2(new_n883), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n769), .B1(new_n692), .B2(new_n790), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n908), .B1(new_n1081), .B2(new_n889), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n874), .A2(new_n1082), .A3(new_n884), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n680), .A2(G330), .A3(new_n786), .A4(new_n889), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1084), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n1070), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n749), .B1(new_n907), .B2(new_n910), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n699), .A2(new_n202), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n714), .A2(new_n279), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT53), .Z(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT54), .B(G143), .Z(new_n1093));
  AOI211_X1 g0893(.A(new_n1090), .B(new_n1092), .C1(new_n725), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(G132), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n722), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(G128), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n247), .B1(new_n719), .B2(new_n804), .C1(new_n1097), .C2(new_n707), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1096), .B(new_n1098), .C1(G159), .C2(new_n993), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G125), .B2(new_n703), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G107), .A2(new_n802), .B1(new_n703), .B2(G294), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n452), .B2(new_n712), .C1(new_n815), .C2(new_n707), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n723), .A2(G116), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n727), .A2(new_n1104), .A3(new_n810), .A4(new_n308), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1103), .A2(new_n1052), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n696), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n825), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1107), .B1(new_n274), .B2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1089), .A2(new_n739), .A3(new_n1109), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1088), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n677), .A2(new_n786), .A3(G330), .A4(new_n679), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n889), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n874), .A2(new_n1082), .A3(new_n884), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1076), .B1(new_n907), .B2(new_n910), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n680), .A2(new_n449), .A3(G330), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n616), .A2(new_n1118), .A3(new_n902), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n913), .B1(new_n1120), .B2(new_n1114), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1081), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1084), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1119), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1117), .A2(new_n1085), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT118), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n658), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1126), .B2(new_n658), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1125), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1131), .A2(KEYINPUT119), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT119), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1125), .A2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n1132), .A2(new_n1134), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1111), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(G378));
  NAND3_X1  g0937(.A1(new_n893), .A2(G330), .A3(new_n897), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n299), .B1(new_n601), .B2(new_n603), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT55), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT55), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(new_n299), .C1(new_n601), .C2(new_n603), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n298), .A2(new_n835), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT56), .Z(new_n1144));
  AND3_X1   g0944(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1149), .A2(G330), .A3(new_n897), .A4(new_n893), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n915), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1148), .A2(new_n1150), .A3(new_n915), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(KEYINPUT120), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n915), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT120), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1119), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1126), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1155), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1126), .A2(new_n1160), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1148), .A2(new_n915), .A3(new_n1150), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n1156), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n1159), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1162), .A2(new_n1166), .A3(new_n658), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1149), .A2(new_n748), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n825), .A2(new_n202), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n722), .A2(new_n1097), .B1(new_n718), .B2(new_n279), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n715), .A2(new_n1093), .B1(new_n725), .B2(G137), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1095), .B2(new_n719), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G125), .C2(new_n708), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT59), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n703), .B2(G124), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G33), .B1(new_n700), .B2(G159), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n202), .B1(new_n302), .B2(G41), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G116), .A2(new_n708), .B1(new_n802), .B2(G97), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n407), .B2(new_n699), .C1(new_n815), .C2(new_n702), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G107), .A2(new_n723), .B1(new_n725), .B2(new_n568), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n994), .A3(new_n1026), .ZN(new_n1182));
  NOR4_X1   g0982(.A1(new_n1180), .A2(G41), .A3(new_n247), .A4(new_n1182), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT58), .Z(new_n1184));
  NAND3_X1  g0984(.A1(new_n1177), .A2(new_n1178), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n739), .B1(new_n1185), .B2(new_n696), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1168), .A2(new_n1169), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1189), .B2(new_n973), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1167), .A2(new_n1190), .ZN(G375));
  AOI21_X1  g0991(.A(new_n1070), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n722), .A2(new_n804), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n707), .A2(new_n1095), .B1(new_n712), .B2(new_n279), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n802), .C2(new_n1093), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n247), .B1(new_n702), .B2(new_n1097), .C1(new_n407), .C2(new_n699), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G50), .B2(new_n993), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(new_n732), .C2(new_n714), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G294), .A2(new_n708), .B1(new_n725), .B2(G107), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n218), .B2(new_n719), .C1(new_n815), .C2(new_n722), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G77), .B2(new_n700), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n714), .A2(new_n452), .B1(new_n702), .B2(new_n536), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT121), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n316), .C2(new_n718), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1198), .B1(new_n1204), .B2(new_n247), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n696), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(G68), .B2(new_n1108), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1113), .B2(new_n748), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1192), .B1(new_n740), .B2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1121), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1209), .B1(new_n1211), .B2(new_n956), .ZN(G381));
  INV_X1    g1012(.A(G396), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1045), .A2(new_n1213), .A3(new_n1046), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(G384), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n974), .A2(new_n1000), .A3(new_n1074), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1167), .A2(new_n1136), .A3(new_n1190), .ZN(new_n1219));
  OR4_X1    g1019(.A1(G381), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(G407));
  OAI211_X1 g1020(.A(G407), .B(G213), .C1(G343), .C2(new_n1219), .ZN(G409));
  INV_X1    g1021(.A(KEYINPUT126), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT62), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G375), .A2(G378), .ZN(new_n1226));
  INV_X1    g1026(.A(G213), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(G343), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1126), .A2(new_n658), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT118), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1126), .A2(new_n1127), .A3(new_n658), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1135), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1088), .A2(new_n1110), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1187), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1155), .A2(new_n973), .A3(new_n1158), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1189), .A2(new_n955), .A3(new_n1163), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1228), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1226), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1210), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT60), .B1(new_n1240), .B2(KEYINPUT122), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT122), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1210), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n658), .A3(new_n1131), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1209), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1216), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(G384), .A2(new_n1209), .A3(new_n1245), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1224), .B(new_n1225), .C1(new_n1239), .C2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1228), .A2(G2897), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1246), .B(G384), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1228), .A2(KEYINPUT124), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  AND4_X1   g1054(.A1(new_n1251), .A2(new_n1247), .A3(new_n1253), .A4(new_n1248), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1239), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1136), .B1(new_n1167), .B2(new_n1190), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1228), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1232), .A2(new_n1233), .A3(new_n1187), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1259), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1264), .A2(new_n1222), .A3(new_n1223), .A4(new_n1252), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1250), .A2(new_n1257), .A3(new_n1258), .A4(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1213), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1218), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1074), .B1(new_n974), .B2(new_n1000), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1268), .B(new_n1214), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G387), .A2(G390), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1272), .B(new_n1218), .C1(new_n1215), .C2(new_n1267), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1266), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT125), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1226), .A2(new_n1238), .A3(KEYINPUT123), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1259), .B2(new_n1263), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1279), .A3(new_n1256), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(KEYINPUT63), .B1(new_n1239), .B2(new_n1249), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1264), .A2(new_n1285), .A3(new_n1252), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT61), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1276), .B1(new_n1283), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1285), .B1(new_n1264), .B2(new_n1252), .ZN(new_n1289));
  NOR4_X1   g1089(.A1(new_n1259), .A2(new_n1263), .A3(KEYINPUT63), .A4(new_n1249), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1258), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1291), .A2(new_n1282), .A3(KEYINPUT125), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1275), .B1(new_n1288), .B2(new_n1292), .ZN(G405));
  XNOR2_X1  g1093(.A(new_n1274), .B(KEYINPUT127), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1226), .A2(new_n1219), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(new_n1249), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1294), .B(new_n1296), .ZN(G402));
endmodule


