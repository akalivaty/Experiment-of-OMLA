

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  AND2_X1 U322 ( .A1(G232GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U323 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n330) );
  XNOR2_X1 U324 ( .A(n331), .B(n330), .ZN(n362) );
  XNOR2_X1 U325 ( .A(n338), .B(n337), .ZN(n339) );
  INV_X1 U326 ( .A(KEYINPUT103), .ZN(n328) );
  XNOR2_X1 U327 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U328 ( .A(n313), .B(n290), .ZN(n314) );
  XNOR2_X1 U329 ( .A(n328), .B(KEYINPUT36), .ZN(n329) );
  XNOR2_X1 U330 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U331 ( .A(n315), .B(n314), .ZN(n319) );
  XNOR2_X1 U332 ( .A(n560), .B(n329), .ZN(n580) );
  XNOR2_X1 U333 ( .A(n347), .B(n346), .ZN(n364) );
  XNOR2_X1 U334 ( .A(G183GAT), .B(KEYINPUT124), .ZN(n454) );
  XNOR2_X1 U335 ( .A(n455), .B(n454), .ZN(G1350GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n292) );
  XNOR2_X1 U337 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n292), .B(n291), .ZN(n300) );
  NAND2_X1 U339 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XOR2_X1 U340 ( .A(G64GAT), .B(G78GAT), .Z(n294) );
  XNOR2_X1 U341 ( .A(G155GAT), .B(G211GAT), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n296) );
  XOR2_X1 U343 ( .A(G183GAT), .B(G127GAT), .Z(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n308) );
  XNOR2_X1 U347 ( .A(G15GAT), .B(G22GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n301), .B(KEYINPUT67), .ZN(n350) );
  XOR2_X1 U349 ( .A(KEYINPUT12), .B(G57GAT), .Z(n303) );
  XNOR2_X1 U350 ( .A(G8GAT), .B(G1GAT), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n350), .B(n304), .ZN(n306) );
  XOR2_X1 U353 ( .A(G71GAT), .B(KEYINPUT69), .Z(n305) );
  XOR2_X1 U354 ( .A(KEYINPUT13), .B(n305), .Z(n338) );
  XOR2_X1 U355 ( .A(n306), .B(n338), .Z(n307) );
  XOR2_X1 U356 ( .A(n308), .B(n307), .Z(n535) );
  XOR2_X1 U357 ( .A(G99GAT), .B(G85GAT), .Z(n336) );
  XOR2_X1 U358 ( .A(G134GAT), .B(KEYINPUT76), .Z(n389) );
  XOR2_X1 U359 ( .A(n336), .B(n389), .Z(n310) );
  XNOR2_X1 U360 ( .A(G190GAT), .B(G218GAT), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n315) );
  XOR2_X1 U362 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n312) );
  XNOR2_X1 U363 ( .A(KEYINPUT75), .B(KEYINPUT65), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U365 ( .A(G92GAT), .B(KEYINPUT74), .Z(n317) );
  XNOR2_X1 U366 ( .A(G29GAT), .B(G106GAT), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n327) );
  XOR2_X1 U369 ( .A(KEYINPUT7), .B(G50GAT), .Z(n321) );
  XNOR2_X1 U370 ( .A(G43GAT), .B(G36GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U372 ( .A(KEYINPUT8), .B(n322), .Z(n354) );
  XOR2_X1 U373 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n324) );
  XNOR2_X1 U374 ( .A(G162GAT), .B(KEYINPUT77), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n354), .B(n325), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n327), .B(n326), .ZN(n560) );
  NAND2_X1 U378 ( .A1(n535), .A2(n580), .ZN(n331) );
  XOR2_X1 U379 ( .A(G64GAT), .B(G92GAT), .Z(n333) );
  XNOR2_X1 U380 ( .A(G176GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n377) );
  XNOR2_X1 U382 ( .A(n377), .B(KEYINPUT32), .ZN(n335) );
  NAND2_X1 U383 ( .A1(G230GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U385 ( .A(G106GAT), .B(G78GAT), .Z(n412) );
  XNOR2_X1 U386 ( .A(n336), .B(n412), .ZN(n337) );
  XOR2_X1 U387 ( .A(n341), .B(KEYINPUT70), .Z(n347) );
  XOR2_X1 U388 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n343) );
  XNOR2_X1 U389 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n342) );
  XOR2_X1 U390 ( .A(n343), .B(n342), .Z(n345) );
  XOR2_X1 U391 ( .A(G120GAT), .B(G57GAT), .Z(n395) );
  XNOR2_X1 U392 ( .A(G148GAT), .B(n395), .ZN(n344) );
  XOR2_X1 U393 ( .A(G169GAT), .B(G8GAT), .Z(n381) );
  XOR2_X1 U394 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n349) );
  XNOR2_X1 U395 ( .A(G197GAT), .B(KEYINPUT66), .ZN(n348) );
  XNOR2_X1 U396 ( .A(n349), .B(n348), .ZN(n351) );
  XOR2_X1 U397 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U398 ( .A(G1GAT), .B(G141GAT), .Z(n353) );
  XNOR2_X1 U399 ( .A(G29GAT), .B(G113GAT), .ZN(n352) );
  XNOR2_X1 U400 ( .A(n353), .B(n352), .ZN(n388) );
  XNOR2_X1 U401 ( .A(n354), .B(n388), .ZN(n355) );
  XNOR2_X1 U402 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U403 ( .A(n381), .B(n357), .Z(n359) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U405 ( .A(n359), .B(n358), .ZN(n568) );
  XOR2_X1 U406 ( .A(n568), .B(KEYINPUT68), .Z(n558) );
  INV_X1 U407 ( .A(n558), .ZN(n360) );
  AND2_X1 U408 ( .A1(n364), .A2(n360), .ZN(n361) );
  AND2_X1 U409 ( .A1(n362), .A2(n361), .ZN(n363) );
  XNOR2_X1 U410 ( .A(n363), .B(KEYINPUT114), .ZN(n370) );
  INV_X1 U411 ( .A(n560), .ZN(n555) );
  INV_X1 U412 ( .A(n535), .ZN(n578) );
  NAND2_X1 U413 ( .A1(n555), .A2(n578), .ZN(n367) );
  XOR2_X1 U414 ( .A(KEYINPUT41), .B(n364), .Z(n546) );
  NOR2_X1 U415 ( .A1(n568), .A2(n546), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n365), .B(KEYINPUT46), .ZN(n366) );
  NOR2_X1 U417 ( .A1(n367), .A2(n366), .ZN(n368) );
  XOR2_X1 U418 ( .A(KEYINPUT47), .B(n368), .Z(n369) );
  NOR2_X1 U419 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U420 ( .A(n371), .B(KEYINPUT48), .ZN(n526) );
  XOR2_X1 U421 ( .A(KEYINPUT18), .B(G190GAT), .Z(n373) );
  XNOR2_X1 U422 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n372) );
  XNOR2_X1 U423 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U424 ( .A(KEYINPUT17), .B(n374), .ZN(n446) );
  XOR2_X1 U425 ( .A(G211GAT), .B(KEYINPUT21), .Z(n376) );
  XNOR2_X1 U426 ( .A(G197GAT), .B(G218GAT), .ZN(n375) );
  XNOR2_X1 U427 ( .A(n376), .B(n375), .ZN(n415) );
  XNOR2_X1 U428 ( .A(n415), .B(n377), .ZN(n385) );
  XOR2_X1 U429 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n379) );
  XNOR2_X1 U430 ( .A(G36GAT), .B(KEYINPUT95), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U432 ( .A(n381), .B(n380), .Z(n383) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U434 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U435 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U436 ( .A(n446), .B(n386), .Z(n517) );
  NOR2_X1 U437 ( .A1(n526), .A2(n517), .ZN(n387) );
  XNOR2_X1 U438 ( .A(n387), .B(KEYINPUT54), .ZN(n565) );
  XOR2_X1 U439 ( .A(n389), .B(n388), .Z(n391) );
  NAND2_X1 U440 ( .A1(G225GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U441 ( .A(n391), .B(n390), .ZN(n403) );
  XOR2_X1 U442 ( .A(KEYINPUT89), .B(KEYINPUT91), .Z(n393) );
  XNOR2_X1 U443 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n392) );
  XNOR2_X1 U444 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U445 ( .A(n394), .B(KEYINPUT90), .Z(n397) );
  XNOR2_X1 U446 ( .A(n395), .B(G85GAT), .ZN(n396) );
  XNOR2_X1 U447 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U448 ( .A(n398), .B(KEYINPUT1), .Z(n401) );
  XNOR2_X1 U449 ( .A(G127GAT), .B(KEYINPUT0), .ZN(n399) );
  XNOR2_X1 U450 ( .A(n399), .B(KEYINPUT80), .ZN(n438) );
  XNOR2_X1 U451 ( .A(n438), .B(KEYINPUT6), .ZN(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U453 ( .A(n403), .B(n402), .ZN(n408) );
  XNOR2_X1 U454 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n404) );
  XNOR2_X1 U455 ( .A(n404), .B(KEYINPUT88), .ZN(n405) );
  XOR2_X1 U456 ( .A(n405), .B(KEYINPUT3), .Z(n407) );
  XNOR2_X1 U457 ( .A(G148GAT), .B(G162GAT), .ZN(n406) );
  XOR2_X1 U458 ( .A(n407), .B(n406), .Z(n423) );
  XNOR2_X1 U459 ( .A(n408), .B(n423), .ZN(n466) );
  XNOR2_X1 U460 ( .A(KEYINPUT92), .B(n466), .ZN(n564) );
  XOR2_X1 U461 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n410) );
  XNOR2_X1 U462 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U464 ( .A(n411), .B(KEYINPUT74), .Z(n414) );
  XNOR2_X1 U465 ( .A(G50GAT), .B(n412), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n414), .B(n413), .ZN(n419) );
  XOR2_X1 U467 ( .A(G141GAT), .B(n415), .Z(n417) );
  NAND2_X1 U468 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U470 ( .A(n419), .B(n418), .Z(n425) );
  XOR2_X1 U471 ( .A(G204GAT), .B(KEYINPUT24), .Z(n421) );
  XNOR2_X1 U472 ( .A(KEYINPUT23), .B(KEYINPUT86), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U474 ( .A(n423), .B(n422), .Z(n424) );
  XNOR2_X1 U475 ( .A(n425), .B(n424), .ZN(n468) );
  INV_X1 U476 ( .A(n468), .ZN(n426) );
  AND2_X1 U477 ( .A1(n564), .A2(n426), .ZN(n427) );
  AND2_X1 U478 ( .A1(n565), .A2(n427), .ZN(n429) );
  XNOR2_X1 U479 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n428) );
  XNOR2_X1 U480 ( .A(n429), .B(n428), .ZN(n449) );
  XOR2_X1 U481 ( .A(G71GAT), .B(G15GAT), .Z(n431) );
  XNOR2_X1 U482 ( .A(G169GAT), .B(G113GAT), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n431), .B(n430), .ZN(n445) );
  XOR2_X1 U484 ( .A(G176GAT), .B(KEYINPUT82), .Z(n433) );
  XNOR2_X1 U485 ( .A(G134GAT), .B(KEYINPUT84), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U487 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n435) );
  XNOR2_X1 U488 ( .A(G120GAT), .B(KEYINPUT83), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U490 ( .A(n437), .B(n436), .Z(n443) );
  XOR2_X1 U491 ( .A(G99GAT), .B(n438), .Z(n440) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n448) );
  INV_X1 U497 ( .A(n446), .ZN(n447) );
  XOR2_X2 U498 ( .A(n448), .B(n447), .Z(n529) );
  NOR2_X1 U499 ( .A1(n449), .A2(n529), .ZN(n450) );
  XOR2_X1 U500 ( .A(KEYINPUT123), .B(n450), .Z(n561) );
  INV_X1 U501 ( .A(n546), .ZN(n531) );
  NAND2_X1 U502 ( .A1(n561), .A2(n531), .ZN(n453) );
  XOR2_X1 U503 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n451) );
  XNOR2_X1 U504 ( .A(n451), .B(G176GAT), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(G1349GAT) );
  NAND2_X1 U506 ( .A1(n535), .A2(n561), .ZN(n455) );
  XOR2_X1 U507 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n457) );
  XNOR2_X1 U508 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(n477) );
  NAND2_X1 U510 ( .A1(n364), .A2(n558), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(KEYINPUT73), .ZN(n489) );
  NOR2_X1 U512 ( .A1(n529), .A2(n517), .ZN(n459) );
  NOR2_X1 U513 ( .A1(n468), .A2(n459), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT25), .ZN(n464) );
  XOR2_X1 U515 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n461) );
  XOR2_X1 U516 ( .A(n517), .B(n461), .Z(n469) );
  NAND2_X1 U517 ( .A1(n529), .A2(n468), .ZN(n462) );
  XOR2_X1 U518 ( .A(n462), .B(KEYINPUT26), .Z(n542) );
  INV_X1 U519 ( .A(n542), .ZN(n567) );
  OR2_X1 U520 ( .A1(n469), .A2(n567), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n467), .B(KEYINPUT97), .ZN(n473) );
  XOR2_X1 U524 ( .A(n468), .B(KEYINPUT28), .Z(n527) );
  INV_X1 U525 ( .A(n527), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n564), .A2(n469), .ZN(n524) );
  NAND2_X1 U527 ( .A1(n524), .A2(n529), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n486) );
  NOR2_X1 U530 ( .A1(n578), .A2(n560), .ZN(n474) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(n474), .Z(n475) );
  NOR2_X1 U532 ( .A1(n486), .A2(n475), .ZN(n502) );
  NAND2_X1 U533 ( .A1(n489), .A2(n502), .ZN(n482) );
  NOR2_X1 U534 ( .A1(n564), .A2(n482), .ZN(n476) );
  XOR2_X1 U535 ( .A(n477), .B(n476), .Z(G1324GAT) );
  NOR2_X1 U536 ( .A1(n517), .A2(n482), .ZN(n478) );
  XOR2_X1 U537 ( .A(G8GAT), .B(n478), .Z(G1325GAT) );
  NOR2_X1 U538 ( .A1(n529), .A2(n482), .ZN(n480) );
  XNOR2_X1 U539 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(n481), .ZN(G1326GAT) );
  NOR2_X1 U542 ( .A1(n527), .A2(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G22GAT), .B(n485), .ZN(G1327GAT) );
  NOR2_X1 U546 ( .A1(n486), .A2(n535), .ZN(n487) );
  NAND2_X1 U547 ( .A1(n580), .A2(n487), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(n488), .ZN(n514) );
  NAND2_X1 U549 ( .A1(n489), .A2(n514), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(KEYINPUT38), .ZN(n498) );
  NOR2_X1 U551 ( .A1(n498), .A2(n564), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(n492), .ZN(G1328GAT) );
  NOR2_X1 U554 ( .A1(n498), .A2(n517), .ZN(n493) );
  XOR2_X1 U555 ( .A(KEYINPUT104), .B(n493), .Z(n494) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  NOR2_X1 U557 ( .A1(n498), .A2(n529), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n527), .A2(n498), .ZN(n499) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT106), .B(n500), .ZN(G1331GAT) );
  NAND2_X1 U564 ( .A1(n531), .A2(n568), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(KEYINPUT107), .ZN(n513) );
  NAND2_X1 U566 ( .A1(n513), .A2(n502), .ZN(n509) );
  NOR2_X1 U567 ( .A1(n564), .A2(n509), .ZN(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n505), .Z(G1332GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n509), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1333GAT) );
  NOR2_X1 U574 ( .A1(n529), .A2(n509), .ZN(n508) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n508), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n527), .A2(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n521) );
  NOR2_X1 U581 ( .A1(n564), .A2(n521), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n517), .A2(n521), .ZN(n518) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n529), .A2(n521), .ZN(n519) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(n519), .Z(n520) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n520), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n527), .A2(n521), .ZN(n522) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(n522), .Z(n523) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  INV_X1 U592 ( .A(n524), .ZN(n525) );
  NOR2_X1 U593 ( .A1(n526), .A2(n525), .ZN(n543) );
  NAND2_X1 U594 ( .A1(n527), .A2(n543), .ZN(n528) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n558), .A2(n539), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U599 ( .A1(n539), .A2(n531), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U601 ( .A(G120GAT), .B(n534), .Z(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n537) );
  NAND2_X1 U603 ( .A1(n539), .A2(n535), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U605 ( .A(G127GAT), .B(n538), .Z(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U607 ( .A1(n539), .A2(n560), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n554) );
  NOR2_X1 U610 ( .A1(n568), .A2(n554), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1344GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n554), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n548) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(KEYINPUT52), .B(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n578), .A2(n554), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT120), .B(n552), .Z(n553) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1351GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n581) );
  INV_X1 U632 ( .A(n581), .ZN(n577) );
  NOR2_X1 U633 ( .A1(n568), .A2(n577), .ZN(n573) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT59), .B(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n364), .A2(n577), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

