

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601;

  XNOR2_X1 U324 ( .A(n327), .B(n292), .ZN(n331) );
  XNOR2_X1 U325 ( .A(n368), .B(KEYINPUT67), .ZN(n379) );
  XNOR2_X1 U326 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U327 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U328 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U329 ( .A(n509), .B(KEYINPUT37), .ZN(n510) );
  XOR2_X1 U330 ( .A(n326), .B(n325), .Z(n292) );
  XOR2_X1 U331 ( .A(n450), .B(n449), .Z(n293) );
  XOR2_X1 U332 ( .A(n356), .B(n426), .Z(n294) );
  XOR2_X1 U333 ( .A(G190GAT), .B(n444), .Z(n295) );
  XOR2_X1 U334 ( .A(KEYINPUT47), .B(n405), .Z(n296) );
  NOR2_X1 U335 ( .A1(n561), .A2(n400), .ZN(n402) );
  NOR2_X1 U336 ( .A1(n497), .A2(n487), .ZN(n474) );
  XNOR2_X1 U337 ( .A(G22GAT), .B(G15GAT), .ZN(n368) );
  INV_X1 U338 ( .A(G36GAT), .ZN(n380) );
  XNOR2_X1 U339 ( .A(n369), .B(KEYINPUT15), .ZN(n370) );
  INV_X1 U340 ( .A(KEYINPUT98), .ZN(n509) );
  XNOR2_X1 U341 ( .A(n451), .B(n293), .ZN(n452) );
  NAND2_X1 U342 ( .A1(n422), .A2(n541), .ZN(n423) );
  XNOR2_X1 U343 ( .A(n383), .B(n382), .ZN(n391) );
  XNOR2_X1 U344 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U345 ( .A(n423), .B(KEYINPUT54), .ZN(n424) );
  XNOR2_X1 U346 ( .A(n511), .B(n510), .ZN(n537) );
  XNOR2_X1 U347 ( .A(n377), .B(n376), .ZN(n593) );
  XNOR2_X1 U348 ( .A(n395), .B(n394), .ZN(n581) );
  XOR2_X1 U349 ( .A(n483), .B(KEYINPUT28), .Z(n553) );
  XNOR2_X1 U350 ( .A(KEYINPUT99), .B(n514), .ZN(n523) );
  XNOR2_X1 U351 ( .A(n470), .B(KEYINPUT58), .ZN(n471) );
  XNOR2_X1 U352 ( .A(n472), .B(n471), .ZN(G1351GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n298) );
  XNOR2_X1 U354 ( .A(KEYINPUT5), .B(KEYINPUT88), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U356 ( .A(KEYINPUT4), .B(n299), .Z(n301) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U359 ( .A(n302), .B(KEYINPUT86), .Z(n309) );
  XOR2_X1 U360 ( .A(G120GAT), .B(G148GAT), .Z(n326) );
  XOR2_X1 U361 ( .A(KEYINPUT85), .B(n326), .Z(n306) );
  XOR2_X1 U362 ( .A(G57GAT), .B(G155GAT), .Z(n304) );
  XNOR2_X1 U363 ( .A(G1GAT), .B(G127GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n304), .B(n303), .ZN(n362) );
  XNOR2_X1 U365 ( .A(G162GAT), .B(n362), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n307), .B(KEYINPUT87), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n311) );
  XNOR2_X1 U369 ( .A(G29GAT), .B(G134GAT), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n310), .B(G85GAT), .ZN(n352) );
  XOR2_X1 U371 ( .A(n311), .B(n352), .Z(n318) );
  XNOR2_X1 U372 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n312), .B(KEYINPUT77), .ZN(n444) );
  XNOR2_X1 U374 ( .A(KEYINPUT2), .B(KEYINPUT83), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n313), .B(KEYINPUT82), .ZN(n314) );
  XOR2_X1 U376 ( .A(n314), .B(KEYINPUT3), .Z(n316) );
  XNOR2_X1 U377 ( .A(G141GAT), .B(KEYINPUT81), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n316), .B(n315), .ZN(n440) );
  XNOR2_X1 U379 ( .A(n444), .B(n440), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n481) );
  XNOR2_X1 U381 ( .A(KEYINPUT89), .B(n481), .ZN(n485) );
  XOR2_X1 U382 ( .A(KEYINPUT32), .B(KEYINPUT68), .Z(n320) );
  XNOR2_X1 U383 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n333) );
  XOR2_X1 U385 ( .A(G71GAT), .B(KEYINPUT13), .Z(n373) );
  XOR2_X1 U386 ( .A(n373), .B(G92GAT), .Z(n322) );
  XOR2_X1 U387 ( .A(G176GAT), .B(G64GAT), .Z(n413) );
  XNOR2_X1 U388 ( .A(G85GAT), .B(n413), .ZN(n321) );
  XNOR2_X1 U389 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U390 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n324) );
  XNOR2_X1 U391 ( .A(KEYINPUT72), .B(KEYINPUT31), .ZN(n323) );
  XNOR2_X1 U392 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U393 ( .A(G99GAT), .B(G106GAT), .Z(n356) );
  XNOR2_X1 U394 ( .A(G78GAT), .B(KEYINPUT70), .ZN(n328) );
  XNOR2_X1 U395 ( .A(n328), .B(G204GAT), .ZN(n426) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U397 ( .A(n294), .B(n329), .ZN(n330) );
  XOR2_X1 U398 ( .A(n333), .B(n332), .Z(n587) );
  INV_X1 U399 ( .A(KEYINPUT7), .ZN(n334) );
  NAND2_X1 U400 ( .A1(G43GAT), .A2(n334), .ZN(n337) );
  INV_X1 U401 ( .A(G43GAT), .ZN(n335) );
  NAND2_X1 U402 ( .A1(n335), .A2(KEYINPUT7), .ZN(n336) );
  NAND2_X1 U403 ( .A1(n337), .A2(n336), .ZN(n339) );
  XNOR2_X1 U404 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n393) );
  XOR2_X1 U406 ( .A(n393), .B(KEYINPUT64), .Z(n341) );
  NAND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U408 ( .A(n341), .B(n340), .ZN(n347) );
  INV_X1 U409 ( .A(n347), .ZN(n345) );
  XOR2_X1 U410 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n343) );
  XNOR2_X1 U411 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n342) );
  XNOR2_X1 U412 ( .A(n343), .B(n342), .ZN(n346) );
  INV_X1 U413 ( .A(n346), .ZN(n344) );
  NAND2_X1 U414 ( .A1(n345), .A2(n344), .ZN(n349) );
  NAND2_X1 U415 ( .A1(n347), .A2(n346), .ZN(n348) );
  NAND2_X1 U416 ( .A1(n349), .A2(n348), .ZN(n354) );
  XOR2_X1 U417 ( .A(G92GAT), .B(G218GAT), .Z(n351) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G190GAT), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n410) );
  XOR2_X1 U420 ( .A(n352), .B(n410), .Z(n353) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U422 ( .A(G50GAT), .B(G162GAT), .Z(n425) );
  XNOR2_X1 U423 ( .A(n355), .B(n425), .ZN(n358) );
  INV_X1 U424 ( .A(n356), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n358), .B(n357), .ZN(n403) );
  XNOR2_X1 U426 ( .A(KEYINPUT74), .B(n403), .ZN(n565) );
  XNOR2_X1 U427 ( .A(KEYINPUT36), .B(n565), .ZN(n598) );
  XOR2_X1 U428 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n360) );
  XNOR2_X1 U429 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n359) );
  XOR2_X1 U430 ( .A(n360), .B(n359), .Z(n377) );
  INV_X1 U431 ( .A(n362), .ZN(n361) );
  XOR2_X1 U432 ( .A(G8GAT), .B(G183GAT), .Z(n416) );
  NAND2_X1 U433 ( .A1(n361), .A2(n416), .ZN(n365) );
  INV_X1 U434 ( .A(n416), .ZN(n363) );
  NAND2_X1 U435 ( .A1(n363), .A2(n362), .ZN(n364) );
  NAND2_X1 U436 ( .A1(n365), .A2(n364), .ZN(n367) );
  NAND2_X1 U437 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U438 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U439 ( .A(n379), .B(KEYINPUT12), .Z(n369) );
  XOR2_X1 U440 ( .A(n373), .B(n372), .Z(n375) );
  XNOR2_X1 U441 ( .A(G211GAT), .B(G78GAT), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n375), .B(n374), .ZN(n376) );
  NOR2_X1 U443 ( .A1(n598), .A2(n593), .ZN(n378) );
  XNOR2_X1 U444 ( .A(KEYINPUT45), .B(n378), .ZN(n396) );
  XOR2_X1 U445 ( .A(G29GAT), .B(n379), .Z(n383) );
  NAND2_X1 U446 ( .A1(G229GAT), .A2(G233GAT), .ZN(n381) );
  XOR2_X1 U447 ( .A(G141GAT), .B(G197GAT), .Z(n385) );
  XNOR2_X1 U448 ( .A(G169GAT), .B(G50GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U450 ( .A(KEYINPUT29), .B(G1GAT), .Z(n387) );
  XNOR2_X1 U451 ( .A(G113GAT), .B(G8GAT), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U455 ( .A(n392), .B(KEYINPUT65), .Z(n395) );
  XNOR2_X1 U456 ( .A(n393), .B(KEYINPUT30), .ZN(n394) );
  NAND2_X1 U457 ( .A1(n396), .A2(n581), .ZN(n397) );
  NOR2_X1 U458 ( .A1(n587), .A2(n397), .ZN(n398) );
  XOR2_X1 U459 ( .A(KEYINPUT113), .B(n398), .Z(n406) );
  XNOR2_X1 U460 ( .A(KEYINPUT111), .B(n593), .ZN(n561) );
  XNOR2_X1 U461 ( .A(KEYINPUT41), .B(n587), .ZN(n571) );
  NOR2_X1 U462 ( .A1(n581), .A2(n571), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n399), .B(KEYINPUT46), .ZN(n400) );
  INV_X1 U464 ( .A(KEYINPUT112), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n402), .B(n401), .ZN(n404) );
  INV_X1 U466 ( .A(n403), .ZN(n576) );
  NOR2_X1 U467 ( .A1(n404), .A2(n576), .ZN(n405) );
  NOR2_X1 U468 ( .A1(n406), .A2(n296), .ZN(n407) );
  XNOR2_X1 U469 ( .A(KEYINPUT48), .B(n407), .ZN(n551) );
  INV_X1 U470 ( .A(n551), .ZN(n422) );
  XOR2_X1 U471 ( .A(G211GAT), .B(KEYINPUT80), .Z(n409) );
  XNOR2_X1 U472 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n430) );
  XNOR2_X1 U474 ( .A(n430), .B(n410), .ZN(n421) );
  XOR2_X1 U475 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n412) );
  XNOR2_X1 U476 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n455) );
  XOR2_X1 U478 ( .A(n455), .B(n413), .Z(n415) );
  NAND2_X1 U479 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U480 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U481 ( .A(n417), .B(n416), .Z(n419) );
  XNOR2_X1 U482 ( .A(G204GAT), .B(KEYINPUT90), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n497) );
  NOR2_X1 U485 ( .A1(n485), .A2(n424), .ZN(n580) );
  XOR2_X1 U486 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U489 ( .A(n429), .B(KEYINPUT79), .Z(n432) );
  XNOR2_X1 U490 ( .A(n430), .B(KEYINPUT22), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U492 ( .A(KEYINPUT84), .B(G155GAT), .Z(n434) );
  XNOR2_X1 U493 ( .A(G218GAT), .B(G106GAT), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U495 ( .A(n436), .B(n435), .Z(n442) );
  XOR2_X1 U496 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n438) );
  XNOR2_X1 U497 ( .A(G22GAT), .B(G148GAT), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n483) );
  NAND2_X1 U501 ( .A1(n580), .A2(n483), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n443), .B(KEYINPUT55), .ZN(n458) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n295), .B(n445), .ZN(n453) );
  XOR2_X1 U505 ( .A(G183GAT), .B(G99GAT), .Z(n447) );
  XNOR2_X1 U506 ( .A(G15GAT), .B(G134GAT), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U508 ( .A(G43GAT), .B(n448), .ZN(n451) );
  XOR2_X1 U509 ( .A(G71GAT), .B(KEYINPUT20), .Z(n450) );
  XNOR2_X1 U510 ( .A(G176GAT), .B(KEYINPUT78), .ZN(n449) );
  XOR2_X1 U511 ( .A(n454), .B(G120GAT), .Z(n457) );
  XNOR2_X1 U512 ( .A(n455), .B(G127GAT), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(n473) );
  NAND2_X1 U514 ( .A1(n458), .A2(n473), .ZN(n469) );
  NOR2_X1 U515 ( .A1(n469), .A2(n581), .ZN(n461) );
  XNOR2_X1 U516 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n459), .B(G169GAT), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n461), .B(n460), .ZN(G1348GAT) );
  INV_X1 U519 ( .A(n469), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n462), .A2(n561), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(G183GAT), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n465), .B(n464), .ZN(G1350GAT) );
  NOR2_X1 U524 ( .A1(n571), .A2(n469), .ZN(n468) );
  XNOR2_X1 U525 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n466), .B(G176GAT), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(G1349GAT) );
  NOR2_X1 U528 ( .A1(n565), .A2(n469), .ZN(n472) );
  INV_X1 U529 ( .A(G190GAT), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n581), .A2(n587), .ZN(n512) );
  INV_X1 U531 ( .A(n473), .ZN(n487) );
  XOR2_X1 U532 ( .A(KEYINPUT92), .B(n474), .Z(n475) );
  NAND2_X1 U533 ( .A1(n483), .A2(n475), .ZN(n477) );
  XNOR2_X1 U534 ( .A(KEYINPUT25), .B(KEYINPUT93), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n480) );
  XOR2_X1 U536 ( .A(n497), .B(KEYINPUT27), .Z(n484) );
  NOR2_X1 U537 ( .A1(n483), .A2(n473), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(KEYINPUT26), .ZN(n579) );
  NAND2_X1 U539 ( .A1(n484), .A2(n579), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n480), .A2(n479), .ZN(n482) );
  NAND2_X1 U541 ( .A1(n482), .A2(n481), .ZN(n490) );
  NAND2_X1 U542 ( .A1(n485), .A2(n484), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT91), .B(n486), .Z(n550) );
  NOR2_X1 U544 ( .A1(n553), .A2(n550), .ZN(n488) );
  NAND2_X1 U545 ( .A1(n488), .A2(n487), .ZN(n489) );
  NAND2_X1 U546 ( .A1(n490), .A2(n489), .ZN(n507) );
  INV_X1 U547 ( .A(n593), .ZN(n491) );
  NAND2_X1 U548 ( .A1(n565), .A2(n491), .ZN(n492) );
  XOR2_X1 U549 ( .A(KEYINPUT16), .B(n492), .Z(n493) );
  NAND2_X1 U550 ( .A1(n507), .A2(n493), .ZN(n494) );
  XOR2_X1 U551 ( .A(KEYINPUT94), .B(n494), .Z(n527) );
  AND2_X1 U552 ( .A1(n512), .A2(n527), .ZN(n502) );
  NAND2_X1 U553 ( .A1(n502), .A2(n485), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT34), .B(n495), .ZN(n496) );
  XNOR2_X1 U555 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  XOR2_X1 U556 ( .A(G8GAT), .B(KEYINPUT95), .Z(n499) );
  INV_X1 U557 ( .A(n497), .ZN(n541) );
  NAND2_X1 U558 ( .A1(n502), .A2(n541), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1325GAT) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .Z(n501) );
  NAND2_X1 U561 ( .A1(n502), .A2(n473), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(G1326GAT) );
  NAND2_X1 U563 ( .A1(n502), .A2(n553), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(KEYINPUT96), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G22GAT), .B(n504), .ZN(G1327GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT97), .B(KEYINPUT100), .Z(n506) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n516) );
  NAND2_X1 U569 ( .A1(n593), .A2(n507), .ZN(n508) );
  NOR2_X1 U570 ( .A1(n598), .A2(n508), .ZN(n511) );
  NAND2_X1 U571 ( .A1(n537), .A2(n512), .ZN(n513) );
  XNOR2_X1 U572 ( .A(n513), .B(KEYINPUT38), .ZN(n514) );
  NAND2_X1 U573 ( .A1(n523), .A2(n485), .ZN(n515) );
  XOR2_X1 U574 ( .A(n516), .B(n515), .Z(G1328GAT) );
  XOR2_X1 U575 ( .A(G36GAT), .B(KEYINPUT101), .Z(n518) );
  NAND2_X1 U576 ( .A1(n523), .A2(n541), .ZN(n517) );
  XNOR2_X1 U577 ( .A(n518), .B(n517), .ZN(G1329GAT) );
  XNOR2_X1 U578 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n522) );
  XOR2_X1 U579 ( .A(KEYINPUT102), .B(KEYINPUT40), .Z(n520) );
  NAND2_X1 U580 ( .A1(n473), .A2(n523), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U582 ( .A(n522), .B(n521), .ZN(G1330GAT) );
  NAND2_X1 U583 ( .A1(n523), .A2(n553), .ZN(n524) );
  XNOR2_X1 U584 ( .A(n524), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n530) );
  INV_X1 U586 ( .A(n581), .ZN(n525) );
  NOR2_X1 U587 ( .A1(n571), .A2(n525), .ZN(n526) );
  XNOR2_X1 U588 ( .A(n526), .B(KEYINPUT104), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n527), .A2(n538), .ZN(n528) );
  XNOR2_X1 U590 ( .A(n528), .B(KEYINPUT105), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n534), .A2(n485), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U593 ( .A(G57GAT), .B(n531), .Z(G1332GAT) );
  NAND2_X1 U594 ( .A1(n541), .A2(n534), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n532), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U596 ( .A1(n534), .A2(n473), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U598 ( .A(G78GAT), .B(KEYINPUT43), .Z(n536) );
  NAND2_X1 U599 ( .A1(n534), .A2(n553), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1335GAT) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n539), .B(KEYINPUT107), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n546), .A2(n485), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G85GAT), .B(n540), .ZN(G1336GAT) );
  NAND2_X1 U605 ( .A1(n541), .A2(n546), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(KEYINPUT108), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G92GAT), .B(n543), .ZN(G1337GAT) );
  XOR2_X1 U608 ( .A(G99GAT), .B(KEYINPUT109), .Z(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n473), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1338GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n548) );
  NAND2_X1 U612 ( .A1(n546), .A2(n553), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U614 ( .A(G106GAT), .B(n549), .Z(G1339GAT) );
  NOR2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT114), .B(n552), .Z(n568) );
  NOR2_X1 U617 ( .A1(n568), .A2(n553), .ZN(n554) );
  NAND2_X1 U618 ( .A1(n473), .A2(n554), .ZN(n564) );
  NOR2_X1 U619 ( .A1(n581), .A2(n564), .ZN(n556) );
  XNOR2_X1 U620 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(G1340GAT) );
  NOR2_X1 U622 ( .A1(n571), .A2(n564), .ZN(n558) );
  XNOR2_X1 U623 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G120GAT), .B(n559), .ZN(G1341GAT) );
  INV_X1 U626 ( .A(n564), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT50), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G127GAT), .B(n563), .ZN(G1342GAT) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1343GAT) );
  INV_X1 U633 ( .A(n568), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n579), .A2(n569), .ZN(n577) );
  NOR2_X1 U635 ( .A1(n581), .A2(n577), .ZN(n570) );
  XOR2_X1 U636 ( .A(G141GAT), .B(n570), .Z(G1344GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n577), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G148GAT), .B(n574), .ZN(G1345GAT) );
  NOR2_X1 U641 ( .A1(n593), .A2(n577), .ZN(n575) );
  XOR2_X1 U642 ( .A(G155GAT), .B(n575), .Z(G1346GAT) );
  NOR2_X1 U643 ( .A1(n403), .A2(n577), .ZN(n578) );
  XOR2_X1 U644 ( .A(G162GAT), .B(n578), .Z(G1347GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n597) );
  NOR2_X1 U646 ( .A1(n581), .A2(n597), .ZN(n586) );
  XOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT122), .Z(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(KEYINPUT121), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(KEYINPUT59), .B(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  INV_X1 U652 ( .A(n587), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n597), .A2(n588), .ZN(n592) );
  XOR2_X1 U654 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n590) );
  XNOR2_X1 U655 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(G1353GAT) );
  NOR2_X1 U658 ( .A1(n593), .A2(n597), .ZN(n595) );
  XNOR2_X1 U659 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n594) );
  XNOR2_X1 U660 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U661 ( .A(G211GAT), .B(n596), .ZN(G1354GAT) );
  NOR2_X1 U662 ( .A1(n598), .A2(n597), .ZN(n600) );
  XNOR2_X1 U663 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n599) );
  XNOR2_X1 U664 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U665 ( .A(G218GAT), .B(n601), .ZN(G1355GAT) );
endmodule

